* NGSPICE file created from lovers_controller.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

.subckt lovers_controller becStatus[0] becStatus[1] becStatus[2] becStatus[3] data_in[0]
+ data_in[10] data_in[11] data_in[12] data_in[13] data_in[14] data_in[15] data_in[16]
+ data_in[17] data_in[18] data_in[19] data_in[1] data_in[20] data_in[21] data_in[22]
+ data_in[23] data_in[24] data_in[25] data_in[26] data_in[27] data_in[28] data_in[29]
+ data_in[2] data_in[30] data_in[31] data_in[3] data_in[4] data_in[5] data_in[6] data_in[7]
+ data_in[8] data_in[9] data_out[0] data_out[10] data_out[11] data_out[12] data_out[13]
+ data_out[14] data_out[15] data_out[16] data_out[17] data_out[18] data_out[19] data_out[1]
+ data_out[20] data_out[21] data_out[22] data_out[23] data_out[24] data_out[25] data_out[26]
+ data_out[27] data_out[28] data_out[29] data_out[2] data_out[30] data_out[31] data_out[3]
+ data_out[4] data_out[5] data_out[6] data_out[7] data_out[8] data_out[9] io_oeb io_out
+ ki la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[3] la_data_in[4] la_data_in[5] la_data_in[6] la_data_in[7]
+ la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[3]
+ la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9]
+ load_data load_status[0] load_status[1] load_status[2] load_status[3] load_status[4]
+ load_status[5] next_key slv_done slv_enable vccd1 vssd1 wb_clk_i wb_rst_i
XFILLER_0_236_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09671_ _18294_/Q hold3545/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09672_/B sky130_fd_sc_hd__mux2_1
X_08622_ _15314_/A hold762/X vssd1 vssd1 vccd1 vccd1 _15933_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_234_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08553_ _12420_/A _08553_/B vssd1 vssd1 vccd1 vccd1 _15900_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08484_ _15163_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _08484_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_175_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09105_ hold2447/X _09106_/B _09104_/Y _12987_/A vssd1 vssd1 vccd1 vccd1 _09105_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09036_ hold245/X hold760/X _09060_/S vssd1 vssd1 vccd1 vccd1 _09037_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold340 hold340/A vssd1 vssd1 vccd1 vccd1 hold340/X sky130_fd_sc_hd__buf_8
XFILLER_0_104_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold351 hold351/A vssd1 vssd1 vccd1 vccd1 input60/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold362 hold362/A vssd1 vssd1 vccd1 vccd1 hold362/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold373 hold47/X vssd1 vssd1 vccd1 vccd1 hold373/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold384 hold384/A vssd1 vssd1 vccd1 vccd1 hold384/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_229_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold395 hold395/A vssd1 vssd1 vccd1 vccd1 hold395/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout820 _10564_/C1 vssd1 vssd1 vccd1 vccd1 _14895_/C1 sky130_fd_sc_hd__buf_4
Xfanout831 _14893_/C1 vssd1 vssd1 vccd1 vccd1 _14769_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_110_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout842 fanout843/X vssd1 vssd1 vccd1 vccd1 _14865_/C1 sky130_fd_sc_hd__clkbuf_4
X_09938_ hold3087/X _16470_/Q _10022_/C vssd1 vssd1 vccd1 vccd1 _09939_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_217_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout853 _11218_/A vssd1 vssd1 vccd1 vccd1 _11206_/A sky130_fd_sc_hd__buf_8
Xfanout864 _15161_/A vssd1 vssd1 vccd1 vccd1 _15215_/A sky130_fd_sc_hd__buf_12
Xfanout875 hold704/X vssd1 vssd1 vccd1 vccd1 _09438_/B sky130_fd_sc_hd__buf_4
XFILLER_0_204_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout886 _15195_/A vssd1 vssd1 vccd1 vccd1 _14461_/A sky130_fd_sc_hd__buf_6
X_09869_ _18360_/Q hold3604/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09870_/B sky130_fd_sc_hd__mux2_1
Xfanout897 _14850_/A vssd1 vssd1 vccd1 vccd1 _15189_/A sky130_fd_sc_hd__clkbuf_16
Xhold1040 _07846_/X vssd1 vssd1 vccd1 vccd1 _15568_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1051 _15811_/Q vssd1 vssd1 vccd1 vccd1 hold1051/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1062 _17516_/Q vssd1 vssd1 vccd1 vccd1 hold1062/X sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ hold1241/X hold4022/X _13796_/S vssd1 vssd1 vccd1 vccd1 _11901_/B sky130_fd_sc_hd__mux2_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1073 _14983_/X vssd1 vssd1 vccd1 vccd1 _18277_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_6_25_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_25_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ hold1909/X _17471_/Q _12916_/S vssd1 vssd1 vccd1 vccd1 _12880_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1084 _15826_/Q vssd1 vssd1 vccd1 vccd1 hold1084/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1095 _18228_/Q vssd1 vssd1 vccd1 vccd1 hold1095/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ hold2966/X hold4343/X _13409_/S vssd1 vssd1 vccd1 vccd1 _11832_/B sky130_fd_sc_hd__mux2_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ hold6062/X _14537_/B hold821/X _13897_/A vssd1 vssd1 vccd1 vccd1 hold822/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11762_/A _11771_/B _12242_/S vssd1 vssd1 vccd1 vccd1 _11762_/X sky130_fd_sc_hd__and3_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ hold5587/X _13883_/B _13500_/X _08347_/A vssd1 vssd1 vccd1 vccd1 _13501_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10713_ _11103_/A _10713_/B vssd1 vssd1 vccd1 vccd1 _10713_/X sky130_fd_sc_hd__or2_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14481_ _15215_/A _14481_/B vssd1 vssd1 vccd1 vccd1 _14481_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_181_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ hold2609/X _17055_/Q _11789_/C vssd1 vssd1 vccd1 vccd1 _11694_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_344_wb_clk_i clkbuf_6_42_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17746_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16220_ _17452_/CLK _16220_/D vssd1 vssd1 vccd1 vccd1 _16220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13432_ hold5819/X _13808_/B _13431_/X _12738_/A vssd1 vssd1 vccd1 vccd1 _13432_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10644_ hold4227/X _10551_/A _10643_/X vssd1 vssd1 vccd1 vccd1 _10644_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16151_ _17491_/CLK _16151_/D vssd1 vssd1 vccd1 vccd1 _16151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10575_ hold4330/X _10986_/A _10574_/X vssd1 vssd1 vccd1 vccd1 _10575_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13363_ hold5502/X _13847_/B _13362_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13363_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15102_ hold6060/X hold340/X hold692/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 hold693/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12314_ _17262_/Q _12356_/B _13481_/S vssd1 vssd1 vccd1 vccd1 _12314_/X sky130_fd_sc_hd__and3_1
X_16082_ _16082_/CLK _16082_/D vssd1 vssd1 vccd1 vccd1 hold567/A sky130_fd_sc_hd__dfxtp_1
X_13294_ _13294_/A _13294_/B vssd1 vssd1 vccd1 vccd1 _13294_/X sky130_fd_sc_hd__or2_1
XFILLER_0_11_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15033_ _14980_/A hold2596/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15034_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12245_ hold2539/X hold4037/X _12371_/C vssd1 vssd1 vccd1 vccd1 _12246_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12176_ hold1825/X hold5137/X _13886_/C vssd1 vssd1 vccd1 vccd1 _12177_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_235_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11127_ _11127_/A _11127_/B vssd1 vssd1 vccd1 vccd1 _11127_/X sky130_fd_sc_hd__or2_1
X_16984_ _17832_/CLK _16984_/D vssd1 vssd1 vccd1 vccd1 _16984_/Q sky130_fd_sc_hd__dfxtp_1
X_15935_ _16120_/CLK _15935_/D vssd1 vssd1 vccd1 vccd1 hold585/A sky130_fd_sc_hd__dfxtp_1
X_11058_ _11136_/A _11058_/B vssd1 vssd1 vccd1 vccd1 _11058_/X sky130_fd_sc_hd__or2_1
XTAP_5160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_60_wb_clk_i clkbuf_6_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18046_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10009_ _11203_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _10009_/Y sky130_fd_sc_hd__nor2_1
XTAP_5193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15866_ _17737_/CLK _15866_/D vssd1 vssd1 vccd1 vccd1 _15866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14817_ hold2027/X _14828_/B _14816_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _14817_/X
+ sky130_fd_sc_hd__o211a_1
X_17605_ _17733_/CLK _17605_/D vssd1 vssd1 vccd1 vccd1 _17605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_231_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15797_ _17728_/CLK _15797_/D vssd1 vssd1 vccd1 vccd1 _15797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17536_ _18372_/CLK _17536_/D vssd1 vssd1 vccd1 vccd1 _17536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14748_ _15195_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14748_/X sky130_fd_sc_hd__or2_1
XFILLER_0_188_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17467_ _17477_/CLK _17467_/D vssd1 vssd1 vccd1 vccd1 _17467_/Q sky130_fd_sc_hd__dfxtp_1
X_14679_ hold1029/X _14666_/B _14678_/X _14697_/C1 vssd1 vssd1 vccd1 vccd1 _14679_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16418_ _18363_/CLK _16418_/D vssd1 vssd1 vccd1 vccd1 _16418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17398_ _18451_/CLK _17398_/D vssd1 vssd1 vccd1 vccd1 _17398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6007 _17554_/Q vssd1 vssd1 vccd1 vccd1 hold6007/X sky130_fd_sc_hd__dlygate4sd3_1
X_16349_ _18262_/CLK _16349_/D vssd1 vssd1 vccd1 vccd1 _16349_/Q sky130_fd_sc_hd__dfxtp_1
Xhold6018 _17551_/Q vssd1 vssd1 vccd1 vccd1 hold6018/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6029 _17557_/Q vssd1 vssd1 vccd1 vccd1 hold6029/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5306 _11989_/X vssd1 vssd1 vccd1 vccd1 _17153_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5317 _16765_/Q vssd1 vssd1 vccd1 vccd1 hold5317/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5328 _10852_/X vssd1 vssd1 vccd1 vccd1 _16774_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5339 _16862_/Q vssd1 vssd1 vccd1 vccd1 hold5339/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4605 _09616_/X vssd1 vssd1 vccd1 vccd1 _16362_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18019_ _18019_/CLK _18019_/D vssd1 vssd1 vccd1 vccd1 _18019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4616 _16779_/Q vssd1 vssd1 vccd1 vccd1 hold4616/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4627 _10453_/X vssd1 vssd1 vccd1 vccd1 _16641_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4638 _16473_/Q vssd1 vssd1 vccd1 vccd1 hold4638/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3904 _09682_/X vssd1 vssd1 vccd1 vccd1 _16384_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4649 _09934_/X vssd1 vssd1 vccd1 vccd1 _16468_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_227_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3915 _16616_/Q vssd1 vssd1 vccd1 vccd1 hold3915/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3926 _09586_/X vssd1 vssd1 vccd1 vccd1 _16352_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3937 _17448_/Q vssd1 vssd1 vccd1 vccd1 hold3937/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3948 _16634_/Q vssd1 vssd1 vccd1 vccd1 hold3948/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3959 _11032_/X vssd1 vssd1 vccd1 vccd1 _16834_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout149 _12749_/S vssd1 vssd1 vccd1 vccd1 _12812_/S sky130_fd_sc_hd__buf_4
X_07984_ _15553_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07984_/X sky130_fd_sc_hd__or2_1
X_09723_ _09981_/A _09723_/B vssd1 vssd1 vccd1 vccd1 _09723_/X sky130_fd_sc_hd__or2_1
XFILLER_0_241_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09654_ _09954_/A _09654_/B vssd1 vssd1 vccd1 vccd1 _09654_/X sky130_fd_sc_hd__or2_1
XFILLER_0_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08605_ hold684/X hold886/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold887/A sky130_fd_sc_hd__mux2_1
X_09585_ _10476_/A _09585_/B vssd1 vssd1 vccd1 vccd1 _09585_/X sky130_fd_sc_hd__or2_1
XFILLER_0_194_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08536_ hold131/X hold735/X _08592_/S vssd1 vssd1 vccd1 vccd1 hold736/A sky130_fd_sc_hd__mux2_1
XFILLER_0_166_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_212_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08467_ hold2246/X _08488_/B _08466_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _08467_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08398_ hold1594/X _08442_/A2 _08397_/X _13417_/C1 vssd1 vssd1 vccd1 vccd1 _08398_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10360_ hold4482/X _10646_/B _10359_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _10360_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09019_ _12426_/A hold776/X vssd1 vssd1 vccd1 vccd1 _16126_/D sky130_fd_sc_hd__and2_1
Xhold5840 _09886_/X vssd1 vssd1 vccd1 vccd1 _16452_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5851 hold6008/X vssd1 vssd1 vccd1 vccd1 _13161_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10291_ hold3284/X _10601_/B _10290_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10291_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5862 output75/X vssd1 vssd1 vccd1 vccd1 data_out[12] sky130_fd_sc_hd__buf_12
XFILLER_0_143_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5873 hold6020/X vssd1 vssd1 vccd1 vccd1 _13225_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12030_ _12285_/A _12030_/B vssd1 vssd1 vccd1 vccd1 _12030_/X sky130_fd_sc_hd__or2_1
Xhold5884 output82/X vssd1 vssd1 vccd1 vccd1 data_out[19] sky130_fd_sc_hd__buf_12
XFILLER_0_130_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5895 _17525_/Q vssd1 vssd1 vccd1 vccd1 hold5895/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold170 hold170/A vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold181 hold181/A vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 hold678/X vssd1 vssd1 vccd1 vccd1 hold679/A sky130_fd_sc_hd__buf_1
XFILLER_0_178_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout650 _12855_/A vssd1 vssd1 vccd1 vccd1 _12873_/A sky130_fd_sc_hd__buf_4
Xfanout661 _12588_/A vssd1 vssd1 vccd1 vccd1 _14364_/A sky130_fd_sc_hd__buf_2
Xfanout672 _08351_/A vssd1 vssd1 vccd1 vccd1 _08373_/A sky130_fd_sc_hd__buf_4
XFILLER_0_233_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout683 _13905_/A vssd1 vssd1 vccd1 vccd1 _14211_/C1 sky130_fd_sc_hd__buf_4
X_13981_ hold2798/X _13986_/B _13980_/Y _13935_/A vssd1 vssd1 vccd1 vccd1 _13981_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout694 _15284_/A vssd1 vssd1 vccd1 vccd1 _12390_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_233_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15720_ _17127_/CLK _15720_/D vssd1 vssd1 vccd1 vccd1 _15720_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ hold4503/X _12931_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12933_/B sky130_fd_sc_hd__mux2_1
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15651_ _17878_/CLK _15651_/D vssd1 vssd1 vccd1 vccd1 _15651_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ hold3353/X _12862_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12864_/B sky130_fd_sc_hd__mux2_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14602_ _15103_/A _14622_/B vssd1 vssd1 vccd1 vccd1 _14602_/X sky130_fd_sc_hd__or2_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ _18370_/CLK _18370_/D vssd1 vssd1 vccd1 vccd1 _18370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11814_ _12198_/A _11814_/B vssd1 vssd1 vccd1 vccd1 _11814_/X sky130_fd_sc_hd__or2_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15582_ _17250_/CLK _15582_/D vssd1 vssd1 vccd1 vccd1 _15582_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ hold3540/X _12793_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12795_/B sky130_fd_sc_hd__mux2_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _17321_/CLK hold148/X vssd1 vssd1 vccd1 vccd1 _17321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14533_ _14604_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14533_/X sky130_fd_sc_hd__or2_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11745_ hold4644/X _12285_/A _11744_/X vssd1 vssd1 vccd1 vccd1 _11745_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17252_ _17908_/CLK _17252_/D vssd1 vssd1 vccd1 vccd1 _17252_/Q sky130_fd_sc_hd__dfxtp_1
X_14464_ hold1027/X _14481_/B _14463_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14464_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11676_ _12243_/A _11676_/B vssd1 vssd1 vccd1 vccd1 _11676_/X sky130_fd_sc_hd__or2_1
XFILLER_0_71_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16203_ _17435_/CLK _16203_/D vssd1 vssd1 vccd1 vccd1 _16203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13415_ hold1594/X hold4963/X _13817_/C vssd1 vssd1 vccd1 vccd1 _13416_/B sky130_fd_sc_hd__mux2_1
X_10627_ _10651_/A _10627_/B vssd1 vssd1 vccd1 vccd1 _10627_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_10_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17183_ _17247_/CLK _17183_/D vssd1 vssd1 vccd1 vccd1 _17183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14395_ _14395_/A _14443_/B vssd1 vssd1 vccd1 vccd1 _14395_/X sky130_fd_sc_hd__or2_1
XFILLER_0_141_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16134_ _17309_/CLK _16134_/D vssd1 vssd1 vccd1 vccd1 hold303/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13346_ hold2367/X hold4230/X _13862_/C vssd1 vssd1 vccd1 vccd1 _13347_/B sky130_fd_sc_hd__mux2_1
X_10558_ hold5163/X _10070_/B _10557_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10558_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16065_ _17320_/CLK _16065_/D vssd1 vssd1 vccd1 vccd1 hold531/A sky130_fd_sc_hd__dfxtp_1
X_13277_ _13276_/X hold3473/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13277_/X sky130_fd_sc_hd__mux2_1
X_10489_ hold4007/X _10619_/B _10488_/X _14853_/C1 vssd1 vssd1 vccd1 vccd1 _10489_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15016_ hold289/A hold510/A vssd1 vssd1 vccd1 vccd1 hold200/A sky130_fd_sc_hd__or2_1
X_12228_ _13482_/A _12228_/B vssd1 vssd1 vccd1 vccd1 _12228_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12159_ _12159_/A _12159_/B vssd1 vssd1 vccd1 vccd1 _12159_/X sky130_fd_sc_hd__or2_1
XFILLER_0_75_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_236_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1809 _17802_/Q vssd1 vssd1 vccd1 vccd1 hold1809/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16967_ _17847_/CLK _16967_/D vssd1 vssd1 vccd1 vccd1 _16967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15918_ _17293_/CLK _15918_/D vssd1 vssd1 vccd1 vccd1 hold473/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16898_ _18064_/CLK _16898_/D vssd1 vssd1 vccd1 vccd1 _16898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15849_ _17734_/CLK _15849_/D vssd1 vssd1 vccd1 vccd1 _15849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_266_wb_clk_i clkbuf_6_56_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18222_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09370_ hold585/X _09367_/A _09392_/C hold803/X vssd1 vssd1 vccd1 vccd1 _09370_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08321_ _15545_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08321_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17519_ _17520_/CLK hold939/X vssd1 vssd1 vccd1 vccd1 _17519_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_157_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08252_ _15531_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08252_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08183_ _14457_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08183_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5103 _16946_/Q vssd1 vssd1 vccd1 vccd1 hold5103/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5114 _11563_/X vssd1 vssd1 vccd1 vccd1 _17011_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5125 _17258_/Q vssd1 vssd1 vccd1 vccd1 hold5125/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5136 _11656_/X vssd1 vssd1 vccd1 vccd1 _17042_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4402 _17573_/Q vssd1 vssd1 vccd1 vccd1 hold4402/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5147 _10096_/X vssd1 vssd1 vccd1 vccd1 _16522_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5158 _10891_/X vssd1 vssd1 vccd1 vccd1 _16787_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4413 _11797_/Y vssd1 vssd1 vccd1 vccd1 _17089_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4424 _17585_/Q vssd1 vssd1 vccd1 vccd1 hold4424/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5169 _17719_/Q vssd1 vssd1 vccd1 vccd1 hold5169/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4435 _12337_/Y vssd1 vssd1 vccd1 vccd1 _17269_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3701 _10147_/X vssd1 vssd1 vccd1 vccd1 _16539_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4446 _12929_/X vssd1 vssd1 vccd1 vccd1 _12930_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3712 _16603_/Q vssd1 vssd1 vccd1 vccd1 hold3712/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4457 _10246_/X vssd1 vssd1 vccd1 vccd1 _16572_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4468 _12941_/X vssd1 vssd1 vccd1 vccd1 _12942_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3723 _12707_/X vssd1 vssd1 vccd1 vccd1 _12708_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3734 _16399_/Q vssd1 vssd1 vccd1 vccd1 hold3734/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4479 _17504_/Q vssd1 vssd1 vccd1 vccd1 hold4479/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3745 _09778_/X vssd1 vssd1 vccd1 vccd1 _16416_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3756 _09754_/X vssd1 vssd1 vccd1 vccd1 _16408_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3767 _17430_/Q vssd1 vssd1 vccd1 vccd1 hold3767/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3778 _09703_/X vssd1 vssd1 vccd1 vccd1 _16391_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3789 _11784_/Y vssd1 vssd1 vccd1 vccd1 _11785_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07967_ hold2068/X _07978_/B _07966_/X _08167_/A vssd1 vssd1 vccd1 vccd1 _07967_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_226_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09706_ hold4775/X _09992_/B _09705_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _09706_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07898_ _15521_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07898_/X sky130_fd_sc_hd__or2_1
X_09637_ hold4656/X _10028_/B _09636_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09637_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09568_ hold3678/X _10046_/B _09567_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09568_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08519_ _17523_/Q _17522_/Q vssd1 vssd1 vccd1 vccd1 _13057_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_33_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09499_ _18461_/Q _12510_/B vssd1 vssd1 vccd1 vccd1 _09499_/Y sky130_fd_sc_hd__nand2_8
XFILLER_0_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11530_ hold4179/X _12299_/B _11529_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _11530_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_1333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11461_ hold5127/X _11165_/B _11460_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _11461_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ _13193_/X _13199_/X _13296_/B1 vssd1 vssd1 vccd1 vccd1 _17543_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_163_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10412_ hold1899/X hold3626/X _10604_/C vssd1 vssd1 vccd1 vccd1 _10413_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11392_ hold4020/X _11786_/B _11391_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _11392_/X
+ sky130_fd_sc_hd__o211a_1
X_14180_ _15145_/A _14204_/B vssd1 vssd1 vccd1 vccd1 _14180_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13131_ _13130_/X hold4636/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13131_/X sky130_fd_sc_hd__mux2_1
X_10343_ hold2485/X hold3814/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10344_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5670 _11431_/X vssd1 vssd1 vccd1 vccd1 _16967_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10274_ hold1209/X _16582_/Q _10625_/C vssd1 vssd1 vccd1 vccd1 _10275_/B sky130_fd_sc_hd__mux2_1
X_13062_ _13062_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13062_/X sky130_fd_sc_hd__or2_1
Xhold5681 _17225_/Q vssd1 vssd1 vccd1 vccd1 hold5681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5692 _11242_/X vssd1 vssd1 vccd1 vccd1 _16904_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12013_ hold5687/X _12299_/B _12012_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _12013_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_218_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4980 _10894_/X vssd1 vssd1 vccd1 vccd1 _16788_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17870_ _17902_/CLK hold522/X vssd1 vssd1 vccd1 vccd1 _17870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4991 _16858_/Q vssd1 vssd1 vccd1 vccd1 hold4991/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16821_ _18024_/CLK _16821_/D vssd1 vssd1 vccd1 vccd1 _16821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout480 _11774_/C vssd1 vssd1 vccd1 vccd1 _12335_/C sky130_fd_sc_hd__clkbuf_8
Xfanout491 _11201_/C vssd1 vssd1 vccd1 vccd1 _09992_/C sky130_fd_sc_hd__buf_6
XFILLER_0_79_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16752_ _18051_/CLK _16752_/D vssd1 vssd1 vccd1 vccd1 _16752_/Q sky130_fd_sc_hd__dfxtp_1
X_13964_ _15525_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13964_/X sky130_fd_sc_hd__or2_1
XFILLER_0_205_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_232_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15703_ _17281_/CLK _15703_/D vssd1 vssd1 vccd1 vccd1 _15703_/Q sky130_fd_sc_hd__dfxtp_1
X_12915_ _12924_/A _12915_/B vssd1 vssd1 vccd1 vccd1 _17481_/D sky130_fd_sc_hd__and2_1
X_16683_ _18081_/CLK _16683_/D vssd1 vssd1 vccd1 vccd1 _16683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13895_ _13895_/A _13895_/B vssd1 vssd1 vccd1 vccd1 _17755_/D sky130_fd_sc_hd__and2_1
XFILLER_0_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18422_ _18424_/CLK _18422_/D vssd1 vssd1 vccd1 vccd1 _18422_/Q sky130_fd_sc_hd__dfxtp_1
X_15634_ _17900_/CLK _15634_/D vssd1 vssd1 vccd1 vccd1 _15634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12846_ _12849_/A _12846_/B vssd1 vssd1 vccd1 vccd1 _17458_/D sky130_fd_sc_hd__and2_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18353_ _18385_/CLK _18353_/D vssd1 vssd1 vccd1 vccd1 _18353_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _17266_/CLK _15565_/D vssd1 vssd1 vccd1 vccd1 _15565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12777_ _12777_/A _12777_/B vssd1 vssd1 vccd1 vccd1 _17435_/D sky130_fd_sc_hd__and2_1
XFILLER_0_68_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _17322_/CLK _17304_/D vssd1 vssd1 vccd1 vccd1 hold349/A sky130_fd_sc_hd__dfxtp_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14516_ hold3019/X _14537_/B _14515_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _14516_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18284_ _18342_/CLK _18284_/D vssd1 vssd1 vccd1 vccd1 _18284_/Q sky130_fd_sc_hd__dfxtp_1
X_11728_ _12301_/A _11728_/B vssd1 vssd1 vccd1 vccd1 _17066_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_232_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15496_ _15498_/A _15496_/B vssd1 vssd1 vccd1 vccd1 _18427_/D sky130_fd_sc_hd__and2_1
XFILLER_0_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17235_ _17897_/CLK _17235_/D vssd1 vssd1 vccd1 vccd1 _17235_/Q sky130_fd_sc_hd__dfxtp_1
X_14447_ _15128_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14447_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_181_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11659_ hold5667/X _11753_/B _11658_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11659_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17166_ _17868_/CLK _17166_/D vssd1 vssd1 vccd1 vccd1 _17166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14378_ _14380_/A hold151/X vssd1 vssd1 vccd1 vccd1 hold152/A sky130_fd_sc_hd__and2_1
XFILLER_0_12_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold906 hold906/A vssd1 vssd1 vccd1 vccd1 hold906/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16117_ _17344_/CLK _16117_/D vssd1 vssd1 vccd1 vccd1 hold264/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold917 hold917/A vssd1 vssd1 vccd1 vccd1 hold917/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold928 hold928/A vssd1 vssd1 vccd1 vccd1 hold928/X sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ _13719_/A _13329_/B vssd1 vssd1 vccd1 vccd1 _13329_/X sky130_fd_sc_hd__or2_1
Xhold939 hold939/A vssd1 vssd1 vccd1 vccd1 hold939/X sky130_fd_sc_hd__dlygate4sd3_1
X_17097_ _17161_/CLK _17097_/D vssd1 vssd1 vccd1 vccd1 _17097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_228_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16048_ _16124_/CLK _16048_/D vssd1 vssd1 vccd1 vccd1 hold261/A sky130_fd_sc_hd__dfxtp_1
Xhold3008 _18331_/Q vssd1 vssd1 vccd1 vccd1 hold3008/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3019 _18054_/Q vssd1 vssd1 vccd1 vccd1 hold3019/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2307 _15222_/X vssd1 vssd1 vccd1 vccd1 _18393_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08870_ hold226/X hold647/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold648/A sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2318 _15578_/Q vssd1 vssd1 vccd1 vccd1 hold2318/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2329 _14458_/X vssd1 vssd1 vccd1 vccd1 _18026_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07821_ _15555_/A hold992/A _15553_/A vssd1 vssd1 vccd1 vccd1 _07824_/C sky130_fd_sc_hd__or3b_1
Xhold1606 _17979_/Q vssd1 vssd1 vccd1 vccd1 hold1606/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1617 _14528_/X vssd1 vssd1 vccd1 vccd1 _18060_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1628 _17782_/Q vssd1 vssd1 vccd1 vccd1 hold1628/X sky130_fd_sc_hd__dlygate4sd3_1
X_17999_ _18054_/CLK _17999_/D vssd1 vssd1 vccd1 vccd1 _17999_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1639 _16174_/Q vssd1 vssd1 vccd1 vccd1 hold1639/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_447_wb_clk_i clkbuf_6_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17628_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_193_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09422_ _09438_/B _16297_/Q vssd1 vssd1 vccd1 vccd1 _09422_/X sky130_fd_sc_hd__or2_1
XFILLER_0_176_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09353_ _15547_/A hold220/A _09359_/C vssd1 vssd1 vccd1 vccd1 _09361_/C sky130_fd_sc_hd__or3_1
XFILLER_0_34_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08304_ hold2897/X _08336_/A2 _08303_/X _08347_/A vssd1 vssd1 vccd1 vccd1 _08304_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09284_ _12777_/A _09284_/B vssd1 vssd1 vccd1 vccd1 _16253_/D sky130_fd_sc_hd__and2_1
XFILLER_0_47_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08235_ hold1935/X _08262_/B _08234_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _08235_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08166_ _15517_/A hold2375/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08167_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08097_ hold1279/X _08097_/A2 _08096_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _08097_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4210 _15253_/X vssd1 vssd1 vccd1 vccd1 _15254_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4221 hold5913/X vssd1 vssd1 vccd1 vccd1 hold5914/A sky130_fd_sc_hd__buf_4
Xhold4232 _13828_/Y vssd1 vssd1 vccd1 vccd1 _17729_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4243 _13821_/Y vssd1 vssd1 vccd1 vccd1 _13822_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4254 _16337_/Q vssd1 vssd1 vccd1 vccd1 _13166_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4265 _10032_/Y vssd1 vssd1 vccd1 vccd1 _10033_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3520 _16911_/Q vssd1 vssd1 vccd1 vccd1 hold3520/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4276 _16328_/Q vssd1 vssd1 vccd1 vccd1 _13094_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3531 _12776_/X vssd1 vssd1 vccd1 vccd1 _12777_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3542 _09967_/X vssd1 vssd1 vccd1 vccd1 _16479_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4287 hold4978/X vssd1 vssd1 vccd1 vccd1 _13832_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3553 _09583_/X vssd1 vssd1 vccd1 vccd1 _16351_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4298 _17104_/Q vssd1 vssd1 vccd1 vccd1 hold4298/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3564 _16363_/Q vssd1 vssd1 vccd1 vccd1 hold3564/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3575 _09817_/X vssd1 vssd1 vccd1 vccd1 _16429_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2830 _16165_/Q vssd1 vssd1 vccd1 vccd1 hold2830/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3586 _16395_/Q vssd1 vssd1 vccd1 vccd1 hold3586/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2841 _07905_/X vssd1 vssd1 vccd1 vccd1 _15596_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2852 _18390_/Q vssd1 vssd1 vccd1 vccd1 hold2852/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08999_ _13046_/C _12445_/B vssd1 vssd1 vccd1 vccd1 _09062_/S sky130_fd_sc_hd__or2_2
Xhold3597 _16515_/Q vssd1 vssd1 vccd1 vccd1 hold3597/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2863 _18435_/Q vssd1 vssd1 vccd1 vccd1 hold2863/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_188_wb_clk_i clkbuf_6_52_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18323_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_138_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2874 _14015_/X vssd1 vssd1 vccd1 vccd1 _17813_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2885 _14063_/X vssd1 vssd1 vccd1 vccd1 _17836_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2896 _08483_/X vssd1 vssd1 vccd1 vccd1 _15870_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_117_wb_clk_i clkbuf_6_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17525_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_173_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10961_ hold2629/X hold4972/X _11153_/C vssd1 vssd1 vccd1 vccd1 _10962_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_211_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12700_ hold2524/X _17411_/Q _12766_/S vssd1 vssd1 vccd1 vccd1 _12700_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13680_ _13776_/A _13680_/B vssd1 vssd1 vccd1 vccd1 _13680_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10892_ hold1955/X _16788_/Q _11186_/C vssd1 vssd1 vccd1 vccd1 _10893_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_210_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12631_ hold2683/X _17388_/Q _12850_/S vssd1 vssd1 vccd1 vccd1 _12631_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15350_ hold872/X _09367_/A _09392_/A hold730/X vssd1 vssd1 vccd1 vccd1 _15350_/X
+ sky130_fd_sc_hd__a22o_1
X_12562_ hold1990/X hold3636/X _12925_/S vssd1 vssd1 vccd1 vccd1 _12562_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_65_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14301_ hold2908/X _14333_/A2 _14300_/X _14552_/C1 vssd1 vssd1 vccd1 vccd1 _14301_/X
+ sky130_fd_sc_hd__o211a_1
X_11513_ hold1873/X _16995_/Q _11774_/C vssd1 vssd1 vccd1 vccd1 _11514_/B sky130_fd_sc_hd__mux2_1
X_15281_ _09412_/B _15477_/A2 _15487_/B1 hold468/X _15280_/X vssd1 vssd1 vccd1 vccd1
+ _15282_/D sky130_fd_sc_hd__a221o_1
X_12493_ hold92/A _12509_/A2 _12501_/A3 _12492_/X _12440_/A vssd1 vssd1 vccd1 vccd1
+ hold66/A sky130_fd_sc_hd__o311a_1
XFILLER_0_149_1250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17020_ _17868_/CLK _17020_/D vssd1 vssd1 vccd1 vccd1 _17020_/Q sky130_fd_sc_hd__dfxtp_1
X_14232_ hold406/X _14502_/B vssd1 vssd1 vccd1 vccd1 _14232_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_145_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11444_ hold2062/X _16972_/Q _11732_/C vssd1 vssd1 vccd1 vccd1 _11445_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14163_ hold330/X _14163_/B vssd1 vssd1 vccd1 vccd1 _14204_/B sky130_fd_sc_hd__or2_4
XFILLER_0_225_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11375_ hold2798/X hold4961/X _11765_/C vssd1 vssd1 vccd1 vccd1 _11376_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13114_ _17565_/Q _17099_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13114_/X sky130_fd_sc_hd__mux2_1
X_10326_ _10542_/A _10326_/B vssd1 vssd1 vccd1 vccd1 _10326_/X sky130_fd_sc_hd__or2_1
X_14094_ _15547_/A _14094_/B vssd1 vssd1 vccd1 vccd1 _14094_/Y sky130_fd_sc_hd__nand2_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _17524_/Q hold923/X _13044_/X _13056_/C _13048_/A vssd1 vssd1 vccd1 vccd1
+ hold924/A sky130_fd_sc_hd__o221a_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _18019_/CLK _17922_/D vssd1 vssd1 vccd1 vccd1 _17922_/Q sky130_fd_sc_hd__dfxtp_1
X_10257_ _10551_/A _10257_/B vssd1 vssd1 vccd1 vccd1 _10257_/X sky130_fd_sc_hd__or2_1
X_10188_ _10560_/A _10188_/B vssd1 vssd1 vccd1 vccd1 _10188_/X sky130_fd_sc_hd__or2_1
X_17853_ _17853_/CLK _17853_/D vssd1 vssd1 vccd1 vccd1 _17853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_233_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16804_ _18039_/CLK _16804_/D vssd1 vssd1 vccd1 vccd1 _16804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14996_ _15103_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14996_/X sky130_fd_sc_hd__or2_1
X_17784_ _17846_/CLK _17784_/D vssd1 vssd1 vccd1 vccd1 _17784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_233_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16735_ _18194_/CLK _16735_/D vssd1 vssd1 vccd1 vccd1 _16735_/Q sky130_fd_sc_hd__dfxtp_1
X_13947_ _14627_/A _14163_/B vssd1 vssd1 vccd1 vccd1 _13994_/B sky130_fd_sc_hd__or2_4
XFILLER_0_205_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16666_ _18224_/CLK _16666_/D vssd1 vssd1 vccd1 vccd1 _16666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13878_ hold3547/X _13791_/A _13877_/X vssd1 vssd1 vccd1 vccd1 _13878_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18405_ _18405_/CLK _18405_/D vssd1 vssd1 vccd1 vccd1 _18405_/Q sky130_fd_sc_hd__dfxtp_1
X_15617_ _17236_/CLK _15617_/D vssd1 vssd1 vccd1 vccd1 _15617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12829_ hold1923/X _17454_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12829_/X sky130_fd_sc_hd__mux2_1
X_16597_ _18233_/CLK _16597_/D vssd1 vssd1 vccd1 vccd1 _16597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_227_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18336_ _18398_/CLK _18336_/D vssd1 vssd1 vccd1 vccd1 _18336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15548_ hold2437/X _15547_/B _15547_/Y _12873_/A vssd1 vssd1 vccd1 vccd1 _15548_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18267_ _18391_/CLK _18267_/D vssd1 vssd1 vccd1 vccd1 _18267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15479_ _17323_/Q _09357_/A _09362_/C hold827/X _15478_/X vssd1 vssd1 vccd1 vccd1
+ _15480_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_142_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08020_ hold2396/X _08029_/B _08019_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _08020_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17218_ _17250_/CLK _17218_/D vssd1 vssd1 vccd1 vccd1 _17218_/Q sky130_fd_sc_hd__dfxtp_1
X_18198_ _18231_/CLK _18198_/D vssd1 vssd1 vccd1 vccd1 _18198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold703 hold711/X vssd1 vssd1 vccd1 vccd1 hold712/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold714 hold714/A vssd1 vssd1 vccd1 vccd1 hold714/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17149_ _17236_/CLK _17149_/D vssd1 vssd1 vccd1 vccd1 _17149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold725 hold725/A vssd1 vssd1 vccd1 vccd1 hold725/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold736 hold736/A vssd1 vssd1 vccd1 vccd1 hold736/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 hold747/A vssd1 vssd1 vccd1 vccd1 hold747/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 hold758/A vssd1 vssd1 vccd1 vccd1 hold758/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09971_ _18394_/Q hold3266/X _10475_/S vssd1 vssd1 vccd1 vccd1 _09972_/B sky130_fd_sc_hd__mux2_1
Xhold769 hold769/A vssd1 vssd1 vccd1 vccd1 hold769/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08922_ hold315/X hold782/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08923_/B sky130_fd_sc_hd__mux2_1
Xhold2104 hold2104/A vssd1 vssd1 vccd1 vccd1 _15145_/A sky130_fd_sc_hd__buf_12
Xhold2115 _18094_/Q vssd1 vssd1 vccd1 vccd1 hold2115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2126 _14225_/X vssd1 vssd1 vccd1 vccd1 _17914_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2137 _18324_/Q vssd1 vssd1 vccd1 vccd1 hold2137/X sky130_fd_sc_hd__dlygate4sd3_1
X_08853_ _12416_/A _08853_/B vssd1 vssd1 vccd1 vccd1 _16045_/D sky130_fd_sc_hd__and2_1
XFILLER_0_224_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1403 _14277_/X vssd1 vssd1 vccd1 vccd1 _17939_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2148 _14099_/X vssd1 vssd1 vccd1 vccd1 _17854_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1414 _18440_/Q vssd1 vssd1 vccd1 vccd1 hold1414/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2159 _16269_/Q vssd1 vssd1 vccd1 vccd1 hold2159/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1425 _15742_/Q vssd1 vssd1 vccd1 vccd1 hold1425/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07804_ _07804_/A _16286_/Q vssd1 vssd1 vccd1 vccd1 _07805_/A sky130_fd_sc_hd__and2_4
Xclkbuf_leaf_281_wb_clk_i clkbuf_6_50_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18023_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1436 _15849_/Q vssd1 vssd1 vccd1 vccd1 hold1436/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 _09091_/X vssd1 vssd1 vccd1 vccd1 _16160_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08784_ _15473_/A hold316/X vssd1 vssd1 vccd1 vccd1 _16012_/D sky130_fd_sc_hd__and2_1
Xhold1458 _13995_/X vssd1 vssd1 vccd1 vccd1 _17804_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_240_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1469 _09123_/X vssd1 vssd1 vccd1 vccd1 _16175_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_210_wb_clk_i clkbuf_6_54_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18298_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09405_ _07804_/A hold5994/X _15284_/A _09404_/X vssd1 vssd1 vccd1 vccd1 _09405_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09336_ hold1309/X _09325_/B _09335_/X _12612_/A vssd1 vssd1 vccd1 vccd1 _09336_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09267_ hold597/X _16245_/Q hold271/X vssd1 vssd1 vccd1 vccd1 hold598/A sky130_fd_sc_hd__mux2_1
XFILLER_0_161_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08218_ hold1489/X _08213_/B _08217_/X _08347_/A vssd1 vssd1 vccd1 vccd1 _08218_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09198_ hold951/X _09206_/B vssd1 vssd1 vccd1 vccd1 _09198_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08149_ _08149_/A _08149_/B vssd1 vssd1 vccd1 vccd1 _15713_/D sky130_fd_sc_hd__and2_1
XFILLER_0_160_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11160_ hold4281/X _11067_/A _11159_/X vssd1 vssd1 vccd1 vccd1 _11160_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4040 _17040_/Q vssd1 vssd1 vccd1 vccd1 hold4040/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10111_ hold3834/X _10589_/B _10110_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10111_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4051 _11422_/X vssd1 vssd1 vccd1 vccd1 _16964_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11091_ _11091_/A _11091_/B vssd1 vssd1 vccd1 vccd1 _11091_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_369_wb_clk_i clkbuf_6_34_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17733_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4062 _12028_/X vssd1 vssd1 vccd1 vccd1 _17166_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4073 _11893_/X vssd1 vssd1 vccd1 vccd1 _17121_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4084 _11521_/X vssd1 vssd1 vccd1 vccd1 _16997_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4095 _16776_/Q vssd1 vssd1 vccd1 vccd1 hold4095/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3350 _17443_/Q vssd1 vssd1 vccd1 vccd1 hold3350/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ _11206_/A _10042_/B vssd1 vssd1 vccd1 vccd1 _16504_/D sky130_fd_sc_hd__nor2_1
Xhold3361 _17469_/Q vssd1 vssd1 vccd1 vccd1 hold3361/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3372 _17405_/Q vssd1 vssd1 vccd1 vccd1 hold3372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3383 _17407_/Q vssd1 vssd1 vccd1 vccd1 hold3383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__buf_4
XFILLER_0_215_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3394 _17428_/Q vssd1 vssd1 vccd1 vccd1 hold3394/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2660 _14703_/X vssd1 vssd1 vccd1 vccd1 _18143_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14850_ _14850_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14850_/X sky130_fd_sc_hd__or2_1
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2671 _15746_/Q vssd1 vssd1 vccd1 vccd1 hold2671/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__buf_1
Xhold2682 _14649_/X vssd1 vssd1 vccd1 vccd1 _18117_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold85 hold7/X vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2693 _18038_/Q vssd1 vssd1 vccd1 vccd1 hold2693/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ hold5006/X _13814_/B _13800_/X _13801_/C1 vssd1 vssd1 vccd1 vccd1 _13801_/X
+ sky130_fd_sc_hd__o211a_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1970 _17807_/Q vssd1 vssd1 vccd1 vccd1 hold1970/X sky130_fd_sc_hd__dlygate4sd3_1
X_14781_ hold2906/X _14772_/B _14780_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14781_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1981 _14867_/X vssd1 vssd1 vccd1 vccd1 _18222_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1992 _16295_/Q vssd1 vssd1 vccd1 vccd1 _09418_/B sky130_fd_sc_hd__dlygate4sd3_1
X_11993_ hold2449/X _17155_/Q _13886_/C vssd1 vssd1 vccd1 vccd1 _11994_/B sky130_fd_sc_hd__mux2_1
X_16520_ _18265_/CLK _16520_/D vssd1 vssd1 vccd1 vccd1 _16520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13732_ hold4733/X _13862_/B _13731_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _13732_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10944_ _11136_/A _10944_/B vssd1 vssd1 vccd1 vccd1 _10944_/X sky130_fd_sc_hd__or2_1
XFILLER_0_211_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16451_ _18396_/CLK _16451_/D vssd1 vssd1 vccd1 vccd1 _16451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13663_ hold5498/X _13874_/B _13662_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13663_/X
+ sky130_fd_sc_hd__o211a_1
X_10875_ _11067_/A _10875_/B vssd1 vssd1 vccd1 vccd1 _10875_/X sky130_fd_sc_hd__or2_1
XFILLER_0_210_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15402_ _15480_/A _15402_/B _15402_/C _15402_/D vssd1 vssd1 vccd1 vccd1 _15402_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_151_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ hold3385/X _12613_/X _12923_/S vssd1 vssd1 vccd1 vccd1 _12614_/X sky130_fd_sc_hd__mux2_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16382_ _18389_/CLK _16382_/D vssd1 vssd1 vccd1 vccd1 _16382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13594_ hold5337/X _13883_/B _13593_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13594_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18121_ _18177_/CLK _18121_/D vssd1 vssd1 vccd1 vccd1 _18121_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_85_wb_clk_i clkbuf_6_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17506_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_137_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15333_ _15490_/A1 _15325_/X _15332_/X _15490_/B1 hold5946/A vssd1 vssd1 vccd1 vccd1
+ _15333_/X sky130_fd_sc_hd__a32o_1
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12545_ hold4534/X _12544_/X _12929_/S vssd1 vssd1 vccd1 vccd1 _12546_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_14_wb_clk_i clkbuf_6_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18451_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18052_ _18052_/CLK _18052_/D vssd1 vssd1 vccd1 vccd1 _18052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15264_ _15414_/A _15264_/B vssd1 vssd1 vccd1 vccd1 _18402_/D sky130_fd_sc_hd__and2_1
X_12476_ _17331_/Q _12506_/B vssd1 vssd1 vccd1 vccd1 _12476_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17003_ _17883_/CLK _17003_/D vssd1 vssd1 vccd1 vccd1 _17003_/Q sky130_fd_sc_hd__dfxtp_1
X_14215_ hold1525/X _14198_/B _14214_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _14215_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_5 _13068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11427_ _11622_/A _11427_/B vssd1 vssd1 vccd1 vccd1 _11427_/X sky130_fd_sc_hd__or2_1
X_15195_ _15195_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15195_/X sky130_fd_sc_hd__or2_1
XFILLER_0_223_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14146_ _15545_/A _14148_/B vssd1 vssd1 vccd1 vccd1 _14146_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11358_ _11553_/A _11358_/B vssd1 vssd1 vccd1 vccd1 _11358_/X sky130_fd_sc_hd__or2_1
X_10309_ hold3757/X _10631_/B _10308_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10309_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14077_ hold1873/X _14107_/A2 _14076_/X _14143_/C1 vssd1 vssd1 vccd1 vccd1 _14077_/X
+ sky130_fd_sc_hd__o211a_1
X_11289_ _11694_/A _11289_/B vssd1 vssd1 vccd1 vccd1 _11289_/X sky130_fd_sc_hd__or2_1
XFILLER_0_197_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13028_ _13029_/B hold905/X hold938/X vssd1 vssd1 vccd1 vccd1 hold939/A sky130_fd_sc_hd__and3b_1
X_17905_ _17905_/CLK _17905_/D vssd1 vssd1 vccd1 vccd1 _17905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17836_ _17887_/CLK _17836_/D vssd1 vssd1 vccd1 vccd1 _17836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17767_ _17799_/CLK _17767_/D vssd1 vssd1 vccd1 vccd1 _17767_/Q sky130_fd_sc_hd__dfxtp_1
X_14979_ hold6076/X hold447/X _14978_/X _15044_/A vssd1 vssd1 vccd1 vccd1 hold448/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_234_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16718_ _18049_/CLK _16718_/D vssd1 vssd1 vccd1 vccd1 _16718_/Q sky130_fd_sc_hd__dfxtp_1
X_17698_ _17730_/CLK _17698_/D vssd1 vssd1 vccd1 vccd1 _17698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16649_ _18235_/CLK _16649_/D vssd1 vssd1 vccd1 vccd1 _16649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09121_ _15555_/A _09121_/B _15553_/A hold992/A vssd1 vssd1 vccd1 vccd1 _09400_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_84_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18319_ _18385_/CLK _18319_/D vssd1 vssd1 vccd1 vccd1 _18319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09052_ hold315/X hold864/X _09060_/S vssd1 vssd1 vccd1 vccd1 _09053_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_163_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08003_ _14457_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08003_/X sky130_fd_sc_hd__or2_1
Xhold500 hold500/A vssd1 vssd1 vccd1 vccd1 hold500/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 hold511/A vssd1 vssd1 vccd1 vccd1 hold511/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 hold522/A vssd1 vssd1 vccd1 vccd1 hold522/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold533 hold533/A vssd1 vssd1 vccd1 vccd1 hold533/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold544 hold544/A vssd1 vssd1 vccd1 vccd1 hold544/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold555 hold555/A vssd1 vssd1 vccd1 vccd1 hold555/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold566 hold566/A vssd1 vssd1 vccd1 vccd1 hold566/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 hold577/A vssd1 vssd1 vccd1 vccd1 input54/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold588 hold588/A vssd1 vssd1 vccd1 vccd1 hold588/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_462_wb_clk_i clkbuf_6_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17434_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09954_ _09954_/A _09954_/B vssd1 vssd1 vccd1 vccd1 _09954_/X sky130_fd_sc_hd__or2_1
XFILLER_0_99_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold599 hold599/A vssd1 vssd1 vccd1 vccd1 hold599/X sky130_fd_sc_hd__dlygate4sd3_1
X_08905_ _12416_/A _08905_/B vssd1 vssd1 vccd1 vccd1 _16070_/D sky130_fd_sc_hd__and2_1
XFILLER_0_176_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09885_ _09981_/A _09885_/B vssd1 vssd1 vccd1 vccd1 _09885_/X sky130_fd_sc_hd__or2_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1200 _15204_/X vssd1 vssd1 vccd1 vccd1 _18384_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1211 _18256_/Q vssd1 vssd1 vccd1 vccd1 hold1211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ hold185/X hold661/X _08860_/S vssd1 vssd1 vccd1 vccd1 hold662/A sky130_fd_sc_hd__mux2_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1222 la_data_in[22] vssd1 vssd1 vccd1 vccd1 hold1222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1233 _17838_/Q vssd1 vssd1 vccd1 vccd1 hold1233/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_225_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1244 _18216_/Q vssd1 vssd1 vccd1 vccd1 hold1244/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1255 _08134_/X vssd1 vssd1 vccd1 vccd1 _08135_/B sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_6_15_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_15_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1266 _14805_/X vssd1 vssd1 vccd1 vccd1 _18192_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08767_ hold245/X hold478/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08768_/B sky130_fd_sc_hd__mux2_1
Xhold1277 _15670_/Q vssd1 vssd1 vccd1 vccd1 hold1277/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1288 _08087_/X vssd1 vssd1 vccd1 vccd1 _15683_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_234_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1299 _18267_/Q vssd1 vssd1 vccd1 vccd1 hold1299/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ _15374_/A hold206/X vssd1 vssd1 vccd1 vccd1 _15970_/D sky130_fd_sc_hd__and2_1
XFILLER_0_67_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10660_ hold5541/X _11732_/B _10659_/X _13895_/A vssd1 vssd1 vccd1 vccd1 _10660_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09319_ _15541_/A _09323_/B vssd1 vssd1 vccd1 vccd1 _09319_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_106_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10591_ _10651_/A _10591_/B vssd1 vssd1 vccd1 vccd1 _16687_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_69_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12330_ hold4722/X _12234_/A _12329_/X vssd1 vssd1 vccd1 vccd1 _12330_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12261_ _13482_/A _12261_/B vssd1 vssd1 vccd1 vccd1 _12261_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14000_ _14681_/A _14163_/B vssd1 vssd1 vccd1 vccd1 _14000_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_181_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11212_ _12331_/A _11212_/B vssd1 vssd1 vccd1 vccd1 _11212_/Y sky130_fd_sc_hd__nor2_1
X_12192_ _13314_/A _12192_/B vssd1 vssd1 vccd1 vccd1 _12192_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_6_54_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_54_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_6010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11143_ _11158_/A _11143_/B vssd1 vssd1 vccd1 vccd1 _11143_/Y sky130_fd_sc_hd__nor2_1
XTAP_6021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput75 _13153_/A vssd1 vssd1 vccd1 vccd1 output75/X sky130_fd_sc_hd__buf_6
Xoutput86 _13233_/A vssd1 vssd1 vccd1 vccd1 output86/X sky130_fd_sc_hd__buf_6
XFILLER_0_235_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_132_wb_clk_i clkbuf_6_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17303_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xoutput97 _13081_/A vssd1 vssd1 vccd1 vccd1 output97/X sky130_fd_sc_hd__buf_6
XTAP_6054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15951_ _17319_/CLK _15951_/D vssd1 vssd1 vccd1 vccd1 hold668/A sky130_fd_sc_hd__dfxtp_1
XTAP_5320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11074_ hold5488/X _11744_/B _11073_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _11074_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3180 _17921_/Q vssd1 vssd1 vccd1 vccd1 hold3180/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10025_ _16499_/Q _10025_/B _10025_/C vssd1 vssd1 vccd1 vccd1 _10025_/X sky130_fd_sc_hd__and3_1
XTAP_6098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14902_ _14972_/A _14910_/B vssd1 vssd1 vccd1 vccd1 _14902_/X sky130_fd_sc_hd__or2_1
Xhold3191 _17973_/Q vssd1 vssd1 vccd1 vccd1 hold3191/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15882_ _17561_/CLK _15882_/D vssd1 vssd1 vccd1 vccd1 _15882_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2490 _14101_/X vssd1 vssd1 vccd1 vccd1 _17855_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ _17653_/CLK _17621_/D vssd1 vssd1 vccd1 vccd1 _17621_/Q sky130_fd_sc_hd__dfxtp_1
X_14833_ hold2096/X _14826_/B _14832_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _14833_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ _18191_/CLK _17552_/D vssd1 vssd1 vccd1 vccd1 _17552_/Q sky130_fd_sc_hd__dfxtp_1
X_14764_ _15103_/A _14780_/B vssd1 vssd1 vccd1 vccd1 _14764_/X sky130_fd_sc_hd__or2_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _12267_/A _11976_/B vssd1 vssd1 vccd1 vccd1 _11976_/X sky130_fd_sc_hd__or2_1
XFILLER_0_187_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16503_ _18392_/CLK _16503_/D vssd1 vssd1 vccd1 vccd1 _16503_/Q sky130_fd_sc_hd__dfxtp_1
X_13715_ hold1568/X hold4756/X _13811_/C vssd1 vssd1 vccd1 vccd1 _13716_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_233_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10927_ hold4063/X _10616_/B _10926_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10927_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17483_ _17484_/CLK _17483_/D vssd1 vssd1 vccd1 vccd1 _17483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14695_ hold2773/X _14718_/B _14694_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14695_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_196_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16434_ _18315_/CLK _16434_/D vssd1 vssd1 vccd1 vccd1 _16434_/Q sky130_fd_sc_hd__dfxtp_1
X_13646_ hold1694/X _17669_/Q _13871_/C vssd1 vssd1 vccd1 vccd1 _13647_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_128_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10858_ hold3724/X _11144_/B _10857_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _10858_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _18382_/CLK _16365_/D vssd1 vssd1 vccd1 vccd1 _16365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13577_ hold2807/X _17646_/Q _13766_/S vssd1 vssd1 vccd1 vccd1 _13578_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_171_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ hold5159/X _11165_/B _10788_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _10789_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15316_ _17335_/Q _15486_/B1 _15485_/B1 _16112_/Q vssd1 vssd1 vccd1 vccd1 _15316_/X
+ sky130_fd_sc_hd__a22o_1
X_18104_ _18156_/CLK _18104_/D vssd1 vssd1 vccd1 vccd1 _18104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12528_ _12984_/A _12528_/B vssd1 vssd1 vccd1 vccd1 _17352_/D sky130_fd_sc_hd__and2_1
XFILLER_0_227_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16296_ _16315_/CLK _16296_/D vssd1 vssd1 vccd1 vccd1 _16296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15247_ hold657/X _15487_/A2 _15484_/B1 hold653/X _15246_/X vssd1 vssd1 vccd1 vccd1
+ _15252_/B sky130_fd_sc_hd__a221o_1
X_18035_ _18058_/CLK _18035_/D vssd1 vssd1 vccd1 vccd1 _18035_/Q sky130_fd_sc_hd__dfxtp_1
X_12459_ hold29/X _08597_/Y _12501_/A3 _12458_/X _15434_/A vssd1 vssd1 vccd1 vccd1
+ hold30/A sky130_fd_sc_hd__o311a_1
XFILLER_0_124_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4809 _17247_/Q vssd1 vssd1 vccd1 vccd1 hold4809/X sky130_fd_sc_hd__dlygate4sd3_1
X_15178_ hold1491/X _15165_/B _15177_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _15178_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14129_ hold2817/X _14148_/B _14128_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _14129_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout309 _09912_/A vssd1 vssd1 vccd1 vccd1 _09948_/A sky130_fd_sc_hd__buf_4
XFILLER_0_120_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09670_ hold3562/X _10052_/B _09669_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09670_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_234_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08621_ hold163/X hold761/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold762/A sky130_fd_sc_hd__mux2_1
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17819_ _18432_/CLK _17819_/D vssd1 vssd1 vccd1 vccd1 _17819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08552_ hold23/X hold411/X _08592_/S vssd1 vssd1 vccd1 vccd1 _08553_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_77_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08483_ hold2895/X _08488_/B _08482_/Y _08139_/A vssd1 vssd1 vccd1 vccd1 _08483_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09104_ _15165_/A _09106_/B vssd1 vssd1 vccd1 vccd1 _09104_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09035_ _15324_/A _09035_/B vssd1 vssd1 vccd1 vccd1 _16134_/D sky130_fd_sc_hd__and2_1
XFILLER_0_131_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold330 hold330/A vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold341 hold341/A vssd1 vssd1 vccd1 vccd1 hold341/X sky130_fd_sc_hd__buf_6
Xhold352 input60/X vssd1 vssd1 vccd1 vccd1 hold352/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_102_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold363 hold363/A vssd1 vssd1 vccd1 vccd1 hold363/X sky130_fd_sc_hd__buf_4
Xhold374 hold374/A vssd1 vssd1 vccd1 vccd1 hold374/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold385 hold385/A vssd1 vssd1 vccd1 vccd1 hold385/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 hold396/A vssd1 vssd1 vccd1 vccd1 hold396/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout810 _15228_/C1 vssd1 vssd1 vccd1 vccd1 _15024_/A sky130_fd_sc_hd__buf_4
XFILLER_0_141_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_217_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout821 _10564_/C1 vssd1 vssd1 vccd1 vccd1 _14841_/C1 sky130_fd_sc_hd__buf_4
X_09937_ hold4754/X _10031_/B _09936_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09937_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout832 _14893_/C1 vssd1 vssd1 vccd1 vccd1 _14807_/C1 sky130_fd_sc_hd__buf_4
Xfanout843 _07787_/Y vssd1 vssd1 vccd1 vccd1 fanout843/X sky130_fd_sc_hd__clkbuf_16
Xfanout854 _11218_/A vssd1 vssd1 vccd1 vccd1 _10603_/A sky130_fd_sc_hd__clkbuf_16
Xfanout865 _07783_/Y vssd1 vssd1 vccd1 vccd1 _15161_/A sky130_fd_sc_hd__clkbuf_16
Xfanout876 hold951/X vssd1 vssd1 vccd1 vccd1 _14413_/A sky130_fd_sc_hd__buf_8
X_09868_ hold3822/X _10052_/B _09867_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _09868_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout887 _15195_/A vssd1 vssd1 vccd1 vccd1 _14980_/A sky130_fd_sc_hd__buf_12
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1030 _14679_/X vssd1 vssd1 vccd1 vccd1 _18132_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout898 _14974_/A vssd1 vssd1 vccd1 vccd1 _14850_/A sky130_fd_sc_hd__buf_12
Xhold1041 _18114_/Q vssd1 vssd1 vccd1 vccd1 hold1041/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08819_ _15244_/A hold838/X vssd1 vssd1 vccd1 vccd1 _16028_/D sky130_fd_sc_hd__and2_1
Xhold1052 _15835_/Q vssd1 vssd1 vccd1 vccd1 hold1052/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1063 _13016_/X vssd1 vssd1 vccd1 vccd1 _17516_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ hold3714/X _10004_/B _09798_/X _08954_/A vssd1 vssd1 vccd1 vccd1 _09799_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1074 hold1145/X vssd1 vssd1 vccd1 vccd1 hold1146/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 _17806_/Q vssd1 vssd1 vccd1 vccd1 hold1085/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1096 _14879_/X vssd1 vssd1 vccd1 vccd1 _18228_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ hold4565/X _13817_/B _11829_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _11830_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _12337_/A _11761_/B vssd1 vssd1 vccd1 vccd1 _11761_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_96_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13500_ _13788_/A _13500_/B vssd1 vssd1 vccd1 vccd1 _13500_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_1303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ hold2094/X hold4531/X _11213_/C vssd1 vssd1 vccd1 vccd1 _10713_/B sky130_fd_sc_hd__mux2_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14480_ hold1799/X _14481_/B _14479_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _14480_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11692_ hold5392/X _12329_/B _11691_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11692_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13431_ _13719_/A _13431_/B vssd1 vssd1 vccd1 vccd1 _13431_/X sky130_fd_sc_hd__or2_1
X_10643_ _16705_/Q _10646_/B _10646_/C vssd1 vssd1 vccd1 vccd1 _10643_/X sky130_fd_sc_hd__and3_1
XFILLER_0_125_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16150_ _17491_/CLK _16150_/D vssd1 vssd1 vccd1 vccd1 _16150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13362_ _13752_/A _13362_/B vssd1 vssd1 vccd1 vccd1 _13362_/X sky130_fd_sc_hd__or2_1
XFILLER_0_51_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10574_ _16682_/Q _11204_/B _11204_/C vssd1 vssd1 vccd1 vccd1 _10574_/X sky130_fd_sc_hd__and3_1
XFILLER_0_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_1350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15101_ hold691/X _15125_/B vssd1 vssd1 vccd1 vccd1 hold692/A sky130_fd_sc_hd__or2_1
XFILLER_0_1_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12313_ _13819_/A _12313_/B vssd1 vssd1 vccd1 vccd1 _17261_/D sky130_fd_sc_hd__nor2_1
X_16081_ _18401_/CLK _16081_/D vssd1 vssd1 vccd1 vccd1 hold516/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_384_wb_clk_i clkbuf_6_33_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17278_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13293_ _13292_/X hold4227/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13293_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15032_ _15054_/A _15032_/B vssd1 vssd1 vccd1 vccd1 _18301_/D sky130_fd_sc_hd__and2_1
X_12244_ _12338_/A _12350_/B _12243_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _12244_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_313_wb_clk_i clkbuf_6_47_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17799_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_210_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12175_ hold4809/X _11798_/B _12174_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _12175_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11126_ hold1951/X hold3958/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11127_/B sky130_fd_sc_hd__mux2_1
X_16983_ _17895_/CLK _16983_/D vssd1 vssd1 vccd1 vccd1 _16983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_236_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_219_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15934_ _17324_/CLK _15934_/D vssd1 vssd1 vccd1 vccd1 hold751/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11057_ hold2127/X _16843_/Q _11153_/C vssd1 vssd1 vccd1 vccd1 _11058_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_200_1280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10008_ _13134_/A _09912_/A _10007_/X vssd1 vssd1 vccd1 vccd1 _10008_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_204_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15865_ _17740_/CLK _15865_/D vssd1 vssd1 vccd1 vccd1 _15865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17604_ _17648_/CLK _17604_/D vssd1 vssd1 vccd1 vccd1 _17604_/Q sky130_fd_sc_hd__dfxtp_1
X_14816_ _15209_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14816_/X sky130_fd_sc_hd__or2_1
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15796_ _17729_/CLK _15796_/D vssd1 vssd1 vccd1 vccd1 _15796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17535_ _17535_/CLK _17535_/D vssd1 vssd1 vccd1 vccd1 _17535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14747_ hold2493/X _14774_/B _14746_/X _14895_/C1 vssd1 vssd1 vccd1 vccd1 _14747_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11959_ hold4032/X _12365_/B _11958_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _11959_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14678_ _14732_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14678_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17466_ _17468_/CLK _17466_/D vssd1 vssd1 vccd1 vccd1 _17466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16417_ _18394_/CLK _16417_/D vssd1 vssd1 vccd1 vccd1 _16417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13629_ _13734_/A _13629_/B vssd1 vssd1 vccd1 vccd1 _13629_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17397_ _18451_/CLK _17397_/D vssd1 vssd1 vccd1 vccd1 _17397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6008 _17539_/Q vssd1 vssd1 vccd1 vccd1 hold6008/X sky130_fd_sc_hd__dlygate4sd3_1
X_16348_ _18389_/CLK _16348_/D vssd1 vssd1 vccd1 vccd1 _16348_/Q sky130_fd_sc_hd__dfxtp_1
Xhold6019 _17555_/Q vssd1 vssd1 vccd1 vccd1 hold6019/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5307 _17007_/Q vssd1 vssd1 vccd1 vccd1 hold5307/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16279_ _17380_/CLK _16279_/D vssd1 vssd1 vccd1 vccd1 _16279_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5318 _10729_/X vssd1 vssd1 vccd1 vccd1 _16733_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5329 _17068_/Q vssd1 vssd1 vccd1 vccd1 hold5329/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4606 _16467_/Q vssd1 vssd1 vccd1 vccd1 hold4606/X sky130_fd_sc_hd__dlygate4sd3_1
X_18018_ _18052_/CLK _18018_/D vssd1 vssd1 vccd1 vccd1 _18018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4617 _10771_/X vssd1 vssd1 vccd1 vccd1 _16747_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4628 _16636_/Q vssd1 vssd1 vccd1 vccd1 hold4628/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4639 _09853_/X vssd1 vssd1 vccd1 vccd1 _16441_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3905 _16703_/Q vssd1 vssd1 vccd1 vccd1 hold3905/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3916 _10282_/X vssd1 vssd1 vccd1 vccd1 _16584_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_240_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3927 _16835_/Q vssd1 vssd1 vccd1 vccd1 hold3927/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3938 _16701_/Q vssd1 vssd1 vccd1 vccd1 hold3938/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3949 _10336_/X vssd1 vssd1 vccd1 vccd1 _16602_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07983_ hold1344/X _07978_/B _07982_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _07983_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09722_ hold2224/X hold4145/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09723_/B sky130_fd_sc_hd__mux2_1
X_09653_ hold1432/X hold3224/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09654_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_222_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_214_1405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08604_ _09440_/B hold626/X vssd1 vssd1 vccd1 vccd1 _15924_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09584_ hold1907/X _13286_/A _10571_/C vssd1 vssd1 vccd1 vccd1 _09585_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_222_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08535_ _12394_/A hold742/X vssd1 vssd1 vccd1 vccd1 _15891_/D sky130_fd_sc_hd__and2_1
XFILLER_0_167_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08466_ _15145_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08466_/X sky130_fd_sc_hd__or2_1
XFILLER_0_212_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08397_ _14166_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08397_/X sky130_fd_sc_hd__or2_1
XFILLER_0_169_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09018_ hold673/X hold775/X _09060_/S vssd1 vssd1 vccd1 vccd1 hold776/A sky130_fd_sc_hd__mux2_1
Xhold5830 _09790_/X vssd1 vssd1 vccd1 vccd1 _16420_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5841 hold6004/X vssd1 vssd1 vccd1 vccd1 _13265_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10290_ _10386_/A _10290_/B vssd1 vssd1 vccd1 vccd1 _10290_/X sky130_fd_sc_hd__or2_1
Xhold5852 output76/X vssd1 vssd1 vccd1 vccd1 data_out[13] sky130_fd_sc_hd__buf_12
Xhold5863 hold6019/X vssd1 vssd1 vccd1 vccd1 _13289_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5874 output85/X vssd1 vssd1 vccd1 vccd1 data_out[21] sky130_fd_sc_hd__buf_12
Xhold160 data_in[11] vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5885 hold6027/X vssd1 vssd1 vccd1 vccd1 _13113_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold171 hold604/X vssd1 vssd1 vccd1 vccd1 hold605/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5896 hold6031/X vssd1 vssd1 vccd1 vccd1 _13089_/A sky130_fd_sc_hd__buf_1
Xhold182 data_in[16] vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold193 hold193/A vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout640 _12199_/C1 vssd1 vssd1 vccd1 vccd1 _12849_/A sky130_fd_sc_hd__buf_4
Xfanout651 _12855_/A vssd1 vssd1 vccd1 vccd1 _12888_/A sky130_fd_sc_hd__buf_2
XFILLER_0_219_1305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout662 fanout739/X vssd1 vssd1 vccd1 vccd1 _12588_/A sky130_fd_sc_hd__clkbuf_8
X_13980_ _15215_/A _13986_/B vssd1 vssd1 vccd1 vccd1 _13980_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_219_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout673 fanout689/X vssd1 vssd1 vccd1 vccd1 _08351_/A sky130_fd_sc_hd__buf_2
Xfanout684 _13905_/A vssd1 vssd1 vccd1 vccd1 _14193_/C1 sky130_fd_sc_hd__buf_4
Xfanout695 _08851_/A vssd1 vssd1 vccd1 vccd1 _15284_/A sky130_fd_sc_hd__buf_4
X_12931_ hold1645/X hold4447/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12931_/X sky130_fd_sc_hd__mux2_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ _17194_/CLK _15650_/D vssd1 vssd1 vccd1 vccd1 _15650_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ hold1130/X hold3288/X _12916_/S vssd1 vssd1 vccd1 vccd1 _12862_/X sky130_fd_sc_hd__mux2_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ hold2115/X _14612_/B _14600_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _14601_/X
+ sky130_fd_sc_hd__o211a_1
X_11813_ hold2883/X hold4373/X _12293_/C vssd1 vssd1 vccd1 vccd1 _11814_/B sky130_fd_sc_hd__mux2_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15581_ _17144_/CLK _15581_/D vssd1 vssd1 vccd1 vccd1 _15581_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12793_ hold3004/X hold3392/X _12838_/S vssd1 vssd1 vccd1 vccd1 _12793_/X sky130_fd_sc_hd__mux2_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17320_ _17320_/CLK hold72/X vssd1 vssd1 vccd1 vccd1 _17320_/Q sky130_fd_sc_hd__dfxtp_1
X_14532_ hold1885/X _14537_/B _14531_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _14532_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _17072_/Q _11744_/B _12317_/C vssd1 vssd1 vccd1 vccd1 _11744_/X sky130_fd_sc_hd__and3_1
XFILLER_0_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _14517_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14463_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17251_ _17749_/CLK _17251_/D vssd1 vssd1 vccd1 vccd1 _17251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11675_ hold2053/X hold5679/X _12242_/S vssd1 vssd1 vccd1 vccd1 _11676_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16202_ _17435_/CLK _16202_/D vssd1 vssd1 vccd1 vccd1 _16202_/Q sky130_fd_sc_hd__dfxtp_1
X_13414_ hold4785/X _13814_/B _13413_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _13414_/X
+ sky130_fd_sc_hd__o211a_1
X_10626_ hold3420/X _10530_/A _10625_/X vssd1 vssd1 vccd1 vccd1 _10626_/Y sky130_fd_sc_hd__a21oi_1
X_17182_ _17278_/CLK _17182_/D vssd1 vssd1 vccd1 vccd1 _17182_/Q sky130_fd_sc_hd__dfxtp_1
X_14394_ hold338/X _14502_/B vssd1 vssd1 vccd1 vccd1 _14443_/B sky130_fd_sc_hd__or2_4
XFILLER_0_10_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16133_ _17328_/CLK _16133_/D vssd1 vssd1 vccd1 vccd1 hold657/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13345_ hold4630/X _13795_/A2 _13344_/X _13729_/C1 vssd1 vssd1 vccd1 vccd1 _13345_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10557_ _11091_/A _10557_/B vssd1 vssd1 vccd1 vccd1 _10557_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16064_ _17314_/CLK _16064_/D vssd1 vssd1 vccd1 vccd1 hold730/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13276_ hold4347/X _13275_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13276_/X sky130_fd_sc_hd__mux2_2
X_10488_ _10524_/A _10488_/B vssd1 vssd1 vccd1 vccd1 _10488_/X sky130_fd_sc_hd__or2_1
X_15015_ hold3051/X hold447/X _15014_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _15015_/X
+ sky130_fd_sc_hd__o211a_1
X_12227_ hold2365/X _17233_/Q _12227_/S vssd1 vssd1 vccd1 vccd1 _12228_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_236_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12158_ hold1082/X _17210_/Q _12332_/C vssd1 vssd1 vccd1 vccd1 _12159_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_235_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_235_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11109_ _11109_/A _11109_/B vssd1 vssd1 vccd1 vccd1 _11109_/X sky130_fd_sc_hd__or2_1
X_12089_ hold2859/X hold4857/X _13886_/C vssd1 vssd1 vccd1 vccd1 _12090_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16966_ _17846_/CLK _16966_/D vssd1 vssd1 vccd1 vccd1 _16966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15917_ _16093_/CLK _15917_/D vssd1 vssd1 vccd1 vccd1 hold498/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16897_ _18070_/CLK _16897_/D vssd1 vssd1 vccd1 vccd1 _16897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ _17707_/CLK _15848_/D vssd1 vssd1 vccd1 vccd1 _15848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15779_ _17678_/CLK _15779_/D vssd1 vssd1 vccd1 vccd1 _15779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08320_ hold2559/X _08323_/B _08319_/Y _08363_/A vssd1 vssd1 vccd1 vccd1 _08320_/X
+ sky130_fd_sc_hd__o211a_1
X_17518_ _17525_/CLK _17518_/D vssd1 vssd1 vccd1 vccd1 hold948/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08251_ hold2762/X _08262_/B _08250_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08251_/X
+ sky130_fd_sc_hd__o211a_1
X_17449_ _17450_/CLK _17449_/D vssd1 vssd1 vccd1 vccd1 _17449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_235_wb_clk_i clkbuf_6_62_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18180_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_144_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08182_ hold2733/X _08209_/B _08181_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _08182_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5104 _11272_/X vssd1 vssd1 vccd1 vccd1 _16914_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5115 _17003_/Q vssd1 vssd1 vccd1 vccd1 hold5115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5126 _12208_/X vssd1 vssd1 vccd1 vccd1 _17226_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5137 _17216_/Q vssd1 vssd1 vccd1 vccd1 hold5137/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4403 _13839_/Y vssd1 vssd1 vccd1 vccd1 _13840_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5148 _17008_/Q vssd1 vssd1 vccd1 vccd1 hold5148/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5159 _16785_/Q vssd1 vssd1 vccd1 vccd1 hold5159/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4414 _16738_/Q vssd1 vssd1 vccd1 vccd1 hold4414/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4425 _13875_/Y vssd1 vssd1 vccd1 vccd1 _13876_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4436 _16566_/Q vssd1 vssd1 vccd1 vccd1 hold4436/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4447 _17488_/Q vssd1 vssd1 vccd1 vccd1 hold4447/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3702 _17166_/Q vssd1 vssd1 vccd1 vccd1 hold3702/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3713 _10243_/X vssd1 vssd1 vccd1 vccd1 _16571_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4458 _17580_/Q vssd1 vssd1 vccd1 vccd1 hold4458/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3724 _16808_/Q vssd1 vssd1 vccd1 vccd1 hold3724/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4469 _16714_/Q vssd1 vssd1 vccd1 vccd1 hold4469/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3735 _09631_/X vssd1 vssd1 vccd1 vccd1 _16367_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3746 _16425_/Q vssd1 vssd1 vccd1 vccd1 hold3746/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3757 _16625_/Q vssd1 vssd1 vccd1 vccd1 hold3757/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3768 _12761_/X vssd1 vssd1 vccd1 vccd1 _12762_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3779 _16569_/Q vssd1 vssd1 vccd1 vccd1 hold3779/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07966_ _09313_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07966_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09705_ _09987_/A _09705_/B vssd1 vssd1 vccd1 vccd1 _09705_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07897_ hold978/X _07918_/B _07896_/X _08135_/A vssd1 vssd1 vccd1 vccd1 hold979/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09636_ _09933_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _09636_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09567_ _09978_/A _09567_/B vssd1 vssd1 vccd1 vccd1 _09567_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08518_ hold2355/X _08503_/Y _08517_/X _08167_/A vssd1 vssd1 vccd1 vccd1 _08518_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09498_ _09498_/A _09498_/B _09498_/C _09498_/D vssd1 vssd1 vccd1 vccd1 _12510_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_0_33_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08449_ _08504_/A hold406/X vssd1 vssd1 vccd1 vccd1 _08498_/B sky130_fd_sc_hd__or2_4
XFILLER_0_37_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ _11556_/A _11460_/B vssd1 vssd1 vccd1 vccd1 _11460_/X sky130_fd_sc_hd__or2_1
Xwire337 wire337/A vssd1 vssd1 vccd1 vccd1 wire337/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_184_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10411_ hold3805/X _10637_/B _10410_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10411_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11391_ _12243_/A _11391_/B vssd1 vssd1 vccd1 vccd1 _11391_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13130_ _17567_/Q _17101_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13130_/X sky130_fd_sc_hd__mux2_1
X_10342_ hold4628/X _10628_/B _10341_/X _14342_/A vssd1 vssd1 vccd1 vccd1 _10342_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13061_ _13060_/X hold5163/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13061_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_131_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5660 _11335_/X vssd1 vssd1 vccd1 vccd1 _16935_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10273_ hold3742/X _10601_/B _10272_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10273_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5671 _17203_/Q vssd1 vssd1 vccd1 vccd1 hold5671/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5682 _12109_/X vssd1 vssd1 vccd1 vccd1 _17193_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5693 _16953_/Q vssd1 vssd1 vccd1 vccd1 hold5693/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12012_ _12210_/A _12012_/B vssd1 vssd1 vccd1 vccd1 _12012_/X sky130_fd_sc_hd__or2_1
Xhold4970 _17189_/Q vssd1 vssd1 vccd1 vccd1 hold4970/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4981 _17621_/Q vssd1 vssd1 vccd1 vccd1 hold4981/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4992 _11008_/X vssd1 vssd1 vccd1 vccd1 _16826_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_39_wb_clk_i clkbuf_6_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18430_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16820_ _18023_/CLK _16820_/D vssd1 vssd1 vccd1 vccd1 _16820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout470 _12371_/C vssd1 vssd1 vccd1 vccd1 _13748_/S sky130_fd_sc_hd__buf_6
Xfanout481 fanout485/X vssd1 vssd1 vccd1 vccd1 _11774_/C sky130_fd_sc_hd__buf_4
XFILLER_0_233_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout492 _10964_/S vssd1 vssd1 vccd1 vccd1 _11201_/C sky130_fd_sc_hd__buf_4
X_16751_ _18019_/CLK _16751_/D vssd1 vssd1 vccd1 vccd1 _16751_/Q sky130_fd_sc_hd__dfxtp_1
X_13963_ hold1658/X _13995_/A2 _13962_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _13963_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_221_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15702_ _17272_/CLK _15702_/D vssd1 vssd1 vccd1 vccd1 _15702_/Q sky130_fd_sc_hd__dfxtp_1
X_12914_ hold3334/X _12913_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12915_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_232_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16682_ _18363_/CLK _16682_/D vssd1 vssd1 vccd1 vccd1 _16682_/Q sky130_fd_sc_hd__dfxtp_1
X_13894_ _14164_/A hold1943/X hold297/X vssd1 vssd1 vccd1 vccd1 _13894_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_216_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18421_ _18421_/CLK _18421_/D vssd1 vssd1 vccd1 vccd1 _18421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12845_ hold3368/X _12844_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12845_/X sky130_fd_sc_hd__mux2_1
X_15633_ _17261_/CLK _15633_/D vssd1 vssd1 vccd1 vccd1 _15633_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18352_ _18352_/CLK _18352_/D vssd1 vssd1 vccd1 vccd1 _18352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12776_ hold3530/X _12775_/X _12839_/S vssd1 vssd1 vccd1 vccd1 _12776_/X sky130_fd_sc_hd__mux2_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _17264_/CLK _15564_/D vssd1 vssd1 vccd1 vccd1 _15564_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _17303_/CLK _17303_/D vssd1 vssd1 vccd1 vccd1 hold518/A sky130_fd_sc_hd__dfxtp_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14515_ _14980_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14515_/X sky130_fd_sc_hd__or2_1
X_11727_ hold4454/X _11631_/A _11726_/X vssd1 vssd1 vccd1 vccd1 _11727_/Y sky130_fd_sc_hd__a21oi_1
X_18283_ _18315_/CLK _18283_/D vssd1 vssd1 vccd1 vccd1 _18283_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15495_ _14166_/A hold1422/X _15505_/S vssd1 vssd1 vccd1 vccd1 _15496_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_84_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17234_ _17266_/CLK _17234_/D vssd1 vssd1 vccd1 vccd1 _17234_/Q sky130_fd_sc_hd__dfxtp_1
X_11658_ _11658_/A _11658_/B vssd1 vssd1 vccd1 vccd1 _11658_/X sky130_fd_sc_hd__or2_1
X_14446_ hold1067/X _14446_/A2 _14445_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _14446_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10609_ _10651_/A _10609_/B vssd1 vssd1 vccd1 vccd1 _16693_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_141_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17165_ _17261_/CLK _17165_/D vssd1 vssd1 vccd1 vccd1 _17165_/Q sky130_fd_sc_hd__dfxtp_1
X_14377_ hold220/A _17988_/Q _14381_/S vssd1 vssd1 vccd1 vccd1 hold151/A sky130_fd_sc_hd__mux2_1
X_11589_ _12219_/A _11589_/B vssd1 vssd1 vccd1 vccd1 _11589_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold907 hold907/A vssd1 vssd1 vccd1 vccd1 hold907/X sky130_fd_sc_hd__buf_4
XFILLER_0_40_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16116_ _17339_/CLK _16116_/D vssd1 vssd1 vccd1 vccd1 hold686/A sky130_fd_sc_hd__dfxtp_1
Xhold918 hold918/A vssd1 vssd1 vccd1 vccd1 hold918/X sky130_fd_sc_hd__dlygate4sd3_1
X_13328_ hold1376/X hold5723/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13329_/B sky130_fd_sc_hd__mux2_1
Xhold929 hold929/A vssd1 vssd1 vccd1 vccd1 hold929/X sky130_fd_sc_hd__dlygate4sd3_1
X_17096_ _17628_/CLK _17096_/D vssd1 vssd1 vccd1 vccd1 _17096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16047_ _18419_/CLK _16047_/D vssd1 vssd1 vccd1 vccd1 hold346/A sky130_fd_sc_hd__dfxtp_1
X_13259_ _13258_/X hold3788/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13259_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3009 _15094_/X vssd1 vssd1 vccd1 vccd1 _18331_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2308 _17902_/Q vssd1 vssd1 vccd1 vccd1 hold2308/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2319 _07866_/X vssd1 vssd1 vccd1 vccd1 _15578_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07820_ hold353/X _14555_/C _14735_/A _09495_/C vssd1 vssd1 vccd1 vccd1 _09122_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_0_224_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1607 _18368_/Q vssd1 vssd1 vccd1 vccd1 hold1607/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1618 _16149_/Q vssd1 vssd1 vccd1 vccd1 hold1618/X sky130_fd_sc_hd__dlygate4sd3_1
X_17998_ _18030_/CLK _17998_/D vssd1 vssd1 vccd1 vccd1 _17998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1629 _13951_/X vssd1 vssd1 vccd1 vccd1 _17782_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16949_ _17831_/CLK _16949_/D vssd1 vssd1 vccd1 vccd1 _16949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09421_ _07804_/A _09463_/B _15284_/A _09420_/X vssd1 vssd1 vccd1 vccd1 _09421_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09352_ hold597/A hold384/A _15182_/A _09352_/D vssd1 vssd1 vccd1 vccd1 _09366_/B
+ sky130_fd_sc_hd__or4_2
Xclkbuf_leaf_416_wb_clk_i clkbuf_6_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17878_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08303_ _14413_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08303_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09283_ _15559_/A hold954/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09284_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_191_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08234_ hold911/X _08280_/B vssd1 vssd1 vccd1 vccd1 _08234_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08165_ _08171_/A _08165_/B vssd1 vssd1 vccd1 vccd1 _15720_/D sky130_fd_sc_hd__and2_1
XFILLER_0_28_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08096_ _14960_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08096_/X sky130_fd_sc_hd__or2_1
Xhold4200 _15313_/X vssd1 vssd1 vccd1 vccd1 _15314_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4211 hold5954/X vssd1 vssd1 vccd1 vccd1 hold5955/A sky130_fd_sc_hd__buf_4
XFILLER_0_105_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4222 _15393_/X vssd1 vssd1 vccd1 vccd1 _15394_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4233 _16340_/Q vssd1 vssd1 vccd1 vccd1 _13190_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4244 _13822_/Y vssd1 vssd1 vccd1 vccd1 _17727_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3510 _16344_/Q vssd1 vssd1 vccd1 vccd1 _13222_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold4255 _10020_/Y vssd1 vssd1 vccd1 vccd1 _10021_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4266 _10033_/Y vssd1 vssd1 vccd1 vccd1 _16501_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3521 _11742_/Y vssd1 vssd1 vccd1 vccd1 _11743_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4277 _09993_/Y vssd1 vssd1 vccd1 vccd1 _09994_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3532 _17434_/Q vssd1 vssd1 vccd1 vccd1 hold3532/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_227_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3543 _16474_/Q vssd1 vssd1 vccd1 vccd1 hold3543/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4288 _13833_/Y vssd1 vssd1 vccd1 vccd1 _13834_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3554 _16508_/Q vssd1 vssd1 vccd1 vccd1 hold3554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4299 _12321_/Y vssd1 vssd1 vccd1 vccd1 _12322_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2820 _15176_/X vssd1 vssd1 vccd1 vccd1 _18371_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3565 _09523_/X vssd1 vssd1 vccd1 vccd1 _16331_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3576 _16459_/Q vssd1 vssd1 vccd1 vccd1 hold3576/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2831 _09101_/X vssd1 vssd1 vccd1 vccd1 _16165_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3587 _09619_/X vssd1 vssd1 vccd1 vccd1 _16363_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08998_ _12440_/A hold687/X vssd1 vssd1 vccd1 vccd1 _16116_/D sky130_fd_sc_hd__and2_1
Xhold2842 _18276_/Q vssd1 vssd1 vccd1 vccd1 hold2842/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2853 _15216_/X vssd1 vssd1 vccd1 vccd1 _18390_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3598 _09979_/X vssd1 vssd1 vccd1 vccd1 _16483_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2864 _15514_/X vssd1 vssd1 vccd1 vccd1 _18435_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2875 _18260_/Q vssd1 vssd1 vccd1 vccd1 hold2875/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07949_ hold2310/X _07991_/A2 _07948_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _07949_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2886 _18091_/Q vssd1 vssd1 vccd1 vccd1 hold2886/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2897 _15785_/Q vssd1 vssd1 vccd1 vccd1 hold2897/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10960_ hold5569/X _11726_/B _10959_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _10960_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_230_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09619_ hold3586/X _10025_/B _09618_/X _15473_/A vssd1 vssd1 vccd1 vccd1 _09619_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10891_ hold5157/X _11171_/B _10890_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _10891_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12630_ _12864_/A _12630_/B vssd1 vssd1 vccd1 vccd1 _17386_/D sky130_fd_sc_hd__and2_1
XFILLER_0_210_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_157_wb_clk_i clkbuf_6_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17338_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_168_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12561_ _12906_/A _12561_/B vssd1 vssd1 vccd1 vccd1 _17363_/D sky130_fd_sc_hd__and2_1
XFILLER_0_93_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14300_ _14980_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14300_/X sky130_fd_sc_hd__or2_1
X_11512_ hold4895/X _11798_/B _11511_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _11512_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15280_ hold620/X _15448_/A2 _15446_/B1 hold772/X vssd1 vssd1 vccd1 vccd1 _15280_/X
+ sky130_fd_sc_hd__a22o_1
X_12492_ _17339_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12492_/X sky130_fd_sc_hd__or2_1
XFILLER_0_135_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14231_ hold2514/X _14216_/Y _14230_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _14231_/X
+ sky130_fd_sc_hd__o211a_1
X_11443_ hold5115/X _11726_/B _11442_/X _13895_/A vssd1 vssd1 vccd1 vccd1 _11443_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14162_ hold330/X _14163_/B vssd1 vssd1 vccd1 vccd1 _14162_/Y sky130_fd_sc_hd__nor2_2
X_11374_ hold5531/X _11195_/B _11373_/X _14462_/C1 vssd1 vssd1 vccd1 vccd1 _11374_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13113_ _13113_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13113_/X sky130_fd_sc_hd__and2_1
X_10325_ hold1712/X _16599_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10326_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14093_ hold2520/X _14094_/B _14092_/Y _13895_/A vssd1 vssd1 vccd1 vccd1 _14093_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ hold937/X hold901/X _13043_/X hold935/X vssd1 vssd1 vccd1 vccd1 _13044_/X
+ sky130_fd_sc_hd__a211o_1
X_17921_ _18049_/CLK _17921_/D vssd1 vssd1 vccd1 vccd1 _17921_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5490 _17703_/Q vssd1 vssd1 vccd1 vccd1 hold5490/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_221_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10256_ hold1815/X hold3987/X _10646_/C vssd1 vssd1 vccd1 vccd1 _10257_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17852_ _17884_/CLK _17852_/D vssd1 vssd1 vccd1 vccd1 _17852_/Q sky130_fd_sc_hd__dfxtp_1
X_10187_ hold2516/X hold3274/X _10475_/S vssd1 vssd1 vccd1 vccd1 _10188_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_205_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16803_ _18036_/CLK _16803_/D vssd1 vssd1 vccd1 vccd1 _16803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_233_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17783_ _18429_/CLK _17783_/D vssd1 vssd1 vccd1 vccd1 _17783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14995_ hold2187/X hold447/X _14994_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _14995_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_234_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16734_ _18065_/CLK _16734_/D vssd1 vssd1 vccd1 vccd1 _16734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13946_ _14627_/A _14163_/B vssd1 vssd1 vccd1 vccd1 _13946_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_233_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_232_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16665_ _18223_/CLK _16665_/D vssd1 vssd1 vccd1 vccd1 _16665_/Q sky130_fd_sc_hd__dfxtp_1
X_13877_ _17746_/Q _13877_/B _13877_/C vssd1 vssd1 vccd1 vccd1 _13877_/X sky130_fd_sc_hd__and3_1
XFILLER_0_18_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18404_ _18404_/CLK _18404_/D vssd1 vssd1 vccd1 vccd1 _18404_/Q sky130_fd_sc_hd__dfxtp_1
X_15616_ _17262_/CLK _15616_/D vssd1 vssd1 vccd1 vccd1 _15616_/Q sky130_fd_sc_hd__dfxtp_1
X_12828_ _12837_/A _12828_/B vssd1 vssd1 vccd1 vccd1 _17452_/D sky130_fd_sc_hd__and2_1
XFILLER_0_232_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16596_ _18166_/CLK _16596_/D vssd1 vssd1 vccd1 vccd1 _16596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18335_ _18377_/CLK hold693/X vssd1 vssd1 vccd1 vccd1 _18335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15547_ _15547_/A _15547_/B vssd1 vssd1 vccd1 vccd1 _15547_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12759_ _12810_/A _12759_/B vssd1 vssd1 vccd1 vccd1 _17429_/D sky130_fd_sc_hd__and2_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18266_ _18298_/CLK _18266_/D vssd1 vssd1 vccd1 vccd1 _18266_/Q sky130_fd_sc_hd__dfxtp_1
X_15478_ hold761/X _09367_/A _09392_/C hold697/X vssd1 vssd1 vccd1 vccd1 _15478_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17217_ _17279_/CLK _17217_/D vssd1 vssd1 vccd1 vccd1 _17217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14429_ _15543_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _14429_/Y sky130_fd_sc_hd__nand2_1
X_18197_ _18197_/CLK _18197_/D vssd1 vssd1 vccd1 vccd1 _18197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold704 hold713/X vssd1 vssd1 vccd1 vccd1 hold704/X sky130_fd_sc_hd__clkbuf_4
X_17148_ _17262_/CLK _17148_/D vssd1 vssd1 vccd1 vccd1 _17148_/Q sky130_fd_sc_hd__dfxtp_1
Xhold715 hold715/A vssd1 vssd1 vccd1 vccd1 hold715/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold726 hold726/A vssd1 vssd1 vccd1 vccd1 hold726/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 hold737/A vssd1 vssd1 vccd1 vccd1 hold737/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold748 hold748/A vssd1 vssd1 vccd1 vccd1 hold748/X sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ hold3886/X _10046_/B _09969_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09970_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold759 hold759/A vssd1 vssd1 vccd1 vccd1 hold759/X sky130_fd_sc_hd__dlygate4sd3_1
X_17079_ _17895_/CLK _17079_/D vssd1 vssd1 vccd1 vccd1 _17079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08921_ _15324_/A hold439/X vssd1 vssd1 vccd1 vccd1 _16078_/D sky130_fd_sc_hd__and2_1
Xhold2105 hold2105/A vssd1 vssd1 vccd1 vccd1 _15199_/A sky130_fd_sc_hd__buf_12
XFILLER_0_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2116 _14601_/X vssd1 vssd1 vccd1 vccd1 _18094_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08852_ hold143/X hold624/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08853_/B sky130_fd_sc_hd__mux2_1
Xhold2127 _18046_/Q vssd1 vssd1 vccd1 vccd1 hold2127/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2138 _15080_/X vssd1 vssd1 vccd1 vccd1 _18324_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_237_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1404 _15761_/Q vssd1 vssd1 vccd1 vccd1 hold1404/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2149 _17913_/Q vssd1 vssd1 vccd1 vccd1 hold2149/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1415 _15524_/X vssd1 vssd1 vccd1 vccd1 _18440_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07803_ _16286_/Q _07801_/B _07802_/Y vssd1 vssd1 vccd1 vccd1 _07803_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_224_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1426 _08212_/X vssd1 vssd1 vccd1 vccd1 _15742_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08783_ hold315/X _16012_/Q _08793_/S vssd1 vssd1 vccd1 vccd1 hold316/A sky130_fd_sc_hd__mux2_1
Xhold1437 _08438_/X vssd1 vssd1 vccd1 vccd1 _15849_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1448 _17966_/Q vssd1 vssd1 vccd1 vccd1 hold1448/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1459 _15612_/Q vssd1 vssd1 vccd1 vccd1 hold1459/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09404_ _09438_/B _09404_/B vssd1 vssd1 vccd1 vccd1 _09404_/X sky130_fd_sc_hd__or2_1
XFILLER_0_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_250_wb_clk_i clkbuf_6_59_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18231_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09335_ _15557_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09335_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09266_ _09272_/A hold573/X vssd1 vssd1 vccd1 vccd1 _16244_/D sky130_fd_sc_hd__and2_1
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08217_ _14330_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08217_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09197_ hold3004/X _09214_/B _09196_/X _12798_/A vssd1 vssd1 vccd1 vccd1 _09197_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08148_ _14726_/A hold2654/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08149_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_6_44_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_44_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08079_ hold2197/X _08088_/B _08078_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _08079_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4030 _17207_/Q vssd1 vssd1 vccd1 vccd1 hold4030/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10110_ _10530_/A _10110_/B vssd1 vssd1 vccd1 vccd1 _10110_/X sky130_fd_sc_hd__or2_1
Xhold4041 _11554_/X vssd1 vssd1 vccd1 vccd1 _17008_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4052 _17456_/Q vssd1 vssd1 vccd1 vccd1 hold4052/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4063 _16831_/Q vssd1 vssd1 vccd1 vccd1 hold4063/X sky130_fd_sc_hd__dlygate4sd3_1
X_11090_ hold2981/X _16854_/Q _11186_/C vssd1 vssd1 vccd1 vccd1 _11091_/B sky130_fd_sc_hd__mux2_1
XTAP_6236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4074 _17408_/Q vssd1 vssd1 vccd1 vccd1 hold4074/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3340 _10303_/X vssd1 vssd1 vccd1 vccd1 _16591_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4085 _16772_/Q vssd1 vssd1 vccd1 vccd1 hold4085/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10041_ _13222_/A _09957_/A _10040_/X vssd1 vssd1 vccd1 vccd1 _10041_/Y sky130_fd_sc_hd__a21oi_1
Xhold4096 _10762_/X vssd1 vssd1 vccd1 vccd1 _16744_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3351 _12800_/X vssd1 vssd1 vccd1 vccd1 _12801_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3362 _17406_/Q vssd1 vssd1 vccd1 vccd1 hold3362/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3373 _17447_/Q vssd1 vssd1 vccd1 vccd1 hold3373/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold81/X vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__buf_4
XFILLER_0_220_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3384 _12692_/X vssd1 vssd1 vccd1 vccd1 _12693_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2650 _15834_/Q vssd1 vssd1 vccd1 vccd1 hold2650/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3395 _12755_/X vssd1 vssd1 vccd1 vccd1 _12756_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__buf_4
XTAP_5568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2661 _15824_/Q vssd1 vssd1 vccd1 vccd1 hold2661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold89/X vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2672 _08220_/X vssd1 vssd1 vccd1 vccd1 _15746_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2683 _18439_/Q vssd1 vssd1 vccd1 vccd1 hold2683/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2694 _14482_/X vssd1 vssd1 vccd1 vccd1 _18038_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1960 _18251_/Q vssd1 vssd1 vccd1 vccd1 hold1960/X sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ _13800_/A _13800_/B vssd1 vssd1 vccd1 vccd1 _13800_/X sky130_fd_sc_hd__or2_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_338_wb_clk_i clkbuf_6_43_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17271_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14780_ _15227_/A _14780_/B vssd1 vssd1 vccd1 vccd1 _14780_/X sky130_fd_sc_hd__or2_1
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11992_ hold5032/X _12374_/B _11991_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _11992_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1971 _14003_/X vssd1 vssd1 vccd1 vccd1 _17807_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1982 hold6122/X vssd1 vssd1 vccd1 vccd1 _09477_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1993 _09419_/X vssd1 vssd1 vccd1 vccd1 _16295_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10943_ hold2796/X _16805_/Q _11153_/C vssd1 vssd1 vccd1 vccd1 _10944_/B sky130_fd_sc_hd__mux2_1
X_13731_ _13737_/A _13731_/B vssd1 vssd1 vccd1 vccd1 _13731_/X sky130_fd_sc_hd__or2_1
XFILLER_0_230_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16450_ _18395_/CLK _16450_/D vssd1 vssd1 vccd1 vccd1 _16450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10874_ hold1772/X _16782_/Q _11162_/C vssd1 vssd1 vccd1 vccd1 _10875_/B sky130_fd_sc_hd__mux2_1
X_13662_ _13758_/A _13662_/B vssd1 vssd1 vccd1 vccd1 _13662_/X sky130_fd_sc_hd__or2_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15401_ _16304_/Q _15477_/A2 _15487_/B1 hold882/X _15400_/X vssd1 vssd1 vccd1 vccd1
+ _15402_/D sky130_fd_sc_hd__a221o_1
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12613_ hold1477/X _17382_/Q _12850_/S vssd1 vssd1 vccd1 vccd1 _12613_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16381_ _18384_/CLK _16381_/D vssd1 vssd1 vccd1 vccd1 _16381_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13593_ _13788_/A _13593_/B vssd1 vssd1 vccd1 vccd1 _13593_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18120_ _18124_/CLK _18120_/D vssd1 vssd1 vccd1 vccd1 _18120_/Q sky130_fd_sc_hd__dfxtp_1
X_15332_ _15489_/A _15332_/B _15332_/C _15332_/D vssd1 vssd1 vccd1 vccd1 _15332_/X
+ sky130_fd_sc_hd__or4_1
X_12544_ hold2926/X hold3381/X _12925_/S vssd1 vssd1 vccd1 vccd1 _12544_/X sky130_fd_sc_hd__mux2_1
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18051_ _18051_/CLK _18051_/D vssd1 vssd1 vccd1 vccd1 _18051_/Q sky130_fd_sc_hd__dfxtp_1
X_12475_ hold172/X _12509_/A2 _12501_/A3 _12474_/X _12410_/A vssd1 vssd1 vccd1 vccd1
+ hold173/A sky130_fd_sc_hd__o311a_1
X_15263_ _15490_/A1 _15255_/X _15262_/X _15490_/B1 hold5920/A vssd1 vssd1 vccd1 vccd1
+ _15263_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_48_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_227_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17002_ _17850_/CLK _17002_/D vssd1 vssd1 vccd1 vccd1 _17002_/Q sky130_fd_sc_hd__dfxtp_1
X_14214_ _15559_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14214_/X sky130_fd_sc_hd__or2_1
X_11426_ hold1481/X _16966_/Q _11717_/C vssd1 vssd1 vccd1 vccd1 _11427_/B sky130_fd_sc_hd__mux2_1
XANTENNA_6 _13068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15194_ hold2948/X _15221_/B _15193_/X _15202_/C1 vssd1 vssd1 vccd1 vccd1 _15194_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_54_wb_clk_i clkbuf_6_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18048_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14145_ hold2481/X _14148_/B _14144_/Y _14211_/C1 vssd1 vssd1 vccd1 vccd1 _14145_/X
+ sky130_fd_sc_hd__o211a_1
X_11357_ hold2532/X hold4877/X _11654_/S vssd1 vssd1 vccd1 vccd1 _11358_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10308_ _10536_/A _10308_/B vssd1 vssd1 vccd1 vccd1 _10308_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14076_ _15203_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14076_/X sky130_fd_sc_hd__or2_1
X_11288_ hold1413/X hold4353/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11289_/B sky130_fd_sc_hd__mux2_1
X_13027_ _13034_/D hold904/X vssd1 vssd1 vccd1 vccd1 _13029_/B sky130_fd_sc_hd__and2_1
XFILLER_0_24_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17904_ _17904_/CLK _17904_/D vssd1 vssd1 vccd1 vccd1 _17904_/Q sky130_fd_sc_hd__dfxtp_1
X_10239_ _10554_/A _10239_/B vssd1 vssd1 vccd1 vccd1 _10239_/X sky130_fd_sc_hd__or2_1
XFILLER_0_219_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17835_ _17867_/CLK _17835_/D vssd1 vssd1 vccd1 vccd1 _17835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_234_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17766_ _17832_/CLK _17766_/D vssd1 vssd1 vccd1 vccd1 _17766_/Q sky130_fd_sc_hd__dfxtp_1
X_14978_ hold423/X _15018_/B vssd1 vssd1 vccd1 vccd1 _14978_/X sky130_fd_sc_hd__or2_1
XFILLER_0_178_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16717_ _18048_/CLK _16717_/D vssd1 vssd1 vccd1 vccd1 _16717_/Q sky130_fd_sc_hd__dfxtp_1
X_13929_ _13929_/A hold554/X vssd1 vssd1 vccd1 vccd1 hold555/A sky130_fd_sc_hd__and2_1
XFILLER_0_77_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17697_ _17697_/CLK _17697_/D vssd1 vssd1 vccd1 vccd1 _17697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16648_ _18265_/CLK _16648_/D vssd1 vssd1 vccd1 vccd1 _16648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16579_ _18233_/CLK _16579_/D vssd1 vssd1 vccd1 vccd1 _16579_/Q sky130_fd_sc_hd__dfxtp_1
X_09120_ _18459_/Q _11158_/A _18462_/Q vssd1 vssd1 vccd1 vccd1 _09120_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_130_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18318_ _18378_/CLK _18318_/D vssd1 vssd1 vccd1 vccd1 _18318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09051_ _12394_/A _09051_/B vssd1 vssd1 vccd1 vccd1 _16142_/D sky130_fd_sc_hd__and2_1
X_18249_ _18379_/CLK _18249_/D vssd1 vssd1 vccd1 vccd1 _18249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08002_ hold2470/X _08033_/B _08001_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _08002_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold501 hold501/A vssd1 vssd1 vccd1 vccd1 hold501/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold512 hold512/A vssd1 vssd1 vccd1 vccd1 hold512/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 hold523/A vssd1 vssd1 vccd1 vccd1 hold523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 hold534/A vssd1 vssd1 vccd1 vccd1 hold534/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold545 hold545/A vssd1 vssd1 vccd1 vccd1 hold545/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold556 hold556/A vssd1 vssd1 vccd1 vccd1 hold556/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold567 hold567/A vssd1 vssd1 vccd1 vccd1 hold567/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 input54/X vssd1 vssd1 vccd1 vccd1 hold578/X sky130_fd_sc_hd__dlymetal6s2s_1
X_09953_ _18388_/Q hold3582/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09954_/B sky130_fd_sc_hd__mux2_1
Xhold589 hold589/A vssd1 vssd1 vccd1 vccd1 hold589/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08904_ hold254/X hold426/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08905_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_0_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09884_ hold2422/X hold5829/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09885_/B sky130_fd_sc_hd__mux2_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1201 _17831_/Q vssd1 vssd1 vccd1 vccd1 hold1201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 _14939_/X vssd1 vssd1 vccd1 vccd1 _18256_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08835_ _12416_/A hold591/X vssd1 vssd1 vccd1 vccd1 _16036_/D sky130_fd_sc_hd__and2_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1223 hold1223/A vssd1 vssd1 vccd1 vccd1 input51/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1234 _14067_/X vssd1 vssd1 vccd1 vccd1 _17838_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1245 _14855_/X vssd1 vssd1 vccd1 vccd1 _18216_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 _15689_/Q vssd1 vssd1 vccd1 vccd1 hold1256/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08766_ _15344_/A _08766_/B vssd1 vssd1 vccd1 vccd1 _16003_/D sky130_fd_sc_hd__and2_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1267 _15774_/Q vssd1 vssd1 vccd1 vccd1 hold1267/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_431_wb_clk_i clkbuf_6_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17729_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1278 _08061_/X vssd1 vssd1 vccd1 vccd1 _15670_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1289 _17793_/Q vssd1 vssd1 vccd1 vccd1 hold1289/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08697_ hold185/X hold205/X _08721_/S vssd1 vssd1 vccd1 vccd1 hold206/A sky130_fd_sc_hd__mux2_1
XFILLER_0_200_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09318_ hold2159/X _09323_/B _09317_/X _12588_/A vssd1 vssd1 vccd1 vccd1 _09318_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10590_ _16527_/Q _10470_/A _10589_/X vssd1 vssd1 vccd1 vccd1 _10590_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09249_ _15525_/A hold2935/X hold271/X vssd1 vssd1 vccd1 vccd1 _09250_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_145_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12260_ hold1865/X hold5036/X _13481_/S vssd1 vssd1 vccd1 vccd1 _12261_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_224_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11211_ hold3512/X _11100_/A _11210_/X vssd1 vssd1 vccd1 vccd1 _11211_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12191_ hold2474/X _17221_/Q _13409_/S vssd1 vssd1 vccd1 vccd1 _12192_/B sky130_fd_sc_hd__mux2_1
XTAP_6000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11142_ hold3442/X _11049_/A _11141_/X vssd1 vssd1 vccd1 vccd1 _11142_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput76 _13161_/A vssd1 vssd1 vccd1 vccd1 output76/X sky130_fd_sc_hd__buf_6
XTAP_6033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput87 _13241_/A vssd1 vssd1 vccd1 vccd1 output87/X sky130_fd_sc_hd__buf_6
XTAP_6044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15950_ _17297_/CLK _15950_/D vssd1 vssd1 vccd1 vccd1 hold102/A sky130_fd_sc_hd__dfxtp_1
XTAP_6055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11073_ _11649_/A _11073_/B vssd1 vssd1 vccd1 vccd1 _11073_/X sky130_fd_sc_hd__or2_1
Xoutput98 _13089_/A vssd1 vssd1 vccd1 vccd1 output98/X sky130_fd_sc_hd__buf_6
XTAP_5321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3170 _14402_/X vssd1 vssd1 vccd1 vccd1 _17999_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14901_ hold2085/X _14896_/Y _14900_/X _15042_/A vssd1 vssd1 vccd1 vccd1 _18238_/D
+ sky130_fd_sc_hd__o211a_1
X_10024_ _11158_/A _10024_/B vssd1 vssd1 vccd1 vccd1 _16498_/D sky130_fd_sc_hd__nor2_1
Xhold3181 _14241_/X vssd1 vssd1 vccd1 vccd1 _17921_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3192 _16335_/Q vssd1 vssd1 vccd1 vccd1 _13150_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15881_ _17222_/CLK _15881_/D vssd1 vssd1 vccd1 vccd1 _15881_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17620_ _17620_/CLK _17620_/D vssd1 vssd1 vccd1 vccd1 _17620_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2480 _09163_/X vssd1 vssd1 vccd1 vccd1 _16194_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2491 _18085_/Q vssd1 vssd1 vccd1 vccd1 hold2491/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14832_ _15225_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14832_/X sky130_fd_sc_hd__or2_1
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_172_wb_clk_i clkbuf_6_48_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18347_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ _18223_/CLK _17551_/D vssd1 vssd1 vccd1 vccd1 _17551_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1790 _15104_/X vssd1 vssd1 vccd1 vccd1 _18336_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_101_wb_clk_i clkbuf_6_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18409_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14763_ hold2111/X _14772_/B _14762_/X _14769_/C1 vssd1 vssd1 vccd1 vccd1 _14763_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11975_ hold1256/X _17149_/Q _12332_/C vssd1 vssd1 vccd1 vccd1 _11976_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_59_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _18325_/CLK _16502_/D vssd1 vssd1 vccd1 vccd1 _16502_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13714_ hold5779/X _13808_/B _13713_/X _12804_/A vssd1 vssd1 vccd1 vccd1 _13714_/X
+ sky130_fd_sc_hd__o211a_1
X_10926_ _11088_/A _10926_/B vssd1 vssd1 vccd1 vccd1 _10926_/X sky130_fd_sc_hd__or2_1
X_17482_ _17484_/CLK _17482_/D vssd1 vssd1 vccd1 vccd1 _17482_/Q sky130_fd_sc_hd__dfxtp_1
X_14694_ _14980_/A _14730_/B vssd1 vssd1 vccd1 vccd1 _14694_/X sky130_fd_sc_hd__or2_1
XFILLER_0_184_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16433_ _18323_/CLK _16433_/D vssd1 vssd1 vccd1 vccd1 _16433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10857_ _11049_/A _10857_/B vssd1 vssd1 vccd1 vccd1 _10857_/X sky130_fd_sc_hd__or2_1
X_13645_ hold5281/X _13856_/B _13644_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13645_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16364_ _18349_/CLK _16364_/D vssd1 vssd1 vccd1 vccd1 _16364_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _11010_/A _10788_/B vssd1 vssd1 vccd1 vccd1 _10788_/X sky130_fd_sc_hd__or2_1
X_13576_ hold3738/X _13795_/A2 _13575_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13576_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _18232_/CLK _18103_/D vssd1 vssd1 vccd1 vccd1 _18103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15315_ hold699/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15315_/X sky130_fd_sc_hd__or2_1
XFILLER_0_171_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12527_ hold3638/X _12526_/X _12929_/S vssd1 vssd1 vccd1 vccd1 _12527_/X sky130_fd_sc_hd__mux2_1
X_16295_ _18460_/CLK _16295_/D vssd1 vssd1 vccd1 vccd1 _16295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18034_ _18126_/CLK _18034_/D vssd1 vssd1 vccd1 vccd1 _18034_/Q sky130_fd_sc_hd__dfxtp_1
X_15246_ _17328_/Q _15486_/B1 _15485_/B1 hold541/X vssd1 vssd1 vccd1 vccd1 _15246_/X
+ sky130_fd_sc_hd__a22o_1
X_12458_ _17322_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12458_/X sky130_fd_sc_hd__or2_1
XFILLER_0_169_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11409_ _12240_/A _11409_/B vssd1 vssd1 vccd1 vccd1 _11409_/X sky130_fd_sc_hd__or2_1
X_15177_ _15231_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15177_/X sky130_fd_sc_hd__or2_1
X_12389_ hold71/X hold805/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12390_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14128_ _14413_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14128_/X sky130_fd_sc_hd__or2_1
XFILLER_0_185_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14059_ hold1742/X _14107_/A2 _14058_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _14059_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08620_ _12420_/A _08620_/B vssd1 vssd1 vccd1 vccd1 _15932_/D sky130_fd_sc_hd__and2_1
XFILLER_0_59_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17818_ _17850_/CLK _17818_/D vssd1 vssd1 vccd1 vccd1 _17818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08551_ _12418_/A hold850/X vssd1 vssd1 vccd1 vccd1 _15899_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17749_ _17749_/CLK _17749_/D vssd1 vssd1 vccd1 vccd1 _17749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08482_ _15541_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _08482_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_203_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09103_ hold2611/X _09102_/B _09102_/Y _12978_/A vssd1 vssd1 vccd1 vccd1 _09103_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09034_ hold254/X hold303/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09035_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold320 hold44/X vssd1 vssd1 vccd1 vccd1 hold320/X sky130_fd_sc_hd__buf_4
Xhold331 hold331/A vssd1 vssd1 vccd1 vccd1 hold331/X sky130_fd_sc_hd__buf_2
Xhold342 hold342/A vssd1 vssd1 vccd1 vccd1 hold342/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 hold353/A vssd1 vssd1 vccd1 vccd1 hold353/X sky130_fd_sc_hd__buf_2
Xhold364 hold364/A vssd1 vssd1 vccd1 vccd1 hold364/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 hold627/X vssd1 vssd1 vccd1 vccd1 hold628/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold386 hold386/A vssd1 vssd1 vccd1 vccd1 hold386/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout800 fanout816/X vssd1 vssd1 vccd1 vccd1 _15160_/C1 sky130_fd_sc_hd__buf_2
Xhold397 hold397/A vssd1 vssd1 vccd1 vccd1 hold397/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 _15228_/C1 vssd1 vssd1 vccd1 vccd1 _15026_/A sky130_fd_sc_hd__buf_4
XFILLER_0_110_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09936_ _09948_/A _09936_/B vssd1 vssd1 vccd1 vccd1 _09936_/X sky130_fd_sc_hd__or2_1
Xfanout822 _10564_/C1 vssd1 vssd1 vccd1 vccd1 _14697_/C1 sky130_fd_sc_hd__buf_2
Xfanout833 fanout843/X vssd1 vssd1 vccd1 vccd1 _14893_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_176_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout844 _13864_/A vssd1 vssd1 vccd1 vccd1 _13819_/A sky130_fd_sc_hd__buf_8
XFILLER_0_42_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout855 _11218_/A vssd1 vssd1 vccd1 vccd1 _10651_/A sky130_fd_sc_hd__buf_8
Xfanout866 _15217_/A vssd1 vssd1 vccd1 vccd1 _15543_/A sky130_fd_sc_hd__clkbuf_16
X_09867_ _09957_/A _09867_/B vssd1 vssd1 vccd1 vccd1 _09867_/X sky130_fd_sc_hd__or2_1
Xfanout877 hold951/X vssd1 vssd1 vccd1 vccd1 _15201_/A sky130_fd_sc_hd__clkbuf_8
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout888 hold1464/X vssd1 vssd1 vccd1 vccd1 hold1465/A sky130_fd_sc_hd__buf_6
Xhold1020 hold913/X vssd1 vssd1 vccd1 vccd1 input48/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1031 _18327_/Q vssd1 vssd1 vccd1 vccd1 hold1031/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout899 hold1579/X vssd1 vssd1 vccd1 vccd1 hold1580/A sky130_fd_sc_hd__buf_6
Xhold1042 _14643_/X vssd1 vssd1 vccd1 vccd1 _18114_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ hold679/X hold837/X _08860_/S vssd1 vssd1 vccd1 vccd1 hold838/A sky130_fd_sc_hd__mux2_1
Xhold1053 _08410_/X vssd1 vssd1 vccd1 vccd1 _15835_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09798_ _09984_/A _09798_/B vssd1 vssd1 vccd1 vccd1 _09798_/X sky130_fd_sc_hd__or2_1
Xhold1064 _18204_/Q vssd1 vssd1 vccd1 vccd1 hold1064/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_240_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1075 hold1147/X vssd1 vssd1 vccd1 vccd1 hold1075/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1086 _13999_/X vssd1 vssd1 vccd1 vccd1 _17806_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 _17775_/Q vssd1 vssd1 vccd1 vccd1 hold1097/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ hold673/X hold779/X _08779_/S vssd1 vssd1 vccd1 vccd1 hold780/A sky130_fd_sc_hd__mux2_1
XFILLER_0_169_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ hold4384/X _11670_/A _11759_/X vssd1 vssd1 vccd1 vccd1 _11760_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_240_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_230_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10711_ hold3960/X _10616_/B _10710_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10711_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _12234_/A _11691_/B vssd1 vssd1 vccd1 vccd1 _11691_/X sky130_fd_sc_hd__or2_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10642_ _10651_/A _10642_/B vssd1 vssd1 vccd1 vccd1 _16704_/D sky130_fd_sc_hd__nor2_1
X_13430_ hold2650/X hold4075/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13431_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_76_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13361_ hold2716/X hold4498/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13362_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10573_ _10603_/A _10573_/B vssd1 vssd1 vccd1 vccd1 _16681_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_183_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15100_ hold2695/X hold341/X _15099_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _15100_/X
+ sky130_fd_sc_hd__o211a_1
X_12312_ hold4343/X _13314_/A _12311_/X vssd1 vssd1 vccd1 vccd1 _12312_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_228_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16080_ _16093_/CLK _16080_/D vssd1 vssd1 vccd1 vccd1 hold468/A sky130_fd_sc_hd__dfxtp_1
X_13292_ hold3476/X _13291_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13292_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15031_ _15193_/A hold2668/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15032_/B sky130_fd_sc_hd__mux2_1
X_12243_ _12243_/A _12243_/B vssd1 vssd1 vccd1 vccd1 _12243_/X sky130_fd_sc_hd__or2_1
XFILLER_0_224_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12174_ _12174_/A _12174_/B vssd1 vssd1 vccd1 vccd1 _12174_/X sky130_fd_sc_hd__or2_1
XFILLER_0_236_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11125_ hold3919/X _11222_/B _11124_/X _14346_/A vssd1 vssd1 vccd1 vccd1 _11125_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_353_wb_clk_i clkbuf_6_40_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17734_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16982_ _17936_/CLK _16982_/D vssd1 vssd1 vccd1 vccd1 _16982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_236_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15933_ _16139_/CLK _15933_/D vssd1 vssd1 vccd1 vccd1 hold761/A sky130_fd_sc_hd__dfxtp_1
X_11056_ hold5626/X _11726_/B _11055_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _11056_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10007_ _16493_/Q _10025_/B _10025_/C vssd1 vssd1 vccd1 vccd1 _10007_/X sky130_fd_sc_hd__and3_1
XFILLER_0_200_1292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_1311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ _17735_/CLK _15864_/D vssd1 vssd1 vccd1 vccd1 _15864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17603_ _17731_/CLK _17603_/D vssd1 vssd1 vccd1 vccd1 _17603_/Q sky130_fd_sc_hd__dfxtp_1
X_14815_ hold2879/X _14826_/B _14814_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14815_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15795_ _17718_/CLK _15795_/D vssd1 vssd1 vccd1 vccd1 _15795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17534_ _17535_/CLK _17534_/D vssd1 vssd1 vccd1 vccd1 _17534_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _15193_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14746_/X sky130_fd_sc_hd__or2_1
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11958_ _12273_/A _11958_/B vssd1 vssd1 vccd1 vccd1 _11958_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17465_ _17468_/CLK _17465_/D vssd1 vssd1 vccd1 vccd1 _17465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10909_ hold5343/X _11195_/B _10908_/X _14462_/C1 vssd1 vssd1 vccd1 vccd1 _10909_/X
+ sky130_fd_sc_hd__o211a_1
X_14677_ hold1519/X _14664_/B _14676_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14677_/X
+ sky130_fd_sc_hd__o211a_1
X_11889_ _13407_/A _11889_/B vssd1 vssd1 vccd1 vccd1 _11889_/X sky130_fd_sc_hd__or2_1
X_16416_ _18361_/CLK _16416_/D vssd1 vssd1 vccd1 vccd1 _16416_/Q sky130_fd_sc_hd__dfxtp_1
X_13628_ hold1218/X _17663_/Q _13829_/C vssd1 vssd1 vccd1 vccd1 _13629_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17396_ _18448_/CLK _17396_/D vssd1 vssd1 vccd1 vccd1 _17396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16347_ _18346_/CLK _16347_/D vssd1 vssd1 vccd1 vccd1 _16347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13559_ hold1134/X _17640_/Q _13841_/C vssd1 vssd1 vccd1 vccd1 _13560_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6009 _17549_/Q vssd1 vssd1 vccd1 vccd1 hold6009/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5308 _11455_/X vssd1 vssd1 vccd1 vccd1 _16975_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16278_ _17380_/CLK _16278_/D vssd1 vssd1 vccd1 vccd1 _16278_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5319 _17668_/Q vssd1 vssd1 vccd1 vccd1 hold5319/X sky130_fd_sc_hd__dlygate4sd3_1
X_18017_ _18048_/CLK _18017_/D vssd1 vssd1 vccd1 vccd1 _18017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15229_ _15229_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15229_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4607 _09835_/X vssd1 vssd1 vccd1 vccd1 _16435_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4618 _16435_/Q vssd1 vssd1 vccd1 vccd1 hold4618/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4629 _10342_/X vssd1 vssd1 vccd1 vccd1 _16604_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3906 _10543_/X vssd1 vssd1 vccd1 vccd1 _16671_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3917 _16769_/Q vssd1 vssd1 vccd1 vccd1 hold3917/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3928 _16879_/Q vssd1 vssd1 vccd1 vccd1 _11165_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3939 _10537_/X vssd1 vssd1 vccd1 vccd1 _16669_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07982_ _14330_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07982_/X sky130_fd_sc_hd__or2_1
X_09721_ hold4567/X _10031_/B _09720_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09721_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09652_ hold4171/X _10052_/B _09651_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09652_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08603_ hold131/X hold625/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold626/A sky130_fd_sc_hd__mux2_1
X_09583_ hold3552/X _10601_/B _09582_/X _15204_/C1 vssd1 vssd1 vccd1 vccd1 _09583_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08534_ hold618/X hold741/X _08592_/S vssd1 vssd1 vccd1 vccd1 hold742/A sky130_fd_sc_hd__mux2_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_212_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08465_ hold1043/X _08488_/B _08464_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _08465_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08396_ hold2043/X _08442_/A2 _08395_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _08396_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09017_ _15491_/A _09017_/B vssd1 vssd1 vccd1 vccd1 _16125_/D sky130_fd_sc_hd__and2_1
XFILLER_0_5_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5820 _13432_/X vssd1 vssd1 vccd1 vccd1 _17597_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5831 _16370_/Q vssd1 vssd1 vccd1 vccd1 hold5831/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5842 output90/X vssd1 vssd1 vccd1 vccd1 data_out[26] sky130_fd_sc_hd__buf_12
Xhold5853 hold6007/X vssd1 vssd1 vccd1 vccd1 _13281_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5864 output93/X vssd1 vssd1 vccd1 vccd1 data_out[29] sky130_fd_sc_hd__buf_12
XFILLER_0_44_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold150 hold219/X vssd1 vssd1 vccd1 vccd1 hold220/A sky130_fd_sc_hd__buf_6
Xhold5875 hold6021/X vssd1 vssd1 vccd1 vccd1 _13105_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 hold1/X vssd1 vssd1 vccd1 vccd1 input7/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5886 hold5886/A vssd1 vssd1 vccd1 vccd1 data_out[7] sky130_fd_sc_hd__buf_12
Xhold5897 output98/X vssd1 vssd1 vccd1 vccd1 data_out[4] sky130_fd_sc_hd__buf_12
Xhold172 hold606/X vssd1 vssd1 vccd1 vccd1 hold172/X sky130_fd_sc_hd__buf_4
Xhold183 hold13/X vssd1 vssd1 vccd1 vccd1 input12/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold194 hold194/A vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout630 _07824_/Y vssd1 vssd1 vccd1 vccd1 _15477_/A2 sky130_fd_sc_hd__buf_8
Xfanout641 _12804_/A vssd1 vssd1 vccd1 vccd1 _12753_/A sky130_fd_sc_hd__buf_4
X_09919_ hold3214/X _10013_/B _09918_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _09919_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout652 fanout739/X vssd1 vssd1 vccd1 vccd1 _12855_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_219_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout663 _13801_/C1 vssd1 vssd1 vccd1 vccd1 _12750_/A sky130_fd_sc_hd__buf_4
Xfanout674 _12289_/C1 vssd1 vssd1 vccd1 vccd1 _08115_/A sky130_fd_sc_hd__buf_4
Xfanout685 fanout689/X vssd1 vssd1 vccd1 vccd1 _13905_/A sky130_fd_sc_hd__clkbuf_4
Xfanout696 _12978_/A vssd1 vssd1 vccd1 vccd1 _14358_/A sky130_fd_sc_hd__buf_4
X_12930_ _12948_/A _12930_/B vssd1 vssd1 vccd1 vccd1 _17486_/D sky130_fd_sc_hd__and2_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _12864_/A _12861_/B vssd1 vssd1 vccd1 vccd1 _17463_/D sky130_fd_sc_hd__and2_1
XFILLER_0_217_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14600_ _15209_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14600_/X sky130_fd_sc_hd__or2_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11812_ hold4931/X _12308_/B _11811_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _11812_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _17280_/CLK _15580_/D vssd1 vssd1 vccd1 vccd1 _15580_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12792_ _12798_/A _12792_/B vssd1 vssd1 vccd1 vccd1 _17440_/D sky130_fd_sc_hd__and2_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _15103_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14531_/X sky130_fd_sc_hd__or2_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _12301_/A _11743_/B vssd1 vssd1 vccd1 vccd1 _11743_/Y sky130_fd_sc_hd__nor2_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17250_ _17250_/CLK _17250_/D vssd1 vssd1 vccd1 vccd1 _17250_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ hold3002/X _14481_/B _14461_/X _14462_/C1 vssd1 vssd1 vccd1 vccd1 _14462_/X
+ sky130_fd_sc_hd__o211a_1
X_11674_ hold4951/X _11789_/B _11673_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _11674_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16201_ _17484_/CLK _16201_/D vssd1 vssd1 vccd1 vccd1 _16201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13413_ _13722_/A _13413_/B vssd1 vssd1 vccd1 vccd1 _13413_/X sky130_fd_sc_hd__or2_1
X_10625_ _16699_/Q _10625_/B _10625_/C vssd1 vssd1 vccd1 vccd1 _10625_/X sky130_fd_sc_hd__and3_1
XFILLER_0_154_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17181_ _17277_/CLK _17181_/D vssd1 vssd1 vccd1 vccd1 _17181_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_3_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_14393_ hold338/X _14502_/B vssd1 vssd1 vccd1 vccd1 _14393_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_183_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16132_ _17331_/CLK _16132_/D vssd1 vssd1 vccd1 vccd1 _16132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10556_ hold2869/X _16676_/Q _11186_/C vssd1 vssd1 vccd1 vccd1 _10557_/B sky130_fd_sc_hd__mux2_1
X_13344_ _13794_/A _13344_/B vssd1 vssd1 vccd1 vccd1 _13344_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16063_ _16082_/CLK _16063_/D vssd1 vssd1 vccd1 vccd1 hold322/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10487_ hold2169/X hold3970/X _10595_/C vssd1 vssd1 vccd1 vccd1 _10488_/B sky130_fd_sc_hd__mux2_1
X_13275_ _13274_/X hold4390/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13275_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15014_ _15229_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _15014_/X sky130_fd_sc_hd__or2_1
XFILLER_0_121_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12226_ hold4855/X _12353_/B _12225_/X _12289_/C1 vssd1 vssd1 vccd1 vccd1 _12226_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_241_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12157_ hold5755/X _12362_/B _12156_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _12157_/X
+ sky130_fd_sc_hd__o211a_1
X_11108_ hold2086/X _16860_/Q _11204_/C vssd1 vssd1 vccd1 vccd1 _11109_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12088_ hold5237/X _12374_/B _12087_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _12088_/X
+ sky130_fd_sc_hd__o211a_1
X_16965_ _17877_/CLK _16965_/D vssd1 vssd1 vccd1 vccd1 _16965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_235_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15916_ _17291_/CLK _15916_/D vssd1 vssd1 vccd1 vccd1 hold763/A sky130_fd_sc_hd__dfxtp_1
X_11039_ hold2501/X hold4614/X _11153_/C vssd1 vssd1 vccd1 vccd1 _11040_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16896_ _18067_/CLK _16896_/D vssd1 vssd1 vccd1 vccd1 _16896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ _17738_/CLK _15847_/D vssd1 vssd1 vccd1 vccd1 _15847_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ _17728_/CLK _15778_/D vssd1 vssd1 vccd1 vccd1 _15778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17517_ _17517_/CLK _17517_/D vssd1 vssd1 vccd1 vccd1 _17517_/Q sky130_fd_sc_hd__dfxtp_1
X_14729_ hold2677/X _14720_/B _14728_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14729_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08250_ _15529_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08250_/X sky130_fd_sc_hd__or2_1
XFILLER_0_145_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17448_ _17452_/CLK _17448_/D vssd1 vssd1 vccd1 vccd1 _17448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08181_ _15515_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08181_/X sky130_fd_sc_hd__or2_1
X_17379_ _17380_/CLK _17379_/D vssd1 vssd1 vccd1 vccd1 _17379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_9_wb_clk_i clkbuf_6_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18445_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_40_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5105 _17051_/Q vssd1 vssd1 vccd1 vccd1 hold5105/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5116 _11443_/X vssd1 vssd1 vccd1 vccd1 _16971_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5127 _17009_/Q vssd1 vssd1 vccd1 vccd1 hold5127/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_275_wb_clk_i clkbuf_6_51_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18106_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_63_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5138 _16955_/Q vssd1 vssd1 vccd1 vccd1 hold5138/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4404 _13840_/Y vssd1 vssd1 vccd1 vccd1 _17733_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5149 _11458_/X vssd1 vssd1 vccd1 vccd1 _16976_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4415 _11223_/Y vssd1 vssd1 vccd1 vccd1 _11224_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4426 _13876_/Y vssd1 vssd1 vccd1 vccd1 _17745_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_204_wb_clk_i clkbuf_6_55_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18392_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4437 _10132_/X vssd1 vssd1 vccd1 vccd1 _16534_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4448 _12935_/X vssd1 vssd1 vccd1 vccd1 _12936_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3703 _11932_/X vssd1 vssd1 vccd1 vccd1 _17134_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3714 _16455_/Q vssd1 vssd1 vccd1 vccd1 hold3714/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4459 _13860_/Y vssd1 vssd1 vccd1 vccd1 _13861_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3725 _10858_/X vssd1 vssd1 vccd1 vccd1 _16776_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3736 _16451_/Q vssd1 vssd1 vccd1 vccd1 hold3736/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3747 _09709_/X vssd1 vssd1 vccd1 vccd1 _16393_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3758 _10309_/X vssd1 vssd1 vccd1 vccd1 _16593_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3769 _17431_/Q vssd1 vssd1 vccd1 vccd1 hold3769/X sky130_fd_sc_hd__dlygate4sd3_1
X_07965_ hold2828/X _07991_/A2 _07964_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _07965_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09704_ hold1399/X hold4679/X _09992_/C vssd1 vssd1 vccd1 vccd1 _09705_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07896_ _15085_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07896_/X sky130_fd_sc_hd__or2_1
XFILLER_0_207_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09635_ hold1157/X hold3620/X _10028_/C vssd1 vssd1 vccd1 vccd1 _09636_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09566_ hold2143/X _13238_/A _10067_/C vssd1 vssd1 vccd1 vccd1 _09567_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08517_ _15521_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08517_/X sky130_fd_sc_hd__or2_1
XFILLER_0_172_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09497_ hold992/A _15169_/A hold597/A _15161_/A vssd1 vssd1 vccd1 vccd1 _09498_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_0_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08448_ _08504_/A hold406/X vssd1 vssd1 vccd1 vccd1 _08448_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_92_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08379_ _08379_/A hold116/X vssd1 vssd1 vccd1 vccd1 hold117/A sky130_fd_sc_hd__and2_1
XFILLER_0_74_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10410_ _10542_/A _10410_/B vssd1 vssd1 vccd1 vccd1 _10410_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11390_ hold1809/X _16954_/Q _11783_/C vssd1 vssd1 vccd1 vccd1 _11391_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_144_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10341_ _10515_/A _10341_/B vssd1 vssd1 vccd1 vccd1 _10341_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13060_ hold5297/X _13059_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13060_/X sky130_fd_sc_hd__mux2_1
Xhold5650 _11338_/X vssd1 vssd1 vccd1 vccd1 _16936_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10272_ _10482_/A _10272_/B vssd1 vssd1 vccd1 vccd1 _10272_/X sky130_fd_sc_hd__or2_1
Xhold5661 _17052_/Q vssd1 vssd1 vccd1 vccd1 hold5661/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5672 _12043_/X vssd1 vssd1 vccd1 vccd1 _17171_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12011_ hold2373/X hold5673/X _12299_/C vssd1 vssd1 vccd1 vccd1 _12012_/B sky130_fd_sc_hd__mux2_1
Xhold5683 _17267_/Q vssd1 vssd1 vccd1 vccd1 hold5683/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5694 _11293_/X vssd1 vssd1 vccd1 vccd1 _16921_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4960 _10906_/X vssd1 vssd1 vccd1 vccd1 _16792_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4971 _12001_/X vssd1 vssd1 vccd1 vccd1 _17157_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4982 _13408_/X vssd1 vssd1 vccd1 vccd1 _17589_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4993 _16823_/Q vssd1 vssd1 vccd1 vccd1 hold4993/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout460 _13868_/C vssd1 vssd1 vccd1 vccd1 _13865_/C sky130_fd_sc_hd__clkbuf_4
Xfanout471 _12371_/C vssd1 vssd1 vccd1 vccd1 _13886_/C sky130_fd_sc_hd__clkbuf_8
X_16750_ _17985_/CLK _16750_/D vssd1 vssd1 vccd1 vccd1 _16750_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout482 _11219_/C vssd1 vssd1 vccd1 vccd1 _11789_/C sky130_fd_sc_hd__clkbuf_8
Xfanout493 _10004_/C vssd1 vssd1 vccd1 vccd1 _10028_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13962_ hold933/X _13998_/B vssd1 vssd1 vccd1 vccd1 _13962_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15701_ _17269_/CLK _15701_/D vssd1 vssd1 vccd1 vccd1 _15701_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_79_wb_clk_i clkbuf_6_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17516_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12913_ hold2633/X hold3312/X _12916_/S vssd1 vssd1 vccd1 vccd1 _12913_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_220_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16681_ _18235_/CLK _16681_/D vssd1 vssd1 vccd1 vccd1 _16681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13893_ hold307/X hold295/X vssd1 vssd1 vccd1 vccd1 hold308/A sky130_fd_sc_hd__nand2_1
XFILLER_0_213_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18420_ _18423_/CLK _18420_/D vssd1 vssd1 vccd1 vccd1 _18420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15632_ _17259_/CLK _15632_/D vssd1 vssd1 vccd1 vccd1 _15632_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ hold1614/X _17459_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12844_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_216_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _18383_/CLK _18351_/D vssd1 vssd1 vccd1 vccd1 _18351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _17899_/CLK _15563_/D vssd1 vssd1 vccd1 vccd1 _15563_/Q sky130_fd_sc_hd__dfxtp_1
X_12775_ hold2625/X _17436_/Q _12838_/S vssd1 vssd1 vccd1 vccd1 _12775_/X sky130_fd_sc_hd__mux2_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _17319_/CLK _17302_/D vssd1 vssd1 vccd1 vccd1 hold489/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_232_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14514_ hold2800/X _14537_/B _14513_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _14514_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ _18378_/CLK _18282_/D vssd1 vssd1 vccd1 vccd1 _18282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _17066_/Q _11726_/B _11726_/C vssd1 vssd1 vccd1 vccd1 _11726_/X sky130_fd_sc_hd__and3_1
XFILLER_0_16_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15494_ _15494_/A _15494_/B vssd1 vssd1 vccd1 vccd1 _18426_/D sky130_fd_sc_hd__and2_1
XFILLER_0_25_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17233_ _17266_/CLK _17233_/D vssd1 vssd1 vccd1 vccd1 _17233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14445_ _14732_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14445_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11657_ hold3061/X hold5113/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11658_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_37_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10608_ hold3488/X _10536_/A _10607_/X vssd1 vssd1 vccd1 vccd1 _10608_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17164_ _17259_/CLK _17164_/D vssd1 vssd1 vccd1 vccd1 _17164_/Q sky130_fd_sc_hd__dfxtp_1
X_14376_ _14376_/A hold787/X vssd1 vssd1 vccd1 vccd1 _17987_/D sky130_fd_sc_hd__and2_1
XFILLER_0_153_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11588_ hold2817/X hold5529/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11589_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16115_ _17338_/CLK _16115_/D vssd1 vssd1 vccd1 vccd1 hold570/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold908 hold908/A vssd1 vssd1 vccd1 vccd1 hold908/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13327_ hold5815/X _13808_/B _13326_/X _13417_/C1 vssd1 vssd1 vccd1 vccd1 _13327_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold919 hold919/A vssd1 vssd1 vccd1 vccd1 hold919/X sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ _10539_/A _10539_/B vssd1 vssd1 vccd1 vccd1 _10539_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17095_ _17127_/CLK _17095_/D vssd1 vssd1 vccd1 vccd1 _17095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16046_ _18418_/CLK _16046_/D vssd1 vssd1 vccd1 vccd1 hold515/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13258_ _17583_/Q _17117_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13258_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12209_ hold1831/X _17227_/Q _12299_/C vssd1 vssd1 vccd1 vccd1 _12210_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_0_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13189_ _13188_/X hold6001/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13189_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2309 _14199_/X vssd1 vssd1 vccd1 vccd1 _17902_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1608 _15170_/X vssd1 vssd1 vccd1 vccd1 _18368_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17997_ _17997_/CLK _17997_/D vssd1 vssd1 vccd1 vccd1 _17997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1619 _09069_/X vssd1 vssd1 vccd1 vccd1 _16149_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16948_ _17862_/CLK _16948_/D vssd1 vssd1 vccd1 vccd1 _16948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16879_ _17825_/CLK _16879_/D vssd1 vssd1 vccd1 vccd1 _16879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_232_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09420_ _09438_/B _16296_/Q vssd1 vssd1 vccd1 vccd1 _09420_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09351_ _09366_/A _09351_/B _09360_/B vssd1 vssd1 vccd1 vccd1 _09351_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08302_ hold2229/X _08336_/A2 _08301_/X _08347_/A vssd1 vssd1 vccd1 vccd1 _08302_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09282_ _12786_/A _09282_/B vssd1 vssd1 vccd1 vccd1 _16252_/D sky130_fd_sc_hd__and2_1
XFILLER_0_173_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08233_ hold1744/X _08262_/B _08232_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08233_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_456_wb_clk_i clkbuf_6_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17725_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08164_ _15515_/A hold2883/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08165_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08095_ hold2503/X _08097_/A2 _08094_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _08095_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_34_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_34_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_144_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4201 hold5907/X vssd1 vssd1 vccd1 vccd1 hold4201/X sky130_fd_sc_hd__buf_4
XFILLER_0_28_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4212 _15453_/X vssd1 vssd1 vccd1 vccd1 _15454_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4223 hold5932/X vssd1 vssd1 vccd1 vccd1 hold5933/A sky130_fd_sc_hd__buf_4
XFILLER_0_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4234 _10029_/Y vssd1 vssd1 vccd1 vccd1 _10030_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3500 _10596_/Y vssd1 vssd1 vccd1 vccd1 _10597_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4245 _16546_/Q vssd1 vssd1 vccd1 vccd1 hold4245/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4256 _10021_/Y vssd1 vssd1 vccd1 vccd1 _16497_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3511 _10041_/Y vssd1 vssd1 vccd1 vccd1 _10042_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4267 _17102_/Q vssd1 vssd1 vccd1 vccd1 hold4267/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3522 _11743_/Y vssd1 vssd1 vccd1 vccd1 _17071_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3533 _12773_/X vssd1 vssd1 vccd1 vccd1 _12774_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4278 _16739_/Q vssd1 vssd1 vccd1 vccd1 hold4278/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3544 _09856_/X vssd1 vssd1 vccd1 vccd1 _16442_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4289 _13834_/Y vssd1 vssd1 vccd1 vccd1 _17731_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3555 _09958_/X vssd1 vssd1 vccd1 vccd1 _16476_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2810 _09225_/X vssd1 vssd1 vccd1 vccd1 _16224_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3566 _16465_/Q vssd1 vssd1 vccd1 vccd1 hold3566/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2821 _17777_/Q vssd1 vssd1 vccd1 vccd1 hold2821/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3577 _09811_/X vssd1 vssd1 vccd1 vccd1 _16427_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2832 _15673_/Q vssd1 vssd1 vccd1 vccd1 hold2832/X sky130_fd_sc_hd__dlygate4sd3_1
X_08997_ hold278/X hold686/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold687/A sky130_fd_sc_hd__mux2_1
Xhold2843 _14981_/X vssd1 vssd1 vccd1 vccd1 _18276_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3588 _16507_/Q vssd1 vssd1 vccd1 vccd1 hold3588/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2854 _18233_/Q vssd1 vssd1 vccd1 vccd1 hold2854/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3599 _17362_/Q vssd1 vssd1 vccd1 vccd1 hold3599/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2865 _18207_/Q vssd1 vssd1 vccd1 vccd1 hold2865/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2876 _14947_/X vssd1 vssd1 vccd1 vccd1 _18260_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07948_ _14457_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07948_/X sky130_fd_sc_hd__or2_1
Xhold2887 _14595_/X vssd1 vssd1 vccd1 vccd1 _18091_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2898 _08304_/X vssd1 vssd1 vccd1 vccd1 _15785_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07879_ _15557_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07879_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09618_ _09912_/A _09618_/B vssd1 vssd1 vccd1 vccd1 _09618_/X sky130_fd_sc_hd__or2_1
XFILLER_0_195_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10890_ _11010_/A _10890_/B vssd1 vssd1 vccd1 vccd1 _10890_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09549_ _09933_/A _09549_/B vssd1 vssd1 vccd1 vccd1 _09549_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12560_ hold4486/X _12559_/X _12929_/S vssd1 vssd1 vccd1 vccd1 _12560_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11511_ _12174_/A _11511_/B vssd1 vssd1 vccd1 vccd1 _11511_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_197_wb_clk_i clkbuf_6_53_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18342_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_109_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12491_ hold53/X _12509_/A2 _12501_/A3 _12490_/X _12426_/A vssd1 vssd1 vccd1 vccd1
+ hold54/A sky130_fd_sc_hd__o311a_1
XFILLER_0_93_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14230_ _15521_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14230_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_126_wb_clk_i clkbuf_6_22_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16086_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_62_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11442_ _11631_/A _11442_/B vssd1 vssd1 vccd1 vccd1 _11442_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14161_ hold6072/X _14148_/B hold580/X _13897_/A vssd1 vssd1 vccd1 vccd1 hold581/A
+ sky130_fd_sc_hd__o211a_1
X_11373_ _11661_/A _11373_/B vssd1 vssd1 vccd1 vccd1 _11373_/X sky130_fd_sc_hd__or2_1
X_13112_ _13105_/X _13111_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17532_/D sky130_fd_sc_hd__o21a_1
X_10324_ hold4465/X _10628_/B _10323_/X _14697_/C1 vssd1 vssd1 vccd1 vccd1 _10324_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14092_ _15545_/A _14094_/B vssd1 vssd1 vccd1 vccd1 _14092_/Y sky130_fd_sc_hd__nand2_1
Xhold5480 _17071_/Q vssd1 vssd1 vccd1 vccd1 hold5480/X sky130_fd_sc_hd__dlygate4sd3_1
X_13043_ _17523_/Q hold907/X _17519_/Q vssd1 vssd1 vccd1 vccd1 _13043_/X sky130_fd_sc_hd__or3_1
X_10255_ hold3803/X _10619_/B _10254_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10255_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17920_ _18048_/CLK _17920_/D vssd1 vssd1 vccd1 vccd1 _17920_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5491 _13654_/X vssd1 vssd1 vccd1 vccd1 _17671_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4790 _11416_/X vssd1 vssd1 vccd1 vccd1 _16962_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17851_ _17883_/CLK _17851_/D vssd1 vssd1 vccd1 vccd1 _17851_/Q sky130_fd_sc_hd__dfxtp_1
X_10186_ hold3688/X _10568_/B _10185_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _10186_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16802_ _18061_/CLK _16802_/D vssd1 vssd1 vccd1 vccd1 _16802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17782_ _17877_/CLK _17782_/D vssd1 vssd1 vccd1 vccd1 _17782_/Q sky130_fd_sc_hd__dfxtp_1
X_14994_ _15209_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14994_/X sky130_fd_sc_hd__or2_1
XFILLER_0_233_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout290 _11100_/A vssd1 vssd1 vccd1 vccd1 _11661_/A sky130_fd_sc_hd__buf_4
XFILLER_0_234_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16733_ _17968_/CLK _16733_/D vssd1 vssd1 vccd1 vccd1 _16733_/Q sky130_fd_sc_hd__dfxtp_1
X_13945_ _15494_/A _13945_/B vssd1 vssd1 vccd1 vccd1 _17780_/D sky130_fd_sc_hd__and2_1
XFILLER_0_117_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_232_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16664_ _18226_/CLK _16664_/D vssd1 vssd1 vccd1 vccd1 _16664_/Q sky130_fd_sc_hd__dfxtp_1
X_13876_ _13888_/A _13876_/B vssd1 vssd1 vccd1 vccd1 _13876_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_186_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18403_ _18406_/CLK _18403_/D vssd1 vssd1 vccd1 vccd1 _18403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15615_ _17590_/CLK _15615_/D vssd1 vssd1 vccd1 vccd1 _15615_/Q sky130_fd_sc_hd__dfxtp_1
X_12827_ hold3377/X _12826_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12827_/X sky130_fd_sc_hd__mux2_1
X_16595_ _18177_/CLK _16595_/D vssd1 vssd1 vccd1 vccd1 _16595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_232_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18334_ _18334_/CLK _18334_/D vssd1 vssd1 vccd1 vccd1 _18334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15546_ hold2472/X _15560_/A2 _15545_/Y _12873_/A vssd1 vssd1 vccd1 vccd1 _15546_/X
+ sky130_fd_sc_hd__o211a_1
X_12758_ hold3226/X _12757_/X _12812_/S vssd1 vssd1 vccd1 vccd1 _12758_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18265_ _18265_/CLK _18265_/D vssd1 vssd1 vccd1 vccd1 _18265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11709_ _12285_/A _11709_/B vssd1 vssd1 vccd1 vccd1 _11709_/X sky130_fd_sc_hd__or2_1
XFILLER_0_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15477_ _07805_/A _15477_/A2 _09365_/B hold823/X vssd1 vssd1 vccd1 vccd1 _15480_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12689_ hold3362/X _12688_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12689_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17216_ _17280_/CLK _17216_/D vssd1 vssd1 vccd1 vccd1 _17216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14428_ hold3031/X _14433_/B _14427_/Y _14354_/A vssd1 vssd1 vccd1 vccd1 _14428_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18196_ _18228_/CLK _18196_/D vssd1 vssd1 vccd1 vccd1 _18196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17147_ _17741_/CLK _17147_/D vssd1 vssd1 vccd1 vccd1 _17147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold705 hold705/A vssd1 vssd1 vccd1 vccd1 hold705/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14359_ hold951/X hold1606/X _14381_/S vssd1 vssd1 vccd1 vccd1 _14360_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_80_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold716 hold716/A vssd1 vssd1 vccd1 vccd1 hold716/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold727 hold727/A vssd1 vssd1 vccd1 vccd1 hold727/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold738 hold738/A vssd1 vssd1 vccd1 vccd1 hold738/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold749 hold749/A vssd1 vssd1 vccd1 vccd1 hold749/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17078_ _17832_/CLK _17078_/D vssd1 vssd1 vccd1 vccd1 _17078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16029_ _17328_/CLK _16029_/D vssd1 vssd1 vccd1 vccd1 hold844/A sky130_fd_sc_hd__dfxtp_1
X_08920_ hold438/X _16078_/Q _08932_/S vssd1 vssd1 vccd1 vccd1 hold439/A sky130_fd_sc_hd__mux2_1
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2106 _07813_/X vssd1 vssd1 vccd1 vccd1 _07817_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2117 _17860_/Q vssd1 vssd1 vccd1 vccd1 hold2117/X sky130_fd_sc_hd__dlygate4sd3_1
X_08851_ _08851_/A hold774/X vssd1 vssd1 vccd1 vccd1 _16044_/D sky130_fd_sc_hd__and2_1
XFILLER_0_97_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2128 _14498_/X vssd1 vssd1 vccd1 vccd1 _18046_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2139 _17944_/Q vssd1 vssd1 vccd1 vccd1 hold2139/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1405 _08253_/X vssd1 vssd1 vccd1 vccd1 _15761_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07802_ _09339_/B _07802_/B vssd1 vssd1 vccd1 vccd1 _07802_/Y sky130_fd_sc_hd__nand2_1
Xhold1416 _17908_/Q vssd1 vssd1 vccd1 vccd1 hold1416/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1427 _15646_/Q vssd1 vssd1 vccd1 vccd1 hold1427/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08782_ _15482_/A _08782_/B vssd1 vssd1 vccd1 vccd1 _16011_/D sky130_fd_sc_hd__and2_1
Xhold1438 _15744_/Q vssd1 vssd1 vccd1 vccd1 hold1438/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1449 _14333_/X vssd1 vssd1 vccd1 vccd1 _17966_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09403_ _07785_/Y _07786_/A _11158_/A vssd1 vssd1 vccd1 vccd1 _09403_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09334_ hold1499/X _09325_/B _09333_/X _12612_/A vssd1 vssd1 vccd1 vccd1 _09334_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09265_ hold384/X hold572/X hold271/X vssd1 vssd1 vccd1 vccd1 hold573/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_290_wb_clk_i clkbuf_6_37_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18021_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_90_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08216_ hold1438/X _08213_/B _08215_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _08216_/X
+ sky130_fd_sc_hd__o211a_1
X_09196_ _15525_/A _09206_/B vssd1 vssd1 vccd1 vccd1 _09196_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08147_ _08153_/A _08147_/B vssd1 vssd1 vccd1 vccd1 _15712_/D sky130_fd_sc_hd__and2_1
XFILLER_0_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08078_ _15537_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08078_/X sky130_fd_sc_hd__or2_1
Xhold4020 _16986_/Q vssd1 vssd1 vccd1 vccd1 hold4020/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4031 _12055_/X vssd1 vssd1 vccd1 vccd1 _17175_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4042 _16420_/Q vssd1 vssd1 vccd1 vccd1 hold4042/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4053 _16809_/Q vssd1 vssd1 vccd1 vccd1 hold4053/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4064 _10927_/X vssd1 vssd1 vccd1 vccd1 _16799_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3330 _16599_/Q vssd1 vssd1 vccd1 vccd1 hold3330/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4075 _17597_/Q vssd1 vssd1 vccd1 vccd1 hold4075/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3341 _18460_/Q vssd1 vssd1 vccd1 vccd1 _07809_/B sky130_fd_sc_hd__buf_4
X_10040_ _16504_/Q _10052_/B _10040_/C vssd1 vssd1 vccd1 vccd1 _10040_/X sky130_fd_sc_hd__and3_1
Xhold4086 _10750_/X vssd1 vssd1 vccd1 vccd1 _16740_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3352 _17472_/Q vssd1 vssd1 vccd1 vccd1 hold3352/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4097 _16960_/Q vssd1 vssd1 vccd1 vccd1 hold4097/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3363 _12689_/X vssd1 vssd1 vccd1 vccd1 _12690_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3374 _12812_/X vssd1 vssd1 vccd1 vccd1 _12813_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__buf_4
XTAP_5547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2640 _13993_/X vssd1 vssd1 vccd1 vccd1 _17803_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3385 _17381_/Q vssd1 vssd1 vccd1 vccd1 hold3385/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2651 _08408_/X vssd1 vssd1 vccd1 vccd1 _15834_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3396 _17439_/Q vssd1 vssd1 vccd1 vccd1 hold3396/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2662 _15674_/Q vssd1 vssd1 vccd1 vccd1 hold2662/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold65 hold91/X vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__buf_6
XFILLER_0_216_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2673 _16214_/Q vssd1 vssd1 vccd1 vccd1 hold2673/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2684 _15522_/X vssd1 vssd1 vccd1 vccd1 _18439_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold8/X vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__buf_4
Xhold2695 _18334_/Q vssd1 vssd1 vccd1 vccd1 hold2695/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1950 _15214_/X vssd1 vssd1 vccd1 vccd1 _18389_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1961 _14929_/X vssd1 vssd1 vccd1 vccd1 _18251_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1972 _18160_/Q vssd1 vssd1 vccd1 vccd1 hold1972/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11991_ _13749_/A _11991_/B vssd1 vssd1 vccd1 vccd1 _11991_/X sky130_fd_sc_hd__or2_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1983 _09431_/X vssd1 vssd1 vccd1 vccd1 _16301_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1994 _18153_/Q vssd1 vssd1 vccd1 vccd1 hold1994/X sky130_fd_sc_hd__dlygate4sd3_1
X_13730_ hold1633/X _17697_/Q _13862_/C vssd1 vssd1 vccd1 vccd1 _13731_/B sky130_fd_sc_hd__mux2_1
X_10942_ hold5515/X _11071_/A2 _10941_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _10942_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13661_ hold1141/X hold5283/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13662_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_378_wb_clk_i clkbuf_6_33_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17584_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10873_ hold4935/X _11162_/B _10872_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _10873_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15400_ hold886/X _15448_/A2 _15446_/B1 hold724/X vssd1 vssd1 vccd1 vccd1 _15400_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12612_ _12612_/A _12612_/B vssd1 vssd1 vccd1 vccd1 _17380_/D sky130_fd_sc_hd__and2_1
X_16380_ _18389_/CLK _16380_/D vssd1 vssd1 vccd1 vccd1 _16380_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_307_wb_clk_i clkbuf_6_45_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17936_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_186_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ hold2229/X _17651_/Q _13883_/C vssd1 vssd1 vccd1 vccd1 _13593_/B sky130_fd_sc_hd__mux2_1
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15331_ _16297_/Q _15477_/A2 _15487_/B1 hold720/X _15330_/X vssd1 vssd1 vccd1 vccd1
+ _15332_/D sky130_fd_sc_hd__a221o_1
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12543_ _12948_/A _12543_/B vssd1 vssd1 vccd1 vccd1 _17357_/D sky130_fd_sc_hd__and2_1
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18050_ _18050_/CLK _18050_/D vssd1 vssd1 vccd1 vccd1 _18050_/Q sky130_fd_sc_hd__dfxtp_1
X_15262_ _15489_/A _15262_/B _15262_/C _15262_/D vssd1 vssd1 vccd1 vccd1 _15262_/X
+ sky130_fd_sc_hd__or4_1
X_12474_ _17330_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12474_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17001_ _17850_/CLK _17001_/D vssd1 vssd1 vccd1 vccd1 _17001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14213_ hold1736/X _14198_/B _14212_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _14213_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11425_ hold5637/X _12305_/B _11424_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _11425_/X
+ sky130_fd_sc_hd__o211a_1
X_15193_ _15193_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15193_/X sky130_fd_sc_hd__or2_1
XFILLER_0_22_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 _13082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14144_ _15543_/A _14148_/B vssd1 vssd1 vccd1 vccd1 _14144_/Y sky130_fd_sc_hd__nand2_1
X_11356_ hold5539/X _11165_/B _11355_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _11356_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10307_ hold2587/X _16593_/Q _10637_/C vssd1 vssd1 vccd1 vccd1 _10308_/B sky130_fd_sc_hd__mux2_1
X_14075_ hold2725/X _14107_/A2 _14074_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _14075_/X
+ sky130_fd_sc_hd__o211a_1
X_11287_ hold4887/X _11765_/B _11286_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _11287_/X
+ sky130_fd_sc_hd__o211a_1
X_13026_ hold937/X hold904/X _17519_/Q vssd1 vssd1 vccd1 vccd1 hold938/A sky130_fd_sc_hd__a21o_1
XFILLER_0_207_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_94_wb_clk_i clkbuf_6_19_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18408_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17903_ _18064_/CLK _17903_/D vssd1 vssd1 vccd1 vccd1 _17903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10238_ hold2073/X _16570_/Q _10640_/C vssd1 vssd1 vccd1 vccd1 _10239_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_218_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_wb_clk_i clkbuf_6_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17484_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_218_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10169_ hold1724/X hold3208/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10170_/B sky130_fd_sc_hd__mux2_1
X_17834_ _17834_/CLK _17834_/D vssd1 vssd1 vccd1 vccd1 _17834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_234_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14977_ hold6079/X hold447/X _14976_/X _15042_/A vssd1 vssd1 vccd1 vccd1 hold977/A
+ sky130_fd_sc_hd__o211a_1
X_17765_ _17831_/CLK _17765_/D vssd1 vssd1 vccd1 vccd1 _17765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_238_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_233_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16716_ _18307_/CLK _16716_/D vssd1 vssd1 vccd1 vccd1 _16716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13928_ hold597/A _17772_/Q hold297/X vssd1 vssd1 vccd1 vccd1 hold554/A sky130_fd_sc_hd__mux2_1
X_17696_ _17728_/CLK _17696_/D vssd1 vssd1 vccd1 vccd1 _17696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16647_ _18205_/CLK _16647_/D vssd1 vssd1 vccd1 vccd1 _16647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13859_ _17740_/Q _13883_/B _13883_/C vssd1 vssd1 vccd1 vccd1 _13859_/X sky130_fd_sc_hd__and3_1
XFILLER_0_186_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16578_ _18168_/CLK _16578_/D vssd1 vssd1 vccd1 vccd1 _16578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18317_ _18381_/CLK _18317_/D vssd1 vssd1 vccd1 vccd1 _18317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15529_ _15529_/A _15549_/B vssd1 vssd1 vccd1 vccd1 _15529_/X sky130_fd_sc_hd__or2_1
XFILLER_0_45_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09050_ hold438/X hold575/X _09060_/S vssd1 vssd1 vccd1 vccd1 _09051_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18248_ _18250_/CLK _18248_/D vssd1 vssd1 vccd1 vccd1 _18248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08001_ _14850_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08001_/X sky130_fd_sc_hd__or2_1
X_18179_ _18215_/CLK _18179_/D vssd1 vssd1 vccd1 vccd1 _18179_/Q sky130_fd_sc_hd__dfxtp_1
Xhold502 hold502/A vssd1 vssd1 vccd1 vccd1 hold502/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold513 hold513/A vssd1 vssd1 vccd1 vccd1 hold513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 hold524/A vssd1 vssd1 vccd1 vccd1 hold524/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold535 hold535/A vssd1 vssd1 vccd1 vccd1 hold535/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 hold546/A vssd1 vssd1 vccd1 vccd1 hold546/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold557 hold557/A vssd1 vssd1 vccd1 vccd1 hold557/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 hold568/A vssd1 vssd1 vccd1 vccd1 hold568/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09952_ hold3578/X _10046_/B _09951_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09952_/X
+ sky130_fd_sc_hd__o211a_1
Xhold579 hold579/A vssd1 vssd1 vccd1 vccd1 hold579/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_229_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08903_ _09440_/B hold725/X vssd1 vssd1 vccd1 vccd1 _16069_/D sky130_fd_sc_hd__and2_1
XFILLER_0_110_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09883_ hold3732/X _10049_/B _09882_/X _15228_/C1 vssd1 vssd1 vccd1 vccd1 _09883_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1202 _14051_/X vssd1 vssd1 vccd1 vccd1 _17831_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ hold180/X hold590/X _08860_/S vssd1 vssd1 vccd1 vccd1 hold591/A sky130_fd_sc_hd__mux2_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1213 _18332_/Q vssd1 vssd1 vccd1 vccd1 hold1213/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 input51/X vssd1 vssd1 vccd1 vccd1 hold1224/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1235 _18295_/Q vssd1 vssd1 vccd1 vccd1 hold1235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 _16177_/Q vssd1 vssd1 vccd1 vccd1 hold1246/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1257 _08099_/X vssd1 vssd1 vccd1 vccd1 _15689_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08765_ hold254/X hold343/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08766_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_174_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1268 _08279_/X vssd1 vssd1 vccd1 vccd1 _15774_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 _15688_/Q vssd1 vssd1 vccd1 vccd1 hold1279/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08696_ _12390_/A hold559/X vssd1 vssd1 vccd1 vccd1 _15969_/D sky130_fd_sc_hd__and2_1
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_400_wb_clk_i clkbuf_6_37_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17890_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09317_ _15539_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09317_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09248_ _12810_/A hold934/X vssd1 vssd1 vccd1 vccd1 _16235_/D sky130_fd_sc_hd__and2_1
XFILLER_0_106_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09179_ hold338/X hold363/X vssd1 vssd1 vccd1 vccd1 _09206_/B sky130_fd_sc_hd__or2_2
XFILLER_0_133_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11210_ _16894_/Q _11210_/B _11210_/C vssd1 vssd1 vccd1 vccd1 _11210_/X sky130_fd_sc_hd__and3_1
X_12190_ hold5323/X _12317_/B _12189_/X _14211_/C1 vssd1 vssd1 vccd1 vccd1 _12190_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11141_ _16871_/Q _11144_/B _11144_/C vssd1 vssd1 vccd1 vccd1 _11141_/X sky130_fd_sc_hd__and3_1
XFILLER_0_102_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput77 _13169_/A vssd1 vssd1 vccd1 vccd1 output77/X sky130_fd_sc_hd__buf_6
XTAP_6034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11072_ hold2129/X _16848_/Q _11738_/C vssd1 vssd1 vccd1 vccd1 _11073_/B sky130_fd_sc_hd__mux2_1
Xoutput88 _13249_/A vssd1 vssd1 vccd1 vccd1 output88/X sky130_fd_sc_hd__buf_6
XTAP_6045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput99 _13097_/A vssd1 vssd1 vccd1 vccd1 output99/X sky130_fd_sc_hd__buf_6
XTAP_6056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3160 _12893_/X vssd1 vssd1 vccd1 vccd1 _12894_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14900_ _14970_/A _14910_/B vssd1 vssd1 vccd1 vccd1 _14900_/X sky130_fd_sc_hd__or2_1
Xhold3171 _18325_/Q vssd1 vssd1 vccd1 vccd1 hold3171/X sky130_fd_sc_hd__dlygate4sd3_1
X_10023_ _13174_/A _09981_/A _10022_/X vssd1 vssd1 vccd1 vccd1 _10023_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3182 _18247_/Q vssd1 vssd1 vccd1 vccd1 hold3182/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15880_ _15886_/CLK _15880_/D vssd1 vssd1 vccd1 vccd1 _15880_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3193 _10014_/Y vssd1 vssd1 vccd1 vccd1 _10015_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2470 _15642_/Q vssd1 vssd1 vccd1 vccd1 hold2470/X sky130_fd_sc_hd__dlygate4sd3_1
X_14831_ hold1311/X _14826_/B _14830_/X _14893_/C1 vssd1 vssd1 vccd1 vccd1 _14831_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2481 _17876_/Q vssd1 vssd1 vccd1 vccd1 hold2481/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2492 _14583_/X vssd1 vssd1 vccd1 vccd1 _18085_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _18223_/CLK _17550_/D vssd1 vssd1 vccd1 vccd1 _17550_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1780 _14905_/X vssd1 vssd1 vccd1 vccd1 _18240_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14762_ _15209_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14762_/X sky130_fd_sc_hd__or2_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1791 _15843_/Q vssd1 vssd1 vccd1 vccd1 hold1791/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_230_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ hold4695/X _12356_/B _11973_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _11974_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16501_ _18382_/CLK _16501_/D vssd1 vssd1 vccd1 vccd1 _16501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ _13722_/A _13713_/B vssd1 vssd1 vccd1 vccd1 _13713_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10925_ hold2997/X _16799_/Q _11183_/C vssd1 vssd1 vccd1 vccd1 _10926_/B sky130_fd_sc_hd__mux2_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17481_ _17481_/CLK _17481_/D vssd1 vssd1 vccd1 vccd1 _17481_/Q sky130_fd_sc_hd__dfxtp_1
X_14693_ hold2685/X _14720_/B _14692_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14693_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16432_ _18345_/CLK _16432_/D vssd1 vssd1 vccd1 vccd1 _16432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_141_wb_clk_i clkbuf_6_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17533_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13644_ _13773_/A _13644_/B vssd1 vssd1 vccd1 vccd1 _13644_/X sky130_fd_sc_hd__or2_1
X_10856_ hold1606/X _16776_/Q _11144_/C vssd1 vssd1 vccd1 vccd1 _10857_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _17533_/CLK _16363_/D vssd1 vssd1 vccd1 vccd1 _16363_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _13794_/A _13575_/B vssd1 vssd1 vccd1 vccd1 _13575_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10787_ hold2701/X hold4575/X _11171_/C vssd1 vssd1 vccd1 vccd1 _10788_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18102_ _18192_/CLK _18102_/D vssd1 vssd1 vccd1 vccd1 _18102_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _15314_/A _15314_/B vssd1 vssd1 vccd1 vccd1 _18407_/D sky130_fd_sc_hd__and2_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ _17515_/Q _17353_/Q _12985_/S vssd1 vssd1 vccd1 vccd1 _12526_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_109_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16294_ _18408_/CLK _16294_/D vssd1 vssd1 vccd1 vccd1 _16294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18033_ _18065_/CLK _18033_/D vssd1 vssd1 vccd1 vccd1 _18033_/Q sky130_fd_sc_hd__dfxtp_1
X_15245_ hold873/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15245_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12457_ hold147/X _12509_/A2 _12501_/A3 _12456_/X _12410_/A vssd1 vssd1 vccd1 vccd1
+ hold148/A sky130_fd_sc_hd__o311a_1
XFILLER_0_125_1306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11408_ hold2209/X hold4097/X _12335_/C vssd1 vssd1 vccd1 vccd1 _11409_/B sky130_fd_sc_hd__mux2_1
X_15176_ hold2819/X _15167_/B _15175_/X _15176_/C1 vssd1 vssd1 vccd1 vccd1 _15176_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_1414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12388_ _15344_/A hold848/X vssd1 vssd1 vccd1 vccd1 _17287_/D sky130_fd_sc_hd__and2_1
XFILLER_0_111_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14127_ hold2607/X _14148_/B _14126_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _14127_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_239_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11339_ hold2627/X _16937_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _11340_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14058_ hold915/X _14106_/B vssd1 vssd1 vccd1 vccd1 _14058_/X sky130_fd_sc_hd__or2_1
XFILLER_0_219_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13009_ _14972_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13009_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17817_ _17850_/CLK _17817_/D vssd1 vssd1 vccd1 vccd1 _17817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_234_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08550_ hold673/X hold849/X _08592_/S vssd1 vssd1 vccd1 vccd1 hold850/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_229_wb_clk_i clkbuf_6_63_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18099_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17748_ _17748_/CLK _17748_/D vssd1 vssd1 vccd1 vccd1 _17748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08481_ hold1720/X _08486_/B _08480_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _08481_/X
+ sky130_fd_sc_hd__o211a_1
X_17679_ _17744_/CLK _17679_/D vssd1 vssd1 vccd1 vccd1 _17679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09102_ _15543_/A _09102_/B vssd1 vssd1 vccd1 vccd1 _09102_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_210_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09033_ _15254_/A hold658/X vssd1 vssd1 vccd1 vccd1 _16133_/D sky130_fd_sc_hd__and2_1
XFILLER_0_116_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_241_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold310 hold310/A vssd1 vssd1 vccd1 vccd1 hold310/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 hold321/A vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold332 hold332/A vssd1 vssd1 vccd1 vccd1 hold332/X sky130_fd_sc_hd__buf_8
Xhold343 hold343/A vssd1 vssd1 vccd1 vccd1 hold343/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold354 hold354/A vssd1 vssd1 vccd1 vccd1 hold354/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold365 hold365/A vssd1 vssd1 vccd1 vccd1 hold365/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold376 hold629/X vssd1 vssd1 vccd1 vccd1 hold630/A sky130_fd_sc_hd__buf_6
Xhold387 hold387/A vssd1 vssd1 vccd1 vccd1 hold387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 hold398/A vssd1 vssd1 vccd1 vccd1 hold398/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 _15019_/C1 vssd1 vssd1 vccd1 vccd1 _15226_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_110_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09935_ hold3108/X hold4711/X _10031_/C vssd1 vssd1 vccd1 vccd1 _09936_/B sky130_fd_sc_hd__mux2_1
Xfanout812 fanout816/X vssd1 vssd1 vccd1 vccd1 _15228_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout823 _14863_/C1 vssd1 vssd1 vccd1 vccd1 _10564_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout834 _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14857_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_141_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout845 _13864_/A vssd1 vssd1 vccd1 vccd1 _12301_/A sky130_fd_sc_hd__buf_8
XFILLER_0_99_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout856 _17754_/Q vssd1 vssd1 vccd1 vccd1 _11218_/A sky130_fd_sc_hd__buf_8
X_09866_ hold1374/X hold3660/X _10040_/C vssd1 vssd1 vccd1 vccd1 _09867_/B sky130_fd_sc_hd__mux2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout867 _15217_/A vssd1 vssd1 vccd1 vccd1 _15163_/A sky130_fd_sc_hd__clkbuf_16
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout878 hold950/X vssd1 vssd1 vccd1 vccd1 hold951/A sky130_fd_sc_hd__buf_6
Xhold1010 _17858_/Q vssd1 vssd1 vccd1 vccd1 hold1010/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 input48/X vssd1 vssd1 vccd1 vccd1 hold914/A sky130_fd_sc_hd__buf_1
XFILLER_0_176_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout889 hold423/X vssd1 vssd1 vccd1 vccd1 _15519_/A sky130_fd_sc_hd__clkbuf_16
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08817_ _15364_/A _08817_/B vssd1 vssd1 vccd1 vccd1 _16027_/D sky130_fd_sc_hd__and2_1
Xhold1032 _15086_/X vssd1 vssd1 vccd1 vccd1 _18327_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1043 _15861_/Q vssd1 vssd1 vccd1 vccd1 hold1043/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ hold1789/X _16423_/Q _10004_/C vssd1 vssd1 vccd1 vccd1 _09798_/B sky130_fd_sc_hd__mux2_1
Xhold1054 _15801_/Q vssd1 vssd1 vccd1 vccd1 hold1054/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1065 _14829_/X vssd1 vssd1 vccd1 vccd1 _18204_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1076 hold1076/A vssd1 vssd1 vccd1 vccd1 _15207_/A sky130_fd_sc_hd__buf_12
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _15414_/A _08748_/B vssd1 vssd1 vccd1 vccd1 _15994_/D sky130_fd_sc_hd__and2_1
Xhold1087 _18438_/Q vssd1 vssd1 vccd1 vccd1 hold1087/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1098 _15809_/Q vssd1 vssd1 vccd1 vccd1 hold1098/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ hold679/X hold851/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold852/A sky130_fd_sc_hd__mux2_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _11088_/A _10710_/B vssd1 vssd1 vccd1 vccd1 _10710_/X sky130_fd_sc_hd__or2_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11690_ hold2308/X hold5257/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11691_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_165_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10641_ hold3459/X _10554_/A _10640_/X vssd1 vssd1 vccd1 vccd1 _10641_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13360_ hold5357/X _13856_/B _13359_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _13360_/X
+ sky130_fd_sc_hd__o211a_1
X_10572_ hold3475/X _10560_/A _10571_/X vssd1 vssd1 vccd1 vccd1 _10573_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_183_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12311_ _12311_/A _12353_/B _13409_/S vssd1 vssd1 vccd1 vccd1 _12311_/X sky130_fd_sc_hd__and3_1
XFILLER_0_161_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13291_ _13290_/X _16929_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13291_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_107_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15030_ _15030_/A _15030_/B vssd1 vssd1 vccd1 vccd1 _18300_/D sky130_fd_sc_hd__and2_1
XFILLER_0_122_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12242_ hold2410/X _17238_/Q _12242_/S vssd1 vssd1 vccd1 vccd1 _12243_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12173_ hold2703/X _17215_/Q _12173_/S vssd1 vssd1 vccd1 vccd1 _12174_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11124_ _11124_/A _11124_/B vssd1 vssd1 vccd1 vccd1 _11124_/X sky130_fd_sc_hd__or2_1
X_16981_ _17831_/CLK _16981_/D vssd1 vssd1 vccd1 vccd1 _16981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15932_ _17325_/CLK _15932_/D vssd1 vssd1 vccd1 vccd1 hold302/A sky130_fd_sc_hd__dfxtp_1
XTAP_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11055_ _11631_/A _11055_/B vssd1 vssd1 vccd1 vccd1 _11055_/X sky130_fd_sc_hd__or2_1
XTAP_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10006_ _11203_/A _10006_/B vssd1 vssd1 vccd1 vccd1 _10006_/Y sky130_fd_sc_hd__nor2_1
XTAP_5174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15863_ _17672_/CLK _15863_/D vssd1 vssd1 vccd1 vccd1 _15863_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_393_wb_clk_i clkbuf_6_36_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17902_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_235_1323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14814_ _15099_/A _14830_/B vssd1 vssd1 vccd1 vccd1 _14814_/X sky130_fd_sc_hd__or2_1
XFILLER_0_203_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17602_ _17730_/CLK _17602_/D vssd1 vssd1 vccd1 vccd1 _17602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15794_ _17661_/CLK _15794_/D vssd1 vssd1 vccd1 vccd1 _15794_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_322_wb_clk_i clkbuf_6_46_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17904_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_192_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ _17533_/CLK _17533_/D vssd1 vssd1 vccd1 vccd1 _17533_/Q sky130_fd_sc_hd__dfxtp_1
X_14745_ hold2485/X _14772_/B _14744_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _14745_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ hold1287/X hold4011/X _12371_/C vssd1 vssd1 vccd1 vccd1 _11958_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_203_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17464_ _17464_/CLK _17464_/D vssd1 vssd1 vccd1 vccd1 _17464_/Q sky130_fd_sc_hd__dfxtp_1
X_10908_ _11661_/A _10908_/B vssd1 vssd1 vccd1 vccd1 _10908_/X sky130_fd_sc_hd__or2_1
X_14676_ _15231_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14676_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11888_ hold1217/X hold4332/X _13886_/C vssd1 vssd1 vccd1 vccd1 _11889_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16415_ _18296_/CLK _16415_/D vssd1 vssd1 vccd1 vccd1 _16415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13627_ hold5024/X _13817_/B _13626_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _13627_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17395_ _18452_/CLK _17395_/D vssd1 vssd1 vccd1 vccd1 _17395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10839_ _11694_/A _10839_/B vssd1 vssd1 vccd1 vccd1 _10839_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16346_ _18361_/CLK _16346_/D vssd1 vssd1 vccd1 vccd1 _16346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13558_ hold5628/X _13880_/B _13557_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _13558_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12509_ hold68/X _12509_/A2 _08868_/X _12508_/X _09061_/A vssd1 vssd1 vccd1 vccd1
+ hold69/A sky130_fd_sc_hd__o311a_1
XFILLER_0_140_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16277_ _17378_/CLK _16277_/D vssd1 vssd1 vccd1 vccd1 _16277_/Q sky130_fd_sc_hd__dfxtp_1
X_13489_ hold5150/X _13871_/B _13488_/X _13675_/C1 vssd1 vssd1 vccd1 vccd1 _13489_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5309 _17023_/Q vssd1 vssd1 vccd1 vccd1 hold5309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15228_ hold2675/X _15219_/B _15227_/X _15228_/C1 vssd1 vssd1 vccd1 vccd1 _15228_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18016_ _18016_/CLK _18016_/D vssd1 vssd1 vccd1 vccd1 _18016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4608 _17598_/Q vssd1 vssd1 vccd1 vccd1 hold4608/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4619 _09739_/X vssd1 vssd1 vccd1 vccd1 _16403_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15159_ _15213_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15159_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3907 _16593_/Q vssd1 vssd1 vccd1 vccd1 hold3907/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3918 _10741_/X vssd1 vssd1 vccd1 vccd1 _16737_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3929 _11071_/X vssd1 vssd1 vccd1 vccd1 _16847_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07981_ hold1817/X _07991_/A2 _07980_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _07981_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_201_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_238_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09720_ _09948_/A _09720_/B vssd1 vssd1 vccd1 vccd1 _09720_/X sky130_fd_sc_hd__or2_1
X_09651_ _09957_/A _09651_/B vssd1 vssd1 vccd1 vccd1 _09651_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08602_ _12418_/A hold768/X vssd1 vssd1 vccd1 vccd1 _15923_/D sky130_fd_sc_hd__and2_1
X_09582_ _10482_/A _09582_/B vssd1 vssd1 vccd1 vccd1 _09582_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08533_ _09057_/A hold227/X vssd1 vssd1 vccd1 vccd1 _15890_/D sky130_fd_sc_hd__and2_1
XFILLER_0_72_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08464_ _14517_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08464_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08395_ _14164_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08395_/X sky130_fd_sc_hd__or2_1
XFILLER_0_18_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09016_ hold452/X hold876/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09017_/B sky130_fd_sc_hd__mux2_1
Xhold5810 _13720_/X vssd1 vssd1 vccd1 vccd1 _17693_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5821 _16430_/Q vssd1 vssd1 vccd1 vccd1 hold5821/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5832 _09544_/X vssd1 vssd1 vccd1 vccd1 _16338_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5843 hold6005/X vssd1 vssd1 vccd1 vccd1 _13177_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5854 output92/X vssd1 vssd1 vccd1 vccd1 data_out[28] sky130_fd_sc_hd__buf_12
XFILLER_0_103_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold140 hold140/A vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5865 hold6018/X vssd1 vssd1 vccd1 vccd1 _13257_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5876 hold5876/A vssd1 vssd1 vccd1 vccd1 data_out[6] sky130_fd_sc_hd__buf_12
Xhold151 hold151/A vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 input7/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5887 hold6028/X vssd1 vssd1 vccd1 vccd1 _13121_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 hold173/A vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5898 hold6032/X vssd1 vssd1 vccd1 vccd1 _13097_/A sky130_fd_sc_hd__buf_1
Xhold184 input12/X vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__buf_1
Xhold195 hold28/X vssd1 vssd1 vccd1 vccd1 input33/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout620 _09351_/Y vssd1 vssd1 vccd1 vccd1 _15448_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_217_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout631 _07824_/Y vssd1 vssd1 vccd1 vccd1 _09362_/A sky130_fd_sc_hd__clkbuf_4
X_09918_ _11061_/A _09918_/B vssd1 vssd1 vccd1 vccd1 _09918_/X sky130_fd_sc_hd__or2_1
Xfanout642 _12804_/A vssd1 vssd1 vccd1 vccd1 _12738_/A sky130_fd_sc_hd__buf_4
Xfanout653 _12597_/A vssd1 vssd1 vccd1 vccd1 _12924_/A sky130_fd_sc_hd__buf_4
Xfanout664 _13801_/C1 vssd1 vssd1 vccd1 vccd1 _13417_/C1 sky130_fd_sc_hd__buf_2
XFILLER_0_176_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout675 _12289_/C1 vssd1 vssd1 vccd1 vccd1 _08137_/A sky130_fd_sc_hd__buf_4
Xfanout686 _14376_/A vssd1 vssd1 vccd1 vccd1 _14352_/A sky130_fd_sc_hd__buf_4
Xfanout697 _12978_/A vssd1 vssd1 vccd1 vccd1 _14362_/A sky130_fd_sc_hd__buf_4
X_09849_ _11109_/A _09849_/B vssd1 vssd1 vccd1 vccd1 _09849_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ hold3360/X _12859_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12861_/B sky130_fd_sc_hd__mux2_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _13797_/A _11811_/B vssd1 vssd1 vccd1 vccd1 _11811_/X sky130_fd_sc_hd__or2_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12791_ hold3534/X _12790_/X _12839_/S vssd1 vssd1 vccd1 vccd1 _12791_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ hold1684/X _14537_/B _14529_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _14530_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11742_ hold3520/X _12219_/A _11741_/X vssd1 vssd1 vccd1 vccd1 _11742_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_230_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _14461_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14461_/X sky130_fd_sc_hd__or2_1
XFILLER_0_113_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11694_/A _11673_/B vssd1 vssd1 vccd1 vccd1 _11673_/X sky130_fd_sc_hd__or2_1
XFILLER_0_154_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16200_ _17484_/CLK _16200_/D vssd1 vssd1 vccd1 vccd1 _16200_/Q sky130_fd_sc_hd__dfxtp_1
X_13412_ hold2043/X hold4781/X _13796_/S vssd1 vssd1 vccd1 vccd1 _13413_/B sky130_fd_sc_hd__mux2_1
X_10624_ _10651_/A _10624_/B vssd1 vssd1 vccd1 vccd1 _16698_/D sky130_fd_sc_hd__nor2_1
X_17180_ _17262_/CLK _17180_/D vssd1 vssd1 vccd1 vccd1 _17180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14392_ _14392_/A _14392_/B vssd1 vssd1 vccd1 vccd1 _17995_/D sky130_fd_sc_hd__and2_1
XFILLER_0_14_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16131_ _17325_/CLK _16131_/D vssd1 vssd1 vccd1 vccd1 hold644/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13343_ hold2826/X hold4262/X _13862_/C vssd1 vssd1 vccd1 vccd1 _13344_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_106_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10555_ hold3347/X _10649_/B _10554_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10555_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16062_ _17293_/CLK _16062_/D vssd1 vssd1 vccd1 vccd1 hold825/A sky130_fd_sc_hd__dfxtp_1
X_13274_ _17585_/Q _17119_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13274_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_224_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ hold3634/X _10625_/B _10485_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _10486_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15013_ hold2699/X _15004_/B _15012_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _15013_/X
+ sky130_fd_sc_hd__o211a_1
X_12225_ _13314_/A _12225_/B vssd1 vssd1 vccd1 vccd1 _12225_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_1322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12156_ _12267_/A _12156_/B vssd1 vssd1 vccd1 vccd1 _12156_/X sky130_fd_sc_hd__or2_1
XFILLER_0_235_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11107_ hold3718/X _11201_/B _11106_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _11107_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12087_ _13749_/A _12087_/B vssd1 vssd1 vccd1 vccd1 _12087_/X sky130_fd_sc_hd__or2_1
X_16964_ _17856_/CLK _16964_/D vssd1 vssd1 vccd1 vccd1 _16964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15915_ _16082_/CLK _15915_/D vssd1 vssd1 vccd1 vccd1 hold470/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11038_ hold4099/X _11071_/A2 _11037_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _11038_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16895_ _18066_/CLK _16895_/D vssd1 vssd1 vccd1 vccd1 _16895_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _17747_/CLK _15846_/D vssd1 vssd1 vccd1 vccd1 _15846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ hold4598/X _12988_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12989_/X sky130_fd_sc_hd__mux2_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15777_ _17734_/CLK _15777_/D vssd1 vssd1 vccd1 vccd1 _15777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17516_ _17516_/CLK _17516_/D vssd1 vssd1 vccd1 vccd1 _17516_/Q sky130_fd_sc_hd__dfxtp_1
X_14728_ _15229_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14728_/X sky130_fd_sc_hd__or2_1
XFILLER_0_185_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14659_ hold2019/X _14666_/B _14658_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _14659_/X
+ sky130_fd_sc_hd__o211a_1
X_17447_ _17450_/CLK _17447_/D vssd1 vssd1 vccd1 vccd1 _17447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08180_ hold1633/X _08209_/B _08179_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _08180_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17378_ _17378_/CLK _17378_/D vssd1 vssd1 vccd1 vccd1 _17378_/Q sky130_fd_sc_hd__dfxtp_1
X_16329_ _18240_/CLK _16329_/D vssd1 vssd1 vccd1 vccd1 _16329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_6_24_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_24_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_28_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5106 _11587_/X vssd1 vssd1 vccd1 vccd1 _17019_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5117 _17148_/Q vssd1 vssd1 vccd1 vccd1 hold5117/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5128 _11461_/X vssd1 vssd1 vccd1 vccd1 _16977_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5139 _11299_/X vssd1 vssd1 vccd1 vccd1 _16923_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4405 _16924_/Q vssd1 vssd1 vccd1 vccd1 hold4405/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4416 _11224_/Y vssd1 vssd1 vccd1 vccd1 _16898_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4427 _16928_/Q vssd1 vssd1 vccd1 vccd1 hold4427/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4438 _17105_/Q vssd1 vssd1 vccd1 vccd1 hold4438/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4449 _16926_/Q vssd1 vssd1 vccd1 vccd1 hold4449/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3704 _16903_/Q vssd1 vssd1 vccd1 vccd1 hold3704/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3715 _09799_/X vssd1 vssd1 vccd1 vccd1 _16423_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3726 _16374_/Q vssd1 vssd1 vccd1 vccd1 hold3726/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3737 _09787_/X vssd1 vssd1 vccd1 vccd1 _16419_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3748 _17505_/Q vssd1 vssd1 vccd1 vccd1 hold3748/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3759 _17494_/Q vssd1 vssd1 vccd1 vccd1 hold3759/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_244_wb_clk_i clkbuf_6_57_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18188_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07964_ _15533_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07964_/X sky130_fd_sc_hd__or2_1
XFILLER_0_215_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09703_ hold3777/X _10004_/B _09702_/X _08954_/A vssd1 vssd1 vccd1 vccd1 _09703_/X
+ sky130_fd_sc_hd__o211a_1
X_07895_ hold2431/X _07918_/B _07894_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _07895_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09634_ hold4801/X _11171_/B _09633_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _09634_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09565_ hold3245/X _10049_/B _09564_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09565_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_1226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08516_ hold1376/X _08503_/Y _08515_/X _13417_/C1 vssd1 vssd1 vccd1 vccd1 _08516_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09496_ _09496_/A hold820/A _15173_/A vssd1 vssd1 vccd1 vccd1 _09498_/C sky130_fd_sc_hd__or3b_1
XFILLER_0_66_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_63_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_63_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_148_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08447_ hold405/A hold509/A hold337/A hold444/A vssd1 vssd1 vccd1 vccd1 hold406/A
+ sky130_fd_sc_hd__or4bb_2
XFILLER_0_149_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08378_ hold97/X _15821_/Q hold115/X vssd1 vssd1 vccd1 vccd1 hold116/A sky130_fd_sc_hd__mux2_1
XFILLER_0_74_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10340_ hold3045/X hold4456/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10341_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5640 _11257_/X vssd1 vssd1 vccd1 vccd1 _16909_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10271_ hold2773/X hold3550/X _10601_/C vssd1 vssd1 vccd1 vccd1 _10272_/B sky130_fd_sc_hd__mux2_1
Xhold5651 _17064_/Q vssd1 vssd1 vccd1 vccd1 hold5651/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5662 _11590_/X vssd1 vssd1 vccd1 vccd1 _17020_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5673 _17161_/Q vssd1 vssd1 vccd1 vccd1 hold5673/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12010_ hold4851/X _13811_/B _12009_/X _08363_/A vssd1 vssd1 vccd1 vccd1 _12010_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5684 _12235_/X vssd1 vssd1 vccd1 vccd1 _17235_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4950 _10804_/X vssd1 vssd1 vccd1 vccd1 _16758_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5695 _17171_/Q vssd1 vssd1 vccd1 vccd1 hold5695/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4961 _16949_/Q vssd1 vssd1 vccd1 vccd1 hold4961/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4972 _16811_/Q vssd1 vssd1 vccd1 vccd1 hold4972/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4983 _17263_/Q vssd1 vssd1 vccd1 vccd1 hold4983/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4994 _10903_/X vssd1 vssd1 vccd1 vccd1 _16791_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout450 _11723_/C vssd1 vssd1 vccd1 vccd1 _11726_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_205_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout461 _13868_/C vssd1 vssd1 vccd1 vccd1 _13841_/C sky130_fd_sc_hd__buf_6
XFILLER_0_156_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout472 fanout485/X vssd1 vssd1 vccd1 vccd1 _12371_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_1259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13961_ hold2788/X _13995_/A2 _13960_/X _13895_/A vssd1 vssd1 vccd1 vccd1 _13961_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout483 _11219_/C vssd1 vssd1 vccd1 vccd1 _11765_/C sky130_fd_sc_hd__clkbuf_8
Xfanout494 _10964_/S vssd1 vssd1 vccd1 vccd1 _10004_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_226_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15700_ _17268_/CLK _15700_/D vssd1 vssd1 vccd1 vccd1 _15700_/Q sky130_fd_sc_hd__dfxtp_1
X_12912_ _12924_/A _12912_/B vssd1 vssd1 vccd1 vccd1 _17480_/D sky130_fd_sc_hd__and2_1
X_16680_ _18265_/CLK _16680_/D vssd1 vssd1 vccd1 vccd1 _16680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13892_ hold361/A hold268/X vssd1 vssd1 vccd1 vccd1 _14163_/B sky130_fd_sc_hd__or2_4
XFILLER_0_119_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12843_ _12843_/A _12843_/B vssd1 vssd1 vccd1 vccd1 _17457_/D sky130_fd_sc_hd__and2_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15631_ _18430_/CLK _15631_/D vssd1 vssd1 vccd1 vccd1 _15631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18350_ _18382_/CLK _18350_/D vssd1 vssd1 vccd1 vccd1 _18350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15562_ _17900_/CLK _15562_/D vssd1 vssd1 vccd1 vccd1 _15562_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12774_ _12777_/A _12774_/B vssd1 vssd1 vccd1 vccd1 _17434_/D sky130_fd_sc_hd__and2_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _17301_/CLK _17301_/D vssd1 vssd1 vccd1 vccd1 hold540/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14513_ _15193_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14513_/X sky130_fd_sc_hd__or2_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_48_wb_clk_i clkbuf_6_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18073_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11725_ _12301_/A _11725_/B vssd1 vssd1 vccd1 vccd1 _17065_/D sky130_fd_sc_hd__nor2_1
X_18281_ _18315_/CLK _18281_/D vssd1 vssd1 vccd1 vccd1 _18281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15493_ _14164_/A hold1813/X _15505_/S vssd1 vssd1 vccd1 vccd1 _15493_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_232_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14444_ hold1342/X _14446_/A2 _14443_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _14444_/X
+ sky130_fd_sc_hd__o211a_1
X_17232_ _17264_/CLK _17232_/D vssd1 vssd1 vccd1 vccd1 _17232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11656_ hold5135/X _11165_/B _11655_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _11656_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10607_ _16693_/Q _10631_/B _10637_/C vssd1 vssd1 vccd1 vccd1 _10607_/X sky130_fd_sc_hd__and3_1
XFILLER_0_142_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17163_ _17878_/CLK _17163_/D vssd1 vssd1 vccd1 vccd1 _17163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14375_ hold597/X hold786/X _14381_/S vssd1 vssd1 vccd1 vccd1 hold787/A sky130_fd_sc_hd__mux2_1
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11587_ hold5105/X _12317_/B _11586_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11587_/X
+ sky130_fd_sc_hd__o211a_1
X_16114_ _17337_/CLK _16114_/D vssd1 vssd1 vccd1 vccd1 hold502/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13326_ _13719_/A _13326_/B vssd1 vssd1 vccd1 vccd1 _13326_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10538_ hold1095/X _16670_/Q _10538_/S vssd1 vssd1 vccd1 vccd1 _10539_/B sky130_fd_sc_hd__mux2_1
Xhold909 hold909/A vssd1 vssd1 vccd1 vccd1 hold909/X sky130_fd_sc_hd__dlygate4sd3_1
X_17094_ _17222_/CLK _17094_/D vssd1 vssd1 vccd1 vccd1 _17094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16045_ _17301_/CLK _16045_/D vssd1 vssd1 vccd1 vccd1 hold624/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13257_ _13257_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13257_/X sky130_fd_sc_hd__and2_1
X_10469_ hold1311/X _16647_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10470_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_122_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_237_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12208_ hold5125/X _12293_/B _12207_/X _12822_/A vssd1 vssd1 vccd1 vccd1 _12208_/X
+ sky130_fd_sc_hd__o211a_1
X_13188_ hold4350/X _13187_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13188_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_236_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12139_ hold5675/X _11771_/B _12138_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _12139_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17996_ _18028_/CLK _17996_/D vssd1 vssd1 vccd1 vccd1 _17996_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1609 _18272_/Q vssd1 vssd1 vccd1 vccd1 hold1609/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16947_ _18065_/CLK _16947_/D vssd1 vssd1 vccd1 vccd1 _16947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16878_ _18049_/CLK _16878_/D vssd1 vssd1 vccd1 vccd1 _16878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15829_ _17624_/CLK _15829_/D vssd1 vssd1 vccd1 vccd1 _15829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09350_ _15543_/A _15541_/A _15182_/A _09352_/D vssd1 vssd1 vccd1 vccd1 _09360_/B
+ sky130_fd_sc_hd__or4_1
X_08301_ _15145_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08301_/X sky130_fd_sc_hd__or2_1
XFILLER_0_158_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09281_ _15557_/A hold973/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09282_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_173_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08232_ hold915/X _08280_/B vssd1 vssd1 vccd1 vccd1 _08232_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08163_ _08163_/A _08163_/B vssd1 vssd1 vccd1 vccd1 _15719_/D sky130_fd_sc_hd__and2_1
XFILLER_0_160_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08094_ _15553_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08094_/X sky130_fd_sc_hd__or2_1
XFILLER_0_113_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4202 _15243_/X vssd1 vssd1 vccd1 vccd1 _15244_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4213 hold5917/X vssd1 vssd1 vccd1 vccd1 hold5918/A sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_425_wb_clk_i clkbuf_6_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17741_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4224 _15383_/X vssd1 vssd1 vccd1 vccd1 _15384_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4235 _10030_/Y vssd1 vssd1 vccd1 vccd1 _16500_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3501 _16525_/Q vssd1 vssd1 vccd1 vccd1 hold3501/X sky130_fd_sc_hd__buf_2
XFILLER_0_11_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4246 _10647_/Y vssd1 vssd1 vccd1 vccd1 _10648_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4257 hold5964/X vssd1 vssd1 vccd1 vccd1 hold5965/A sky130_fd_sc_hd__buf_4
Xhold3512 _16734_/Q vssd1 vssd1 vccd1 vccd1 hold3512/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3523 _16720_/Q vssd1 vssd1 vccd1 vccd1 hold3523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4268 _12315_/Y vssd1 vssd1 vccd1 vccd1 _12316_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4279 _11226_/Y vssd1 vssd1 vccd1 vccd1 _11227_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3534 _17440_/Q vssd1 vssd1 vccd1 vccd1 hold3534/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3545 _16381_/Q vssd1 vssd1 vccd1 vccd1 hold3545/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2800 _18053_/Q vssd1 vssd1 vccd1 vccd1 hold2800/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2811 _15671_/Q vssd1 vssd1 vccd1 vccd1 hold2811/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3556 _16622_/Q vssd1 vssd1 vccd1 vccd1 hold3556/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3567 _09829_/X vssd1 vssd1 vccd1 vccd1 _16433_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08996_ _12426_/A _08996_/B vssd1 vssd1 vccd1 vccd1 _16115_/D sky130_fd_sc_hd__and2_1
Xhold2822 _15734_/Q vssd1 vssd1 vccd1 vccd1 hold2822/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3578 _16506_/Q vssd1 vssd1 vccd1 vccd1 hold3578/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2833 _08067_/X vssd1 vssd1 vccd1 vccd1 _15673_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3589 _09955_/X vssd1 vssd1 vccd1 vccd1 _16475_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2844 _17881_/Q vssd1 vssd1 vccd1 vccd1 hold2844/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2855 _14889_/X vssd1 vssd1 vccd1 vccd1 _18233_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2866 _14835_/X vssd1 vssd1 vccd1 vccd1 _18207_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07947_ hold2691/X _07991_/A2 _07946_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _07947_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2877 _15668_/Q vssd1 vssd1 vccd1 vccd1 hold2877/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2888 _18195_/Q vssd1 vssd1 vccd1 vccd1 hold2888/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2899 _15860_/Q vssd1 vssd1 vccd1 vccd1 hold2899/X sky130_fd_sc_hd__dlygate4sd3_1
X_07878_ hold1356/X _07865_/B _07877_/X _14211_/C1 vssd1 vssd1 vccd1 vccd1 _07878_/X
+ sky130_fd_sc_hd__o211a_1
X_09617_ hold2842/X hold3564/X _10025_/C vssd1 vssd1 vccd1 vccd1 _09618_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_190_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09548_ hold3065/X _13190_/A _10028_/C vssd1 vssd1 vccd1 vccd1 _09549_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09479_ _09483_/B _09483_/C vssd1 vssd1 vccd1 vccd1 _09481_/C sky130_fd_sc_hd__or2_1
XFILLER_0_135_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11510_ hold2725/X hold4789/X _12173_/S vssd1 vssd1 vccd1 vccd1 _11511_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12490_ _17338_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12490_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11441_ hold2960/X _16971_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _11442_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14160_ hold579/X _14160_/B vssd1 vssd1 vccd1 vccd1 hold580/A sky130_fd_sc_hd__or2_1
XFILLER_0_61_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11372_ hold2131/X _16948_/Q _11660_/S vssd1 vssd1 vccd1 vccd1 _11373_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13111_ _13199_/A1 _13109_/X _13110_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13111_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_21_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10323_ _10515_/A _10323_/B vssd1 vssd1 vccd1 vccd1 _10323_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14091_ hold2871/X _14094_/B _14090_/Y _15506_/A vssd1 vssd1 vccd1 vccd1 _14091_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_166_wb_clk_i clkbuf_6_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18377_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_219_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13042_ _13046_/C _13046_/D hold922/X vssd1 vssd1 vccd1 vccd1 hold923/A sky130_fd_sc_hd__nor3_1
Xhold5470 _17612_/Q vssd1 vssd1 vccd1 vccd1 hold5470/X sky130_fd_sc_hd__dlygate4sd3_1
X_10254_ _10524_/A _10254_/B vssd1 vssd1 vccd1 vccd1 _10254_/X sky130_fd_sc_hd__or2_1
Xhold5481 _11647_/X vssd1 vssd1 vccd1 vccd1 _17039_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5492 _17743_/Q vssd1 vssd1 vccd1 vccd1 hold5492/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4780 _13633_/X vssd1 vssd1 vccd1 vccd1 _17664_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_56_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17850_ _17850_/CLK _17850_/D vssd1 vssd1 vccd1 vccd1 _17850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10185_ _10476_/A _10185_/B vssd1 vssd1 vccd1 vccd1 _10185_/X sky130_fd_sc_hd__or2_1
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4791 _17200_/Q vssd1 vssd1 vccd1 vccd1 hold4791/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16801_ _18036_/CLK _16801_/D vssd1 vssd1 vccd1 vccd1 _16801_/Q sky130_fd_sc_hd__dfxtp_1
X_17781_ _18427_/CLK _17781_/D vssd1 vssd1 vccd1 vccd1 _17781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14993_ hold1157/X _15004_/B _14992_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _14993_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout280 _13599_/A vssd1 vssd1 vccd1 vccd1 _13758_/A sky130_fd_sc_hd__buf_2
Xfanout291 fanout299/X vssd1 vssd1 vccd1 vccd1 _11100_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16732_ _18031_/CLK _16732_/D vssd1 vssd1 vccd1 vccd1 _16732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13944_ _15559_/A hold1238/X hold297/X vssd1 vssd1 vccd1 vccd1 _13945_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_202_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16663_ _18221_/CLK _16663_/D vssd1 vssd1 vccd1 vccd1 _16663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13875_ hold4424/X _13758_/A _13874_/X vssd1 vssd1 vccd1 vccd1 _13875_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18402_ _18409_/CLK _18402_/D vssd1 vssd1 vccd1 vccd1 _18402_/Q sky130_fd_sc_hd__dfxtp_1
X_15614_ _17268_/CLK _15614_/D vssd1 vssd1 vccd1 vccd1 _15614_/Q sky130_fd_sc_hd__dfxtp_1
X_12826_ hold2557/X _17453_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12826_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_186_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16594_ _18124_/CLK _16594_/D vssd1 vssd1 vccd1 vccd1 _16594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18333_ _18379_/CLK _18333_/D vssd1 vssd1 vccd1 vccd1 _18333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12757_ hold2330/X _17430_/Q _12811_/S vssd1 vssd1 vccd1 vccd1 _12757_/X sky130_fd_sc_hd__mux2_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15545_ _15545_/A _15547_/B vssd1 vssd1 vccd1 vccd1 _15545_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_155_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11708_ hold1416/X hold5199/X _12317_/C vssd1 vssd1 vccd1 vccd1 _11709_/B sky130_fd_sc_hd__mux2_1
X_18264_ _18296_/CLK hold241/X vssd1 vssd1 vccd1 vccd1 _18264_/Q sky130_fd_sc_hd__dfxtp_1
X_15476_ hold347/X _09392_/B _09386_/D hold542/X _15475_/X vssd1 vssd1 vccd1 vccd1
+ _15480_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_56_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12688_ hold1643/X _17407_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12688_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_127_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14427_ _15541_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _14427_/Y sky130_fd_sc_hd__nand2_1
X_17215_ _17247_/CLK _17215_/D vssd1 vssd1 vccd1 vccd1 _17215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11639_ hold2215/X hold5577/X _11738_/C vssd1 vssd1 vccd1 vccd1 _11640_/B sky130_fd_sc_hd__mux2_1
X_18195_ _18221_/CLK _18195_/D vssd1 vssd1 vccd1 vccd1 _18195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14358_ _14358_/A _14358_/B vssd1 vssd1 vccd1 vccd1 _17978_/D sky130_fd_sc_hd__and2_1
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17146_ _17576_/CLK _17146_/D vssd1 vssd1 vccd1 vccd1 _17146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold706 hold706/A vssd1 vssd1 vccd1 vccd1 hold706/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 hold717/A vssd1 vssd1 vccd1 vccd1 hold717/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13309_ _13308_/X hold3208/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13309_/X sky130_fd_sc_hd__mux2_1
Xhold728 hold728/A vssd1 vssd1 vccd1 vccd1 hold728/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17077_ _17861_/CLK _17077_/D vssd1 vssd1 vccd1 vccd1 _17077_/Q sky130_fd_sc_hd__dfxtp_1
Xhold739 hold739/A vssd1 vssd1 vccd1 vccd1 hold739/X sky130_fd_sc_hd__buf_1
XFILLER_0_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14289_ hold2139/X _14333_/A2 _14288_/X _14354_/A vssd1 vssd1 vccd1 vccd1 _14289_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16028_ _17284_/CLK _16028_/D vssd1 vssd1 vccd1 vccd1 hold837/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08850_ hold92/X hold773/X _08866_/S vssd1 vssd1 vccd1 vccd1 hold774/A sky130_fd_sc_hd__mux2_1
Xhold2107 _09366_/A vssd1 vssd1 vccd1 vccd1 _09400_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2118 _14113_/X vssd1 vssd1 vccd1 vccd1 _17860_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2129 _18051_/Q vssd1 vssd1 vccd1 vccd1 hold2129/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07801_ _09342_/A _07801_/B vssd1 vssd1 vccd1 vccd1 _07802_/B sky130_fd_sc_hd__and2_1
Xhold1406 _17990_/Q vssd1 vssd1 vccd1 vccd1 hold1406/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08781_ hold438/X hold458/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08782_/B sky130_fd_sc_hd__mux2_1
Xhold1417 _14211_/X vssd1 vssd1 vccd1 vccd1 _17908_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17979_ _17981_/CLK _17979_/D vssd1 vssd1 vccd1 vccd1 _17979_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1428 _08010_/X vssd1 vssd1 vccd1 vccd1 _15646_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1439 _08216_/X vssd1 vssd1 vccd1 vccd1 _15744_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_237_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09402_ _12412_/A _09402_/B vssd1 vssd1 vccd1 vccd1 _16286_/D sky130_fd_sc_hd__and2_1
XFILLER_0_153_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09333_ _15555_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09333_/X sky130_fd_sc_hd__or2_1
XFILLER_0_177_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09264_ _12750_/A _09264_/B vssd1 vssd1 vccd1 vccd1 _16243_/D sky130_fd_sc_hd__and2_1
XFILLER_0_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08215_ _15549_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08215_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09195_ hold986/X _09218_/B _09194_/X _12798_/A vssd1 vssd1 vccd1 vccd1 hold987/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08146_ _14330_/A hold1217/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08147_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222_1303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08077_ hold1275/X _08088_/B _08076_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _08077_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4010 _10384_/X vssd1 vssd1 vccd1 vccd1 _16618_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4021 _11392_/X vssd1 vssd1 vccd1 vccd1 _16954_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_222_1347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4032 _17175_/Q vssd1 vssd1 vccd1 vccd1 hold4032/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4043 _09694_/X vssd1 vssd1 vccd1 vccd1 _16388_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4054 _16632_/Q vssd1 vssd1 vccd1 vccd1 hold4054/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3320 _16591_/Q vssd1 vssd1 vccd1 vccd1 hold3320/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4065 _17436_/Q vssd1 vssd1 vccd1 vccd1 hold4065/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3331 _10231_/X vssd1 vssd1 vccd1 vccd1 _16567_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4076 _13336_/X vssd1 vssd1 vccd1 vccd1 _17565_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3342 _09391_/X vssd1 vssd1 vccd1 vccd1 _16283_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4087 _17039_/Q vssd1 vssd1 vccd1 vccd1 hold4087/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3353 _17464_/Q vssd1 vssd1 vccd1 vccd1 hold3353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4098 _11314_/X vssd1 vssd1 vccd1 vccd1 _16928_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3364 _17480_/Q vssd1 vssd1 vccd1 vccd1 hold3364/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__buf_4
XFILLER_0_216_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2630 _14432_/X vssd1 vssd1 vccd1 vccd1 _18014_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3375 _17390_/Q vssd1 vssd1 vccd1 vccd1 hold3375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2641 _18353_/Q vssd1 vssd1 vccd1 vccd1 hold2641/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3386 _12614_/X vssd1 vssd1 vccd1 vccd1 _12615_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__buf_4
XTAP_5559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08979_ hold53/X hold753/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08980_/B sky130_fd_sc_hd__mux2_1
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2652 _18104_/Q vssd1 vssd1 vccd1 vccd1 hold2652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3397 _12788_/X vssd1 vssd1 vccd1 vccd1 _12789_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2663 _08069_/X vssd1 vssd1 vccd1 vccd1 _15674_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2674 _09205_/X vssd1 vssd1 vccd1 vccd1 _16214_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2685 _18138_/Q vssd1 vssd1 vccd1 vccd1 hold2685/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1940 _14239_/X vssd1 vssd1 vccd1 vccd1 _17920_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__clkbuf_4
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1951 _18069_/Q vssd1 vssd1 vccd1 vccd1 hold1951/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2696 _15100_/X vssd1 vssd1 vccd1 vccd1 _18334_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ hold2470/X _17154_/Q _13748_/S vssd1 vssd1 vccd1 vccd1 _11991_/B sky130_fd_sc_hd__mux2_1
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1962 _17887_/Q vssd1 vssd1 vccd1 vccd1 hold1962/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1973 _14739_/X vssd1 vssd1 vccd1 vccd1 _18160_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1984 _18096_/Q vssd1 vssd1 vccd1 vccd1 hold1984/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1995 _14723_/X vssd1 vssd1 vccd1 vccd1 _18153_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10941_ _11655_/A _10941_/B vssd1 vssd1 vccd1 vccd1 _10941_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13660_ hold5608/X _13880_/B _13659_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13660_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10872_ _11067_/A _10872_/B vssd1 vssd1 vccd1 vccd1 _10872_/X sky130_fd_sc_hd__or2_1
XFILLER_0_97_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ hold3268/X _12610_/X _12923_/S vssd1 vssd1 vccd1 vccd1 _12611_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ hold5504/X _13880_/B _13590_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _17650_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15330_ hold473/X _15448_/A2 _15446_/B1 hold825/X vssd1 vssd1 vccd1 vccd1 _15330_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ hold4517/X _12541_/X _12929_/S vssd1 vssd1 vccd1 vccd1 _12542_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_213_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15261_ _16290_/Q _15477_/A2 _15487_/B1 _16078_/Q _15260_/X vssd1 vssd1 vccd1 vccd1
+ _15262_/D sky130_fd_sc_hd__a221o_1
X_12473_ hold59/X _12445_/A _12445_/B _12472_/X _12394_/A vssd1 vssd1 vccd1 vccd1
+ hold60/A sky130_fd_sc_hd__o311a_1
XFILLER_0_191_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_347_wb_clk_i clkbuf_6_42_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17747_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17000_ _17847_/CLK _17000_/D vssd1 vssd1 vccd1 vccd1 _17000_/Q sky130_fd_sc_hd__dfxtp_1
X_14212_ _15557_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14212_/X sky130_fd_sc_hd__or2_1
X_11424_ _12093_/A _11424_/B vssd1 vssd1 vccd1 vccd1 _11424_/X sky130_fd_sc_hd__or2_1
X_15192_ hold2349/X _15219_/B _15191_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _15192_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_8 _13100_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14143_ hold3039/X _14142_/B _14142_/Y _14143_/C1 vssd1 vssd1 vccd1 vccd1 _14143_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11355_ _11556_/A _11355_/B vssd1 vssd1 vccd1 vccd1 _11355_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10306_ hold3753/X _10598_/B _10305_/X _15218_/C1 vssd1 vssd1 vccd1 vccd1 _10306_/X
+ sky130_fd_sc_hd__o211a_1
X_14074_ _14413_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14074_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11286_ _11670_/A _11286_/B vssd1 vssd1 vccd1 vccd1 _11286_/X sky130_fd_sc_hd__or2_1
X_13025_ hold905/X _13025_/B _13025_/C vssd1 vssd1 vccd1 vccd1 _17518_/D sky130_fd_sc_hd__and3_1
XFILLER_0_219_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17902_ _17902_/CLK _17902_/D vssd1 vssd1 vccd1 vccd1 _17902_/Q sky130_fd_sc_hd__dfxtp_1
X_10237_ hold3272/X _10637_/B _10236_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10237_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_238_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17833_ _17894_/CLK _17833_/D vssd1 vssd1 vccd1 vccd1 _17833_/Q sky130_fd_sc_hd__dfxtp_1
X_10168_ hold4543/X _10628_/B _10167_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _10168_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_234_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_233_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_238_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17764_ _17894_/CLK _17764_/D vssd1 vssd1 vccd1 vccd1 _17764_/Q sky130_fd_sc_hd__dfxtp_1
X_10099_ hold3247/X _10577_/B _10098_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _10099_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_221_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14976_ hold945/X _15018_/B vssd1 vssd1 vccd1 vccd1 _14976_/X sky130_fd_sc_hd__or2_1
XFILLER_0_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_63_wb_clk_i clkbuf_6_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18047_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16715_ _18072_/CLK _16715_/D vssd1 vssd1 vccd1 vccd1 _16715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13927_ _13927_/A hold385/X vssd1 vssd1 vccd1 vccd1 _17771_/D sky130_fd_sc_hd__and2_1
XFILLER_0_221_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17695_ _17730_/CLK _17695_/D vssd1 vssd1 vccd1 vccd1 _17695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16646_ _18172_/CLK _16646_/D vssd1 vssd1 vccd1 vccd1 _16646_/Q sky130_fd_sc_hd__dfxtp_1
X_13858_ _13873_/A _13858_/B vssd1 vssd1 vccd1 vccd1 _13858_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_201_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12809_ hold3230/X _12808_/X _12839_/S vssd1 vssd1 vccd1 vccd1 _12809_/X sky130_fd_sc_hd__mux2_1
X_16577_ _18232_/CLK _16577_/D vssd1 vssd1 vccd1 vccd1 _16577_/Q sky130_fd_sc_hd__dfxtp_1
X_13789_ hold5545/X _13883_/B _13788_/X _08347_/A vssd1 vssd1 vccd1 vccd1 _13789_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18316_ _18372_/CLK _18316_/D vssd1 vssd1 vccd1 vccd1 _18316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15528_ hold1350/X _15547_/B _15527_/X _12849_/A vssd1 vssd1 vccd1 vccd1 _15528_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18247_ _18375_/CLK _18247_/D vssd1 vssd1 vccd1 vccd1 _18247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15459_ hold732/X _09386_/A _09357_/A _17321_/Q _15458_/X vssd1 vssd1 vccd1 vccd1
+ _15462_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_127_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08000_ hold1966/X _08033_/B _07999_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _08000_/X
+ sky130_fd_sc_hd__o211a_1
X_18178_ _18188_/CLK _18178_/D vssd1 vssd1 vccd1 vccd1 _18178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold503 hold503/A vssd1 vssd1 vccd1 vccd1 hold503/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 hold514/A vssd1 vssd1 vccd1 vccd1 hold514/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17129_ _17161_/CLK _17129_/D vssd1 vssd1 vccd1 vccd1 _17129_/Q sky130_fd_sc_hd__dfxtp_1
Xhold525 hold525/A vssd1 vssd1 vccd1 vccd1 hold525/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold536 hold536/A vssd1 vssd1 vccd1 vccd1 hold536/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 hold547/A vssd1 vssd1 vccd1 vccd1 hold547/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09951_ _09978_/A _09951_/B vssd1 vssd1 vccd1 vccd1 _09951_/X sky130_fd_sc_hd__or2_1
Xhold558 hold558/A vssd1 vssd1 vccd1 vccd1 hold558/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 hold569/A vssd1 vssd1 vccd1 vccd1 hold569/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08902_ hold185/X hold724/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold725/A sky130_fd_sc_hd__mux2_1
XFILLER_0_141_1378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09882_ _09954_/A _09882_/B vssd1 vssd1 vccd1 vccd1 _09882_/X sky130_fd_sc_hd__or2_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _15314_/A _08833_/B vssd1 vssd1 vccd1 vccd1 _16035_/D sky130_fd_sc_hd__and2_1
XFILLER_0_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 _15787_/Q vssd1 vssd1 vccd1 vccd1 hold1203/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 _15096_/X vssd1 vssd1 vccd1 vccd1 _18332_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1225 _09332_/X vssd1 vssd1 vccd1 vccd1 _16276_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1236 _15019_/X vssd1 vssd1 vccd1 vccd1 _18295_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08764_ _15414_/A hold564/X vssd1 vssd1 vccd1 vccd1 _16002_/D sky130_fd_sc_hd__and2_1
Xhold1247 _09129_/X vssd1 vssd1 vccd1 vccd1 _16177_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1258 _17844_/Q vssd1 vssd1 vccd1 vccd1 hold1258/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1269 _16229_/Q vssd1 vssd1 vccd1 vccd1 hold1269/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08695_ hold180/X hold558/X _08721_/S vssd1 vssd1 vccd1 vccd1 hold559/A sky130_fd_sc_hd__mux2_1
XFILLER_0_95_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09316_ hold2145/X _09323_/B _09315_/X _12588_/A vssd1 vssd1 vccd1 vccd1 _09316_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09247_ hold933/X _16235_/Q _09283_/S vssd1 vssd1 vccd1 vccd1 hold934/A sky130_fd_sc_hd__mux2_1
XFILLER_0_7_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_440_wb_clk_i clkbuf_6_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17561_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_91_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09178_ hold338/X hold363/X vssd1 vssd1 vccd1 vccd1 _09178_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_44_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08129_ _08145_/A _08129_/B vssd1 vssd1 vccd1 vccd1 _15703_/D sky130_fd_sc_hd__and2_1
XFILLER_0_82_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11140_ hold4079/X _11732_/B _11139_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _11140_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput78 _13177_/A vssd1 vssd1 vccd1 vccd1 output78/X sky130_fd_sc_hd__buf_6
XTAP_6035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11071_ _11165_/A _11071_/A2 _11070_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _11071_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput89 _13257_/A vssd1 vssd1 vccd1 vccd1 output89/X sky130_fd_sc_hd__buf_6
XTAP_5312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3150 _12851_/X vssd1 vssd1 vccd1 vccd1 _12852_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10022_ _16498_/Q _10022_/B _10022_/C vssd1 vssd1 vccd1 vccd1 _10022_/X sky130_fd_sc_hd__and3_1
Xhold3161 _17422_/Q vssd1 vssd1 vccd1 vccd1 hold3161/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3172 _15082_/X vssd1 vssd1 vccd1 vccd1 _18325_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3183 _14921_/X vssd1 vssd1 vccd1 vccd1 _18247_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3194 _10015_/Y vssd1 vssd1 vccd1 vccd1 _16495_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2460 _17878_/Q vssd1 vssd1 vccd1 vccd1 hold2460/X sky130_fd_sc_hd__dlygate4sd3_1
X_14830_ _15169_/A _14830_/B vssd1 vssd1 vccd1 vccd1 _14830_/X sky130_fd_sc_hd__or2_1
XTAP_5378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2471 _08002_/X vssd1 vssd1 vccd1 vccd1 _15642_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2482 _14145_/X vssd1 vssd1 vccd1 vccd1 _17876_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2493 _18164_/Q vssd1 vssd1 vccd1 vccd1 hold2493/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1770 _15776_/Q vssd1 vssd1 vccd1 vccd1 hold1770/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1781 _18179_/Q vssd1 vssd1 vccd1 vccd1 hold1781/X sky130_fd_sc_hd__dlygate4sd3_1
X_14761_ hold2867/X _14772_/B _14760_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14761_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11973_ _13482_/A _11973_/B vssd1 vssd1 vccd1 vccd1 _11973_/X sky130_fd_sc_hd__or2_1
XFILLER_0_203_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1792 _08426_/X vssd1 vssd1 vccd1 vccd1 _15843_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16500_ _18381_/CLK _16500_/D vssd1 vssd1 vccd1 vccd1 _16500_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10924_ hold4147/X _11753_/B _10923_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _10924_/X
+ sky130_fd_sc_hd__o211a_1
X_13712_ hold2589/X hold4660/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13713_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_196_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14692_ _15193_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14692_/X sky130_fd_sc_hd__or2_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17480_ _17481_/CLK _17480_/D vssd1 vssd1 vccd1 vccd1 _17480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16431_ _18376_/CLK _16431_/D vssd1 vssd1 vccd1 vccd1 _16431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10855_ hold3850/X _11144_/B _10854_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _10855_/X
+ sky130_fd_sc_hd__o211a_1
X_13643_ hold1054/X _17668_/Q _13871_/C vssd1 vssd1 vccd1 vccd1 _13644_/B sky130_fd_sc_hd__mux2_1
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16362_ _18371_/CLK _16362_/D vssd1 vssd1 vccd1 vccd1 _16362_/Q sky130_fd_sc_hd__dfxtp_1
X_13574_ hold2971/X _17645_/Q _13766_/S vssd1 vssd1 vccd1 vccd1 _13575_/B sky130_fd_sc_hd__mux2_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ hold4138/X _11744_/B _10785_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _10786_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18101_ _18191_/CLK _18101_/D vssd1 vssd1 vccd1 vccd1 _18101_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15313_ _15490_/A1 _15305_/X _15312_/X _15481_/B1 hold4199/X vssd1 vssd1 vccd1 vccd1
+ _15313_/X sky130_fd_sc_hd__a32o_1
X_12525_ _12984_/A _12525_/B vssd1 vssd1 vccd1 vccd1 _17351_/D sky130_fd_sc_hd__and2_1
XFILLER_0_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16293_ _18404_/CLK _16293_/D vssd1 vssd1 vccd1 vccd1 _16293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_181_wb_clk_i clkbuf_6_51_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18389_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18032_ _18059_/CLK _18032_/D vssd1 vssd1 vccd1 vccd1 _18032_/Q sky130_fd_sc_hd__dfxtp_1
X_12456_ _17321_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12456_/X sky130_fd_sc_hd__or2_1
X_15244_ _15244_/A _15244_/B vssd1 vssd1 vccd1 vccd1 _18400_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_110_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17336_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ hold5313/X _11789_/B _11406_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _11407_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15175_ _15229_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15175_/X sky130_fd_sc_hd__or2_1
X_12387_ hold684/X hold847/X _12441_/S vssd1 vssd1 vccd1 vccd1 hold848/A sky130_fd_sc_hd__mux2_1
XFILLER_0_105_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14126_ _15525_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14126_/X sky130_fd_sc_hd__or2_1
X_11338_ hold5649/X _11717_/B _11337_/X _12588_/A vssd1 vssd1 vccd1 vccd1 _11338_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_238_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14057_ hold2090/X _14107_/A2 _14056_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _14057_/X
+ sky130_fd_sc_hd__o211a_1
X_11269_ hold5537/X _12323_/B _11268_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11269_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13008_ hold1811/X _13003_/Y _13007_/X _12984_/A vssd1 vssd1 vccd1 vccd1 _13008_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17816_ _18429_/CLK _17816_/D vssd1 vssd1 vccd1 vccd1 _17816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_238_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_234_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17747_ _17747_/CLK _17747_/D vssd1 vssd1 vccd1 vccd1 _17747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14959_ hold2838/X _14946_/B _14958_/X _15228_/C1 vssd1 vssd1 vccd1 vccd1 _14959_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08480_ _14604_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08480_/X sky130_fd_sc_hd__or2_1
XFILLER_0_221_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17678_ _17678_/CLK _17678_/D vssd1 vssd1 vccd1 vccd1 _17678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16629_ _18233_/CLK _16629_/D vssd1 vssd1 vccd1 vccd1 _16629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_269_wb_clk_i clkbuf_6_57_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18162_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_186_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09101_ hold2830/X _09102_/B _09100_/Y _12978_/A vssd1 vssd1 vccd1 vccd1 _09101_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09032_ hold185/X hold657/X _09056_/S vssd1 vssd1 vccd1 vccd1 hold658/A sky130_fd_sc_hd__mux2_1
XFILLER_0_25_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold300 hold300/A vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold311 hold311/A vssd1 vssd1 vccd1 vccd1 hold311/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold322 hold322/A vssd1 vssd1 vccd1 vccd1 hold322/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold333 hold333/A vssd1 vssd1 vccd1 vccd1 hold333/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold344 hold344/A vssd1 vssd1 vccd1 vccd1 hold344/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold355 hold355/A vssd1 vssd1 vccd1 vccd1 hold355/X sky130_fd_sc_hd__buf_4
Xhold366 hold929/X vssd1 vssd1 vccd1 vccd1 hold930/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 hold377/A vssd1 vssd1 vccd1 vccd1 hold377/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold388 hold388/A vssd1 vssd1 vccd1 vccd1 hold388/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout802 _15019_/C1 vssd1 vssd1 vccd1 vccd1 _15218_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_141_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold399 hold399/A vssd1 vssd1 vccd1 vccd1 hold399/X sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ hold4648/X _10028_/B _09933_/X _15048_/A vssd1 vssd1 vccd1 vccd1 _09934_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout813 _15204_/C1 vssd1 vssd1 vccd1 vccd1 _15212_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout824 _14390_/A vssd1 vssd1 vccd1 vccd1 _14344_/A sky130_fd_sc_hd__buf_4
Xfanout835 _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14853_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_176_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout846 _17754_/Q vssd1 vssd1 vccd1 vccd1 _13864_/A sky130_fd_sc_hd__buf_8
X_09865_ hold3652/X _10049_/B _09864_/X _15212_/C1 vssd1 vssd1 vccd1 vccd1 _09865_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout857 _13312_/B1 vssd1 vssd1 vccd1 vccd1 _13048_/A sky130_fd_sc_hd__buf_6
Xhold1000 _18263_/Q vssd1 vssd1 vccd1 vccd1 hold1000/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout868 _07782_/Y vssd1 vssd1 vccd1 vccd1 _15217_/A sky130_fd_sc_hd__buf_8
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout879 _15145_/A vssd1 vssd1 vccd1 vccd1 _15525_/A sky130_fd_sc_hd__buf_12
Xhold1011 _14107_/X vssd1 vssd1 vccd1 vccd1 _17858_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1022 hold914/X vssd1 vssd1 vccd1 vccd1 hold1022/X sky130_fd_sc_hd__buf_8
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ hold29/X hold440/X _08866_/S vssd1 vssd1 vccd1 vccd1 _08817_/B sky130_fd_sc_hd__mux2_1
Xhold1033 _18178_/Q vssd1 vssd1 vccd1 vccd1 hold1033/X sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ hold5177/X _09992_/B _09795_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _09796_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1044 _08465_/X vssd1 vssd1 vccd1 vccd1 _15861_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1055 _08336_/X vssd1 vssd1 vccd1 vccd1 _15801_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 _15822_/Q vssd1 vssd1 vccd1 vccd1 hold1066/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08747_ hold452/X hold873/X _08779_/S vssd1 vssd1 vccd1 vccd1 _08748_/B sky130_fd_sc_hd__mux2_1
Xhold1077 _13918_/X vssd1 vssd1 vccd1 vccd1 _13919_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1088 _15520_/X vssd1 vssd1 vccd1 vccd1 _18438_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1099 _15731_/Q vssd1 vssd1 vccd1 vccd1 hold1099/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08678_ _15434_/A _08678_/B vssd1 vssd1 vccd1 vccd1 _15960_/D sky130_fd_sc_hd__and2_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ _16704_/Q _10649_/B _10640_/C vssd1 vssd1 vccd1 vccd1 _10640_/X sky130_fd_sc_hd__and3_1
XFILLER_0_53_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10571_ _10571_/A _10571_/B _10571_/C vssd1 vssd1 vccd1 vccd1 _10571_/X sky130_fd_sc_hd__and3_1
XFILLER_0_91_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12310_ _13819_/A _12310_/B vssd1 vssd1 vccd1 vccd1 _12310_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_134_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13290_ _17587_/Q _17121_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13290_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12241_ hold5384/X _12335_/B _12240_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _12241_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12172_ hold5771/X _12362_/B _12171_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _12172_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11123_ hold1127/X hold3858/X _11219_/C vssd1 vssd1 vccd1 vccd1 _11124_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16980_ _17862_/CLK _16980_/D vssd1 vssd1 vccd1 vccd1 _16980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15931_ _16090_/CLK _15931_/D vssd1 vssd1 vccd1 vccd1 hold859/A sky130_fd_sc_hd__dfxtp_1
XTAP_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11054_ hold878/X hold5569/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11055_/B sky130_fd_sc_hd__mux2_1
XTAP_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10005_ _13126_/A _09984_/A _10004_/X vssd1 vssd1 vccd1 vccd1 _10005_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15862_ _17739_/CLK _15862_/D vssd1 vssd1 vccd1 vccd1 _15862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2290 _09189_/X vssd1 vssd1 vccd1 vccd1 _16206_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17601_ _17729_/CLK _17601_/D vssd1 vssd1 vccd1 vccd1 _17601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14813_ hold1495/X _14828_/B _14812_/X _14895_/C1 vssd1 vssd1 vccd1 vccd1 _14813_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ _17724_/CLK _15793_/D vssd1 vssd1 vccd1 vccd1 _15793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17532_ _17533_/CLK _17532_/D vssd1 vssd1 vccd1 vccd1 _17532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14744_ _15191_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14744_/X sky130_fd_sc_hd__or2_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ hold4863/X _11771_/B _11955_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _11956_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17463_ _17464_/CLK _17463_/D vssd1 vssd1 vccd1 vccd1 _17463_/Q sky130_fd_sc_hd__dfxtp_1
X_10907_ hold1927/X hold5335/X _11660_/S vssd1 vssd1 vccd1 vccd1 _10908_/B sky130_fd_sc_hd__mux2_1
X_14675_ hold2643/X _14666_/B _14674_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14675_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_362_wb_clk_i clkbuf_6_35_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17608_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11887_ hold5121/X _11798_/B _11886_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11887_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16414_ _18327_/CLK _16414_/D vssd1 vssd1 vccd1 vccd1 _16414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13626_ _13722_/A _13626_/B vssd1 vssd1 vccd1 vccd1 _13626_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10838_ hold3191/X hold4117/X _11789_/C vssd1 vssd1 vccd1 vccd1 _10839_/B sky130_fd_sc_hd__mux2_1
X_17394_ _18452_/CLK _17394_/D vssd1 vssd1 vccd1 vccd1 _17394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16345_ _18352_/CLK _16345_/D vssd1 vssd1 vccd1 vccd1 _16345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10769_ hold2908/X _16747_/Q _11153_/C vssd1 vssd1 vccd1 vccd1 _10770_/B sky130_fd_sc_hd__mux2_1
X_13557_ _13599_/A _13557_/B vssd1 vssd1 vccd1 vccd1 _13557_/X sky130_fd_sc_hd__or2_1
XFILLER_0_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12508_ _17347_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12508_/X sky130_fd_sc_hd__or2_1
Xclkbuf_6_14_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_14_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_125_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13488_ _13776_/A _13488_/B vssd1 vssd1 vccd1 vccd1 _13488_/X sky130_fd_sc_hd__or2_1
X_16276_ _17380_/CLK _16276_/D vssd1 vssd1 vccd1 vccd1 _16276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18015_ _18047_/CLK _18015_/D vssd1 vssd1 vccd1 vccd1 _18015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12439_ hold495/X hold695/X _12441_/S vssd1 vssd1 vccd1 vccd1 hold696/A sky130_fd_sc_hd__mux2_1
X_15227_ _15227_/A _15227_/B vssd1 vssd1 vccd1 vccd1 _15227_/X sky130_fd_sc_hd__or2_1
XFILLER_0_152_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4609 _13339_/X vssd1 vssd1 vccd1 vccd1 _17566_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15158_ hold6064/X _15165_/B hold631/X _15024_/A vssd1 vssd1 vccd1 vccd1 hold632/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3908 _10213_/X vssd1 vssd1 vccd1 vccd1 _16561_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3919 _16897_/Q vssd1 vssd1 vccd1 vccd1 hold3919/X sky130_fd_sc_hd__dlygate4sd3_1
X_14109_ _14789_/A _14163_/B vssd1 vssd1 vccd1 vccd1 _14140_/B sky130_fd_sc_hd__or2_4
X_15089_ _15197_/A _15119_/B vssd1 vssd1 vccd1 vccd1 _15089_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07980_ _15549_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07980_/X sky130_fd_sc_hd__or2_1
XFILLER_0_227_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09650_ hold2009/X hold3726/X _10040_/C vssd1 vssd1 vccd1 vccd1 _09651_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_207_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08601_ hold618/X hold767/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold768/A sky130_fd_sc_hd__mux2_1
XFILLER_0_222_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09581_ _18264_/Q _13278_/A _10601_/C vssd1 vssd1 vccd1 vccd1 _09582_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_222_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08532_ hold226/X _15890_/Q _08594_/S vssd1 vssd1 vccd1 vccd1 hold227/A sky130_fd_sc_hd__mux2_1
XFILLER_0_54_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_53_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_53_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_188_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08463_ hold2899/X _08488_/B _08462_/X _13675_/C1 vssd1 vssd1 vccd1 vccd1 _08463_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08394_ _08504_/A hold445/X vssd1 vssd1 vccd1 vccd1 _08445_/B sky130_fd_sc_hd__or2_4
XFILLER_0_147_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09015_ _15434_/A hold756/X vssd1 vssd1 vccd1 vccd1 _16124_/D sky130_fd_sc_hd__and2_1
XFILLER_0_143_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5800 _11872_/X vssd1 vssd1 vccd1 vccd1 _17114_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5811 _16324_/Q vssd1 vssd1 vccd1 vccd1 _13062_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5822 _09724_/X vssd1 vssd1 vccd1 vccd1 _16398_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5833 _16502_/Q vssd1 vssd1 vccd1 vccd1 hold5833/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5844 output78/X vssd1 vssd1 vccd1 vccd1 data_out[15] sky130_fd_sc_hd__buf_12
Xhold130 input27/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 hold16/X vssd1 vssd1 vccd1 vccd1 input21/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5855 hold6011/X vssd1 vssd1 vccd1 vccd1 _13169_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5866 output89/X vssd1 vssd1 vccd1 vccd1 data_out[25] sky130_fd_sc_hd__buf_12
Xhold5877 hold6023/X vssd1 vssd1 vccd1 vccd1 _13217_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold152 hold152/A vssd1 vssd1 vccd1 vccd1 hold152/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5888 hold5888/A vssd1 vssd1 vccd1 vccd1 data_out[8] sky130_fd_sc_hd__buf_12
XFILLER_0_229_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold163 hold2/X vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__clkbuf_8
Xhold5899 output99/X vssd1 vssd1 vccd1 vccd1 data_out[5] sky130_fd_sc_hd__buf_12
Xhold174 hold174/A vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold185 hold14/X vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__buf_4
XFILLER_0_106_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold196 input33/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 _15485_/B1 vssd1 vssd1 vccd1 vccd1 _09362_/D sky130_fd_sc_hd__buf_6
Xfanout621 _09351_/Y vssd1 vssd1 vccd1 vccd1 _09367_/A sky130_fd_sc_hd__clkbuf_8
Xfanout632 _12445_/A vssd1 vssd1 vccd1 vccd1 _12509_/A2 sky130_fd_sc_hd__clkbuf_8
X_09917_ hold1847/X _16463_/Q _10964_/S vssd1 vssd1 vccd1 vccd1 _09918_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_217_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout643 _12804_/A vssd1 vssd1 vccd1 vccd1 _08361_/A sky130_fd_sc_hd__buf_2
Xfanout654 _12597_/A vssd1 vssd1 vccd1 vccd1 _12612_/A sky130_fd_sc_hd__buf_2
XFILLER_0_226_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout665 _13801_/C1 vssd1 vssd1 vccd1 vccd1 _09272_/A sky130_fd_sc_hd__buf_4
XFILLER_0_176_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout676 fanout689/X vssd1 vssd1 vccd1 vccd1 _12289_/C1 sky130_fd_sc_hd__buf_2
X_09848_ hold2641/X hold3755/X _10985_/S vssd1 vssd1 vccd1 vccd1 _09849_/B sky130_fd_sc_hd__mux2_1
Xfanout687 _14376_/A vssd1 vssd1 vccd1 vccd1 _13901_/A sky130_fd_sc_hd__buf_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout698 _08851_/A vssd1 vssd1 vccd1 vccd1 _12978_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_198_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09779_ hold2257/X _16417_/Q _10067_/C vssd1 vssd1 vccd1 vccd1 _09780_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ hold2999/X hold4745/X _13796_/S vssd1 vssd1 vccd1 vccd1 _11811_/B sky130_fd_sc_hd__mux2_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ hold986/X _17441_/Q _12838_/S vssd1 vssd1 vccd1 vccd1 _12790_/X sky130_fd_sc_hd__mux2_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _17071_/Q _11741_/B _11741_/C vssd1 vssd1 vccd1 vccd1 _11741_/X sky130_fd_sc_hd__and3_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ hold2601/X _14481_/B _14459_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14460_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ hold1534/X _17048_/Q _11789_/C vssd1 vssd1 vccd1 vccd1 _11673_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_37_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10623_ hold3503/X _10554_/A _10622_/X vssd1 vssd1 vccd1 vccd1 _10623_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_181_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13411_ hold4879/X _13829_/B _13410_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13411_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14391_ _14732_/A hold1014/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14392_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16130_ _17325_/CLK _16130_/D vssd1 vssd1 vccd1 vccd1 hold344/A sky130_fd_sc_hd__dfxtp_1
X_13342_ hold3763/X _13795_/A2 _13341_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _13342_/X
+ sky130_fd_sc_hd__o211a_1
X_10554_ _10554_/A _10554_/B vssd1 vssd1 vccd1 vccd1 _10554_/X sky130_fd_sc_hd__or2_1
XFILLER_0_91_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13273_ _13273_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13273_/X sky130_fd_sc_hd__and2_1
X_16061_ _18417_/CLK _16061_/D vssd1 vssd1 vccd1 vccd1 hold806/A sky130_fd_sc_hd__dfxtp_1
X_10485_ _10530_/A _10485_/B vssd1 vssd1 vccd1 vccd1 _10485_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15012_ _15227_/A hold510/A vssd1 vssd1 vccd1 vccd1 _15012_/X sky130_fd_sc_hd__or2_1
X_12224_ hold2993/X _17232_/Q _13409_/S vssd1 vssd1 vccd1 vccd1 _12225_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_121_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12155_ hold2537/X hold5745/X _12362_/C vssd1 vssd1 vccd1 vccd1 _12156_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11106_ _11106_/A _11106_/B vssd1 vssd1 vccd1 vccd1 _11106_/X sky130_fd_sc_hd__or2_1
XFILLER_0_235_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12086_ hold2760/X hold5032/X _13748_/S vssd1 vssd1 vccd1 vccd1 _12087_/B sky130_fd_sc_hd__mux2_1
X_16963_ _17907_/CLK _16963_/D vssd1 vssd1 vccd1 vccd1 _16963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_217_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15914_ _16058_/CLK _15914_/D vssd1 vssd1 vccd1 vccd1 hold785/A sky130_fd_sc_hd__dfxtp_1
X_11037_ _11655_/A _11037_/B vssd1 vssd1 vccd1 vccd1 _11037_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16894_ _18065_/CLK _16894_/D vssd1 vssd1 vccd1 vccd1 _16894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15845_ _17608_/CLK _15845_/D vssd1 vssd1 vccd1 vccd1 _15845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15776_ _17702_/CLK _15776_/D vssd1 vssd1 vccd1 vccd1 _15776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12988_ hold1974/X _17507_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12988_/X sky130_fd_sc_hd__mux2_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17515_ _17516_/CLK hold947/X vssd1 vssd1 vccd1 vccd1 _17515_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14727_ hold2815/X _14718_/B _14726_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14727_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11939_ hold2783/X _17137_/Q _12329_/C vssd1 vssd1 vccd1 vccd1 _11940_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_75_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17446_ _17446_/CLK _17446_/D vssd1 vssd1 vccd1 vccd1 _17446_/Q sky130_fd_sc_hd__dfxtp_1
X_14658_ _15213_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14658_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13609_ hold3952/X _13817_/B _13608_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _13609_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17377_ _17378_/CLK _17377_/D vssd1 vssd1 vccd1 vccd1 _17377_/Q sky130_fd_sc_hd__dfxtp_1
X_14589_ hold1012/X _14612_/B _14588_/X _14895_/C1 vssd1 vssd1 vccd1 vccd1 _14589_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16328_ _18373_/CLK _16328_/D vssd1 vssd1 vccd1 vccd1 _16328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5107 _17282_/Q vssd1 vssd1 vccd1 vccd1 hold5107/X sky130_fd_sc_hd__dlygate4sd3_1
X_16259_ _17360_/CLK _16259_/D vssd1 vssd1 vccd1 vccd1 _16259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5118 _11878_/X vssd1 vssd1 vccd1 vccd1 _17116_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5129 _17167_/Q vssd1 vssd1 vccd1 vccd1 hold5129/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4406 _11781_/Y vssd1 vssd1 vccd1 vccd1 _11782_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4417 _16910_/Q vssd1 vssd1 vccd1 vccd1 hold4417/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4428 _11793_/Y vssd1 vssd1 vccd1 vccd1 _11794_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4439 _12324_/Y vssd1 vssd1 vccd1 vccd1 _12325_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_65_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3705 _11718_/Y vssd1 vssd1 vccd1 vccd1 _11719_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3716 _16357_/Q vssd1 vssd1 vccd1 vccd1 hold3716/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3727 _09556_/X vssd1 vssd1 vccd1 vccd1 _16342_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3738 _17677_/Q vssd1 vssd1 vccd1 vccd1 hold3738/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3749 _12986_/X vssd1 vssd1 vccd1 vccd1 _12987_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07963_ hold1382/X _07978_/B _07962_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _07963_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09702_ _09984_/A _09702_/B vssd1 vssd1 vccd1 vccd1 _09702_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07894_ _14457_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07894_/X sky130_fd_sc_hd__or2_1
XFILLER_0_177_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09633_ _11106_/A _09633_/B vssd1 vssd1 vccd1 vccd1 _09633_/X sky130_fd_sc_hd__or2_1
XFILLER_0_223_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_284_wb_clk_i clkbuf_6_50_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18363_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09564_ _10386_/A _09564_/B vssd1 vssd1 vccd1 vccd1 _09564_/X sky130_fd_sc_hd__or2_1
XFILLER_0_222_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_213_wb_clk_i clkbuf_6_60_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18174_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_214_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08515_ _15519_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08515_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09495_ _14555_/B _14555_/C _09495_/C vssd1 vssd1 vccd1 vccd1 _09498_/B sky130_fd_sc_hd__or3_1
XFILLER_0_81_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08446_ hold1143/X _08433_/B _08445_/X _13675_/C1 vssd1 vssd1 vccd1 vccd1 _08446_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08377_ _08377_/A hold221/X vssd1 vssd1 vccd1 vccd1 hold222/A sky130_fd_sc_hd__and2_1
XFILLER_0_34_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_225_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_225_1367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5630 _17061_/Q vssd1 vssd1 vccd1 vccd1 hold5630/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_10270_ hold5042/X _10070_/B _10269_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _10270_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5641 _17227_/Q vssd1 vssd1 vccd1 vccd1 hold5641/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5652 _11626_/X vssd1 vssd1 vccd1 vccd1 _17032_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5663 _17066_/Q vssd1 vssd1 vccd1 vccd1 hold5663/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5674 _11917_/X vssd1 vssd1 vccd1 vccd1 _17129_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5685 _17085_/Q vssd1 vssd1 vccd1 vccd1 hold5685/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4940 _11671_/X vssd1 vssd1 vccd1 vccd1 _17047_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5696 _11947_/X vssd1 vssd1 vccd1 vccd1 _17139_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4951 _17080_/Q vssd1 vssd1 vccd1 vccd1 hold4951/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4962 _11281_/X vssd1 vssd1 vccd1 vccd1 _16917_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4973 _10867_/X vssd1 vssd1 vccd1 vccd1 _16779_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4984 _12223_/X vssd1 vssd1 vccd1 vccd1 _17231_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4995 _16773_/Q vssd1 vssd1 vccd1 vccd1 hold4995/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout440 fanout485/X vssd1 vssd1 vccd1 vccd1 _13721_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_233_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout451 _11723_/C vssd1 vssd1 vccd1 vccd1 _11732_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_233_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout462 _12332_/C vssd1 vssd1 vccd1 vccd1 _12362_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_205_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout473 _11783_/C vssd1 vssd1 vccd1 vccd1 _12329_/C sky130_fd_sc_hd__clkbuf_8
X_13960_ _15521_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13960_/X sky130_fd_sc_hd__or2_1
Xfanout484 fanout485/X vssd1 vssd1 vccd1 vccd1 _11219_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_219_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout495 _10025_/C vssd1 vssd1 vccd1 vccd1 _10031_/C sky130_fd_sc_hd__buf_6
X_12911_ hold3364/X _12910_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12912_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_213_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13891_ hold361/A hold268/X vssd1 vssd1 vccd1 vccd1 hold295/A sky130_fd_sc_hd__nor2_1
XFILLER_0_201_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15630_ _17194_/CLK _15630_/D vssd1 vssd1 vccd1 vccd1 _15630_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12842_ hold3366/X _12841_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12842_/X sky130_fd_sc_hd__mux2_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _17229_/CLK _15561_/D vssd1 vssd1 vccd1 vccd1 _15561_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12773_ hold3532/X _12772_/X _12839_/S vssd1 vssd1 vccd1 vccd1 _12773_/X sky130_fd_sc_hd__mux2_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _17300_/CLK _17300_/D vssd1 vssd1 vccd1 vccd1 hold800/A sky130_fd_sc_hd__dfxtp_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14512_ hold2316/X _14537_/B _14511_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _14512_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18280_ _18349_/CLK _18280_/D vssd1 vssd1 vccd1 vccd1 _18280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ hold3538/X _11043_/A _11723_/X vssd1 vssd1 vccd1 vccd1 _11724_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _15492_/A hold295/X vssd1 vssd1 vccd1 vccd1 _15505_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_230_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17899_/CLK _17231_/D vssd1 vssd1 vccd1 vccd1 _17231_/Q sky130_fd_sc_hd__dfxtp_1
X_11655_ _11655_/A _11655_/B vssd1 vssd1 vccd1 vccd1 _11655_/X sky130_fd_sc_hd__or2_1
X_14443_ _14443_/A _14443_/B vssd1 vssd1 vccd1 vccd1 _14443_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10606_ _11206_/A _10606_/B vssd1 vssd1 vccd1 vccd1 _16692_/D sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_88_wb_clk_i clkbuf_6_17_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17284_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17162_ _17194_/CLK _17162_/D vssd1 vssd1 vccd1 vccd1 _17162_/Q sky130_fd_sc_hd__dfxtp_1
X_14374_ _14376_/A hold784/X vssd1 vssd1 vccd1 vccd1 _17986_/D sky130_fd_sc_hd__and2_1
X_11586_ _12285_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11586_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16113_ _17336_/CLK _16113_/D vssd1 vssd1 vccd1 vccd1 hold100/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10537_ hold3938/X _10631_/B _10536_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10537_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13325_ hold2335/X hold5720/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13326_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_17_wb_clk_i clkbuf_6_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18437_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17093_ _17093_/CLK _17093_/D vssd1 vssd1 vccd1 vccd1 _17093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16044_ _17300_/CLK _16044_/D vssd1 vssd1 vccd1 vccd1 hold773/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13256_ _13249_/X _13255_/X _13296_/B1 vssd1 vssd1 vccd1 vccd1 _17550_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_204_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10468_ hold3848/X _10568_/B _10467_/X _14895_/C1 vssd1 vssd1 vccd1 vccd1 _10468_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ _13716_/A _12207_/B vssd1 vssd1 vccd1 vccd1 _12207_/X sky130_fd_sc_hd__or2_1
X_13187_ _13186_/X _16916_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13187_/X sky130_fd_sc_hd__mux2_1
X_10399_ hold3337/X _10589_/B _10398_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10399_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12138_ _12243_/A _12138_/B vssd1 vssd1 vccd1 vccd1 _12138_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17995_ _18059_/CLK _17995_/D vssd1 vssd1 vccd1 vccd1 _17995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_236_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12069_ _13482_/A _12069_/B vssd1 vssd1 vccd1 vccd1 _12069_/X sky130_fd_sc_hd__or2_1
X_16946_ _17859_/CLK _16946_/D vssd1 vssd1 vccd1 vccd1 _16946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16877_ _18048_/CLK _16877_/D vssd1 vssd1 vccd1 vccd1 _16877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15828_ _17719_/CLK _15828_/D vssd1 vssd1 vccd1 vccd1 _15828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15759_ _17678_/CLK _15759_/D vssd1 vssd1 vccd1 vccd1 _15759_/Q sky130_fd_sc_hd__dfxtp_1
X_08300_ hold1037/X _08336_/A2 _08299_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _08300_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09280_ _12810_/A hold981/X vssd1 vssd1 vccd1 vccd1 _16251_/D sky130_fd_sc_hd__and2_1
XFILLER_0_74_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08231_ hold1694/X _08268_/B _08230_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08231_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17429_ _17429_/CLK _17429_/D vssd1 vssd1 vccd1 vccd1 _17429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08162_ _15513_/A hold2999/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08163_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08093_ hold1056/X _08088_/B _08092_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _08093_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4203 hold5951/X vssd1 vssd1 vccd1 vccd1 hold5952/A sky130_fd_sc_hd__buf_4
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4214 _15323_/X vssd1 vssd1 vccd1 vccd1 _15324_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4225 _16540_/Q vssd1 vssd1 vccd1 vccd1 hold4225/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4236 _16330_/Q vssd1 vssd1 vccd1 vccd1 _13110_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3502 _10584_/Y vssd1 vssd1 vccd1 vccd1 _10585_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4247 _10648_/Y vssd1 vssd1 vccd1 vccd1 _16706_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4258 _15443_/X vssd1 vssd1 vccd1 vccd1 _15444_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3513 _11211_/Y vssd1 vssd1 vccd1 vccd1 _11212_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3524 _11169_/Y vssd1 vssd1 vccd1 vccd1 _11170_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4269 _12316_/Y vssd1 vssd1 vccd1 vccd1 _17262_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3535 _12791_/X vssd1 vssd1 vccd1 vccd1 _12792_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3546 _09577_/X vssd1 vssd1 vccd1 vccd1 _16349_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2801 _14514_/X vssd1 vssd1 vccd1 vccd1 _18053_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3557 _10300_/X vssd1 vssd1 vccd1 vccd1 _16590_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2812 _08063_/X vssd1 vssd1 vccd1 vccd1 _15671_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08995_ hold320/X hold570/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08996_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3568 _16694_/Q vssd1 vssd1 vccd1 vccd1 _10610_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2823 _08196_/X vssd1 vssd1 vccd1 vccd1 _15734_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_465_wb_clk_i clkbuf_6_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17446_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_103_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2834 _16260_/Q vssd1 vssd1 vccd1 vccd1 hold2834/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3579 _09952_/X vssd1 vssd1 vccd1 vccd1 _16474_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2845 _14155_/X vssd1 vssd1 vccd1 vccd1 _17881_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2856 _18299_/Q vssd1 vssd1 vccd1 vccd1 hold2856/X sky130_fd_sc_hd__dlygate4sd3_1
X_07946_ _14850_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07946_/X sky130_fd_sc_hd__or2_1
Xhold2867 _18171_/Q vssd1 vssd1 vccd1 vccd1 hold2867/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2878 _08057_/X vssd1 vssd1 vccd1 vccd1 _15668_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2889 _14811_/X vssd1 vssd1 vccd1 vccd1 _18195_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_214_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07877_ _15555_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07877_/X sky130_fd_sc_hd__or2_1
XFILLER_0_230_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09616_ hold4604/X _11162_/B _09615_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _09616_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_1352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09547_ hold3560/X _10025_/B _09546_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09547_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09478_ _09483_/C _09478_/B _09478_/C vssd1 vssd1 vccd1 vccd1 _16320_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_47_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08429_ _15163_/A _08433_/B vssd1 vssd1 vccd1 vccd1 _08429_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_191_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11440_ hold5484/X _11726_/B _11439_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _11440_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11371_ hold5261/X _11753_/B _11370_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11371_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10322_ hold2677/X _16598_/Q _10628_/C vssd1 vssd1 vccd1 vccd1 _10323_/B sky130_fd_sc_hd__mux2_1
X_13110_ _13110_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13110_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14090_ _15543_/A _14094_/B vssd1 vssd1 vccd1 vccd1 _14090_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_225_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ hold907/X hold921/X _17523_/Q vssd1 vssd1 vccd1 vccd1 hold922/A sky130_fd_sc_hd__or3b_1
Xhold5460 _17681_/Q vssd1 vssd1 vccd1 vccd1 hold5460/X sky130_fd_sc_hd__dlygate4sd3_1
X_10253_ hold2113/X hold3322/X _10595_/C vssd1 vssd1 vccd1 vccd1 _10254_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_221_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5471 _13381_/X vssd1 vssd1 vccd1 vccd1 _17580_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5482 _17716_/Q vssd1 vssd1 vccd1 vccd1 hold5482/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5493 _13774_/X vssd1 vssd1 vccd1 vccd1 _17711_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4770 _17507_/Q vssd1 vssd1 vccd1 vccd1 hold4770/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10184_ hold2765/X hold3616/X _10571_/C vssd1 vssd1 vccd1 vccd1 _10185_/B sky130_fd_sc_hd__mux2_1
Xhold4781 _17591_/Q vssd1 vssd1 vccd1 vccd1 hold4781/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4792 _12034_/X vssd1 vssd1 vccd1 vccd1 _17168_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16800_ _18067_/CLK _16800_/D vssd1 vssd1 vccd1 vccd1 _16800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17780_ _18428_/CLK _17780_/D vssd1 vssd1 vccd1 vccd1 _17780_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_135_wb_clk_i clkbuf_6_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17341_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14992_ _15207_/A hold510/A vssd1 vssd1 vccd1 vccd1 _14992_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout270 _11556_/A vssd1 vssd1 vccd1 vccd1 _11655_/A sky130_fd_sc_hd__buf_4
Xfanout281 _13599_/A vssd1 vssd1 vccd1 vccd1 _13791_/A sky130_fd_sc_hd__buf_4
X_16731_ _18347_/CLK _16731_/D vssd1 vssd1 vccd1 vccd1 _16731_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout292 _11697_/A vssd1 vssd1 vccd1 vccd1 _12174_/A sky130_fd_sc_hd__buf_4
XFILLER_0_205_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13943_ _13943_/A _13943_/B vssd1 vssd1 vccd1 vccd1 _17779_/D sky130_fd_sc_hd__and2_1
XFILLER_0_199_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16662_ _18188_/CLK _16662_/D vssd1 vssd1 vccd1 vccd1 _16662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13874_ _17745_/Q _13874_/B _13874_/C vssd1 vssd1 vccd1 vccd1 _13874_/X sky130_fd_sc_hd__and3_1
XFILLER_0_198_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18401_ _18401_/CLK _18401_/D vssd1 vssd1 vccd1 vccd1 _18401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15613_ _17209_/CLK _15613_/D vssd1 vssd1 vccd1 vccd1 _15613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12825_ _12837_/A _12825_/B vssd1 vssd1 vccd1 vccd1 _17451_/D sky130_fd_sc_hd__and2_1
X_16593_ _18197_/CLK _16593_/D vssd1 vssd1 vccd1 vccd1 _16593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18332_ _18396_/CLK _18332_/D vssd1 vssd1 vccd1 vccd1 _18332_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15544_ hold2565/X _15547_/B _15543_/Y _12873_/A vssd1 vssd1 vccd1 vccd1 _15544_/X
+ sky130_fd_sc_hd__o211a_1
X_12756_ _12810_/A _12756_/B vssd1 vssd1 vccd1 vccd1 _17428_/D sky130_fd_sc_hd__and2_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18263_ _18393_/CLK _18263_/D vssd1 vssd1 vccd1 vccd1 _18263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ hold5620/X _12335_/B _11706_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _11707_/X
+ sky130_fd_sc_hd__o211a_1
X_15475_ hold851/X _09386_/A _09362_/D hold433/X vssd1 vssd1 vccd1 vccd1 _15475_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12687_ _12849_/A _12687_/B vssd1 vssd1 vccd1 vccd1 _17405_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17214_ _17278_/CLK _17214_/D vssd1 vssd1 vccd1 vccd1 _17214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14426_ hold1933/X _14433_/B _14425_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _14426_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18194_ _18194_/CLK _18194_/D vssd1 vssd1 vccd1 vccd1 _18194_/Q sky130_fd_sc_hd__dfxtp_1
X_11638_ hold5329/X _11732_/B _11637_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _11638_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17145_ _17743_/CLK _17145_/D vssd1 vssd1 vccd1 vccd1 _17145_/Q sky130_fd_sc_hd__dfxtp_1
X_14357_ _15199_/A hold3067/X _14381_/S vssd1 vssd1 vccd1 vccd1 _14358_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11569_ hold5239/X _11765_/B _11568_/X _14346_/A vssd1 vssd1 vccd1 vccd1 _11569_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold707 hold817/X vssd1 vssd1 vccd1 vccd1 hold818/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 hold718/A vssd1 vssd1 vccd1 vccd1 hold718/X sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ hold4278/X _13307_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13308_/X sky130_fd_sc_hd__mux2_2
Xhold729 hold729/A vssd1 vssd1 vccd1 vccd1 hold729/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17076_ _17894_/CLK _17076_/D vssd1 vssd1 vccd1 vccd1 _17076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14288_ hold927/X _14338_/B vssd1 vssd1 vccd1 vccd1 _14288_/X sky130_fd_sc_hd__or2_1
X_16027_ _18425_/CLK _16027_/D vssd1 vssd1 vccd1 vccd1 hold440/A sky130_fd_sc_hd__dfxtp_1
X_13239_ _13311_/A1 _13237_/X _13238_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13239_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2108 _09401_/X vssd1 vssd1 vccd1 vccd1 _09402_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2119 _17911_/Q vssd1 vssd1 vccd1 vccd1 hold2119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07800_ _18461_/Q _18459_/Q vssd1 vssd1 vccd1 vccd1 _07801_/B sky130_fd_sc_hd__nor2_1
X_08780_ _15414_/A _08780_/B vssd1 vssd1 vccd1 vccd1 _16010_/D sky130_fd_sc_hd__and2_1
XFILLER_0_139_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1407 _18036_/Q vssd1 vssd1 vccd1 vccd1 hold1407/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1418 hold6113/X vssd1 vssd1 vccd1 vccd1 hold1418/X sky130_fd_sc_hd__buf_1
X_17978_ _17978_/CLK _17978_/D vssd1 vssd1 vccd1 vccd1 _17978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1429 _15586_/Q vssd1 vssd1 vccd1 vccd1 hold1429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16929_ _17843_/CLK _16929_/D vssd1 vssd1 vccd1 vccd1 _16929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09401_ _15231_/A _16286_/Q _09401_/S vssd1 vssd1 vccd1 vccd1 _09401_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_172_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09332_ hold6067/X _09325_/B _09331_/X _12612_/A vssd1 vssd1 vccd1 vccd1 _09332_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_220_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09263_ _15539_/A hold1668/X hold271/X vssd1 vssd1 vccd1 vccd1 _09264_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08214_ hold2398/X _08213_/B _08213_/Y _08385_/A vssd1 vssd1 vccd1 vccd1 _08214_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09194_ hold933/X _09230_/B vssd1 vssd1 vccd1 vccd1 _09194_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08145_ _08145_/A _08145_/B vssd1 vssd1 vccd1 vccd1 _15711_/D sky130_fd_sc_hd__and2_1
XFILLER_0_161_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08076_ _14529_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08076_/X sky130_fd_sc_hd__or2_1
XFILLER_0_222_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4000 _10144_/X vssd1 vssd1 vccd1 vccd1 _16538_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4011 _17143_/Q vssd1 vssd1 vccd1 vccd1 hold4011/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4022 _17124_/Q vssd1 vssd1 vccd1 vccd1 hold4022/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_222_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4033 _11959_/X vssd1 vssd1 vccd1 vccd1 _17143_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4044 _17271_/Q vssd1 vssd1 vccd1 vccd1 _12341_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3310 _16844_/Q vssd1 vssd1 vccd1 vccd1 hold3310/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4055 _10330_/X vssd1 vssd1 vccd1 vccd1 _16600_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3321 _10207_/X vssd1 vssd1 vccd1 vccd1 _16559_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4066 _17626_/Q vssd1 vssd1 vccd1 vccd1 hold4066/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4077 _17608_/Q vssd1 vssd1 vccd1 vccd1 hold4077/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3332 _17479_/Q vssd1 vssd1 vccd1 vccd1 hold3332/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3343 _17392_/Q vssd1 vssd1 vccd1 vccd1 hold3343/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4088 _11551_/X vssd1 vssd1 vccd1 vccd1 _17007_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3354 _17476_/Q vssd1 vssd1 vccd1 vccd1 hold3354/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4099 _16868_/Q vssd1 vssd1 vccd1 vccd1 hold4099/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2620 _18229_/Q vssd1 vssd1 vccd1 vccd1 hold2620/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3365 _17371_/Q vssd1 vssd1 vccd1 vccd1 hold3365/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__clkbuf_4
XTAP_5538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2631 _18339_/Q vssd1 vssd1 vccd1 vccd1 hold2631/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3376 _17404_/Q vssd1 vssd1 vccd1 vccd1 hold3376/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3387 hold5962/X vssd1 vssd1 vccd1 vccd1 hold5963/A sky130_fd_sc_hd__buf_6
Xhold2642 _15140_/X vssd1 vssd1 vccd1 vccd1 _18353_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _12394_/A _08978_/B vssd1 vssd1 vccd1 vccd1 _16106_/D sky130_fd_sc_hd__and2_1
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2653 _14621_/X vssd1 vssd1 vccd1 vccd1 _18104_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3398 _17459_/Q vssd1 vssd1 vccd1 vccd1 hold3398/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__buf_4
Xhold2664 _18190_/Q vssd1 vssd1 vccd1 vccd1 hold2664/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2675 _18396_/Q vssd1 vssd1 vccd1 vccd1 hold2675/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1930 _09223_/X vssd1 vssd1 vccd1 vccd1 _16223_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1941 _18322_/Q vssd1 vssd1 vccd1 vccd1 hold1941/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2686 _14693_/X vssd1 vssd1 vccd1 vccd1 _18138_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ hold1602/X _07924_/B _07928_/X _12822_/A vssd1 vssd1 vccd1 vccd1 _07929_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_231_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2697 _15590_/Q vssd1 vssd1 vccd1 vccd1 hold2697/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1952 _14546_/X vssd1 vssd1 vccd1 vccd1 _18069_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1963 _14169_/X vssd1 vssd1 vccd1 vccd1 _17887_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1974 _16170_/Q vssd1 vssd1 vccd1 vccd1 hold1974/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1985 _14605_/X vssd1 vssd1 vccd1 vccd1 _18096_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10940_ hold1897/X hold5364/X _11738_/C vssd1 vssd1 vccd1 vccd1 _10941_/B sky130_fd_sc_hd__mux2_1
Xhold1996 _16267_/Q vssd1 vssd1 vccd1 vccd1 hold1996/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10871_ hold1587/X hold4837/X _11162_/C vssd1 vssd1 vccd1 vccd1 _10872_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_210_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ hold1297/X _17381_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12610_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _13791_/A _13590_/B vssd1 vssd1 vccd1 vccd1 _13590_/X sky130_fd_sc_hd__or2_1
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12541_ hold1473/X _17358_/Q _12925_/S vssd1 vssd1 vccd1 vccd1 _12541_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_108_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15260_ _15911_/Q _15448_/A2 _15446_/B1 hold187/X vssd1 vssd1 vccd1 vccd1 _15260_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12472_ _17329_/Q _12506_/B vssd1 vssd1 vccd1 vccd1 _12472_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14211_ hold1416/X _14198_/B _14210_/X _14211_/C1 vssd1 vssd1 vccd1 vccd1 _14211_/X
+ sky130_fd_sc_hd__o211a_1
X_11423_ hold2873/X hold5591/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11424_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_105_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15191_ _15191_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15191_/X sky130_fd_sc_hd__or2_1
XFILLER_0_152_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_9 _13116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14142_ _15215_/A _14142_/B vssd1 vssd1 vccd1 vccd1 _14142_/Y sky130_fd_sc_hd__nand2_1
X_11354_ hold1787/X hold5390/X _11654_/S vssd1 vssd1 vccd1 vccd1 _11355_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_387_wb_clk_i clkbuf_6_35_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17236_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_127_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10305_ _10563_/A _10305_/B vssd1 vssd1 vccd1 vccd1 _10305_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14073_ hold2244/X _14107_/A2 _14072_/X _14143_/C1 vssd1 vssd1 vccd1 vccd1 _14073_/X
+ sky130_fd_sc_hd__o211a_1
X_11285_ _17767_/Q hold4337/X _11765_/C vssd1 vssd1 vccd1 vccd1 _11286_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_316_wb_clk_i clkbuf_6_47_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18036_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_120_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5290 _13648_/X vssd1 vssd1 vccd1 vccd1 _17669_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13024_ hold937/X hold904/A vssd1 vssd1 vccd1 vccd1 _13025_/C sky130_fd_sc_hd__nand2_1
X_10236_ _10542_/A _10236_/B vssd1 vssd1 vccd1 vccd1 _10236_/X sky130_fd_sc_hd__or2_1
XFILLER_0_197_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17901_ _17901_/CLK _17901_/D vssd1 vssd1 vccd1 vccd1 _17901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17832_ _17832_/CLK _17832_/D vssd1 vssd1 vccd1 vccd1 _17832_/Q sky130_fd_sc_hd__dfxtp_1
X_10167_ _10515_/A _10167_/B vssd1 vssd1 vccd1 vccd1 _10167_/X sky130_fd_sc_hd__or2_1
XFILLER_0_233_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17763_ _17892_/CLK _17763_/D vssd1 vssd1 vccd1 vccd1 _17763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_238_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10098_ _10482_/A _10098_/B vssd1 vssd1 vccd1 vccd1 _10098_/X sky130_fd_sc_hd__or2_1
X_14975_ hold6075/X hold447/X _14974_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _14975_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16714_ _18045_/CLK _16714_/D vssd1 vssd1 vccd1 vccd1 _16714_/Q sky130_fd_sc_hd__dfxtp_1
X_13926_ hold384/X _17771_/Q hold297/X vssd1 vssd1 vccd1 vccd1 hold385/A sky130_fd_sc_hd__mux2_1
X_17694_ _17726_/CLK _17694_/D vssd1 vssd1 vccd1 vccd1 _17694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_236_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16645_ _18203_/CLK _16645_/D vssd1 vssd1 vccd1 vccd1 _16645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13857_ hold4408/X _13752_/A _13856_/X vssd1 vssd1 vccd1 vccd1 _13857_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_202_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12808_ hold1572/X _17447_/Q _12811_/S vssd1 vssd1 vccd1 vccd1 _12808_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16576_ _18166_/CLK _16576_/D vssd1 vssd1 vccd1 vccd1 _16576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13788_ _13788_/A _13788_/B vssd1 vssd1 vccd1 vccd1 _13788_/X sky130_fd_sc_hd__or2_1
XFILLER_0_128_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18315_ _18315_/CLK hold237/X vssd1 vssd1 vccd1 vccd1 _18315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15527_ hold951/X _15559_/B vssd1 vssd1 vccd1 vccd1 _15527_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_wb_clk_i clkbuf_6_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18045_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12739_ hold572/X hold3173/X _12811_/S vssd1 vssd1 vccd1 vccd1 _12739_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_155_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18246_ _18334_/CLK _18246_/D vssd1 vssd1 vccd1 vccd1 _18246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15458_ hold859/X _09367_/A _09362_/C hold794/X vssd1 vssd1 vccd1 vccd1 _15458_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14409_ _14517_/A _14443_/B vssd1 vssd1 vccd1 vccd1 _14409_/X sky130_fd_sc_hd__or2_1
X_18177_ _18177_/CLK _18177_/D vssd1 vssd1 vccd1 vccd1 _18177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ hold869/X _09365_/B _09392_/C hold656/X _15388_/X vssd1 vssd1 vccd1 vccd1
+ _15392_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_170_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold504 hold504/A vssd1 vssd1 vccd1 vccd1 hold504/X sky130_fd_sc_hd__dlygate4sd3_1
X_17128_ _17628_/CLK _17128_/D vssd1 vssd1 vccd1 vccd1 _17128_/Q sky130_fd_sc_hd__dfxtp_1
Xhold515 hold515/A vssd1 vssd1 vccd1 vccd1 hold515/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold526 hold526/A vssd1 vssd1 vccd1 vccd1 hold526/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 hold537/A vssd1 vssd1 vccd1 vccd1 hold537/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold548 hold576/X vssd1 vssd1 vccd1 vccd1 hold577/A sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ hold1869/X hold3543/X _10067_/C vssd1 vssd1 vccd1 vccd1 _09951_/B sky130_fd_sc_hd__mux2_1
Xhold559 hold559/A vssd1 vssd1 vccd1 vccd1 hold559/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17059_ _17907_/CLK _17059_/D vssd1 vssd1 vccd1 vccd1 _17059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08901_ _09440_/B hold729/X vssd1 vssd1 vccd1 vccd1 _16068_/D sky130_fd_sc_hd__and2_1
X_09881_ hold1503/X _16451_/Q _10049_/C vssd1 vssd1 vccd1 vccd1 _09882_/B sky130_fd_sc_hd__mux2_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ hold172/X hold890/X _08866_/S vssd1 vssd1 vccd1 vccd1 _08833_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_237_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1204 _08308_/X vssd1 vssd1 vccd1 vccd1 _15787_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1215 _15800_/Q vssd1 vssd1 vccd1 vccd1 hold1215/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 _15823_/Q vssd1 vssd1 vccd1 vccd1 hold1226/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1237 _16242_/Q vssd1 vssd1 vccd1 vccd1 hold1237/X sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ hold185/X hold563/X _08779_/S vssd1 vssd1 vccd1 vccd1 hold564/A sky130_fd_sc_hd__mux2_1
Xhold1248 _16213_/Q vssd1 vssd1 vccd1 vccd1 hold1248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1259 _14079_/X vssd1 vssd1 vccd1 vccd1 _17844_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ _12410_/A _08694_/B vssd1 vssd1 vccd1 vccd1 _15968_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09315_ _15103_/A _09315_/B vssd1 vssd1 vccd1 vccd1 _09315_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09246_ _12786_/A _09246_/B vssd1 vssd1 vccd1 vccd1 _16234_/D sky130_fd_sc_hd__and2_1
XFILLER_0_173_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09177_ hold1319/X _09177_/A2 _09176_/X _12924_/A vssd1 vssd1 vccd1 vccd1 _09177_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08128_ _15533_/A hold2622/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08129_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08059_ hold2705/X _08097_/A2 _08058_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _08059_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11070_ _11556_/A _11070_/B vssd1 vssd1 vccd1 vccd1 _11070_/X sky130_fd_sc_hd__or2_1
XTAP_6025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput79 _13185_/A vssd1 vssd1 vccd1 vccd1 output79/X sky130_fd_sc_hd__buf_6
XTAP_6036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3140 _12632_/X vssd1 vssd1 vccd1 vccd1 _12633_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10021_ _10603_/A _10021_/B vssd1 vssd1 vccd1 vccd1 _10021_/Y sky130_fd_sc_hd__nor2_1
XTAP_5313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3151 _17398_/Q vssd1 vssd1 vccd1 vccd1 hold3151/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3162 _12737_/X vssd1 vssd1 vccd1 vccd1 _12738_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3173 _17424_/Q vssd1 vssd1 vccd1 vccd1 hold3173/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3184 _18351_/Q vssd1 vssd1 vccd1 vccd1 hold3184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3195 _16351_/Q vssd1 vssd1 vccd1 vccd1 _13278_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2450 _08004_/X vssd1 vssd1 vccd1 vccd1 _15643_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2461 _14149_/X vssd1 vssd1 vccd1 vccd1 _17878_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2472 _18451_/Q vssd1 vssd1 vccd1 vccd1 hold2472/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2483 _18215_/Q vssd1 vssd1 vccd1 vccd1 hold2483/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2494 _14747_/X vssd1 vssd1 vccd1 vccd1 _18164_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1760 _15868_/Q vssd1 vssd1 vccd1 vccd1 hold1760/X sky130_fd_sc_hd__dlygate4sd3_1
X_14760_ _15099_/A _14780_/B vssd1 vssd1 vccd1 vccd1 _14760_/X sky130_fd_sc_hd__or2_1
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1771 _08286_/X vssd1 vssd1 vccd1 vccd1 _15776_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1782 _14777_/X vssd1 vssd1 vccd1 vccd1 _18179_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11972_ hold1279/X _17148_/Q _13481_/S vssd1 vssd1 vccd1 vccd1 _11973_/B sky130_fd_sc_hd__mux2_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1793 _15765_/Q vssd1 vssd1 vccd1 vccd1 hold1793/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13711_ hold5783/X _13808_/B _13710_/X _12738_/A vssd1 vssd1 vccd1 vccd1 _13711_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10923_ _11100_/A _10923_/B vssd1 vssd1 vccd1 vccd1 _10923_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_230_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14691_ hold2518/X _14718_/B _14690_/X _14691_/C1 vssd1 vssd1 vccd1 vccd1 _14691_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16430_ _18375_/CLK _16430_/D vssd1 vssd1 vccd1 vccd1 _16430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13642_ hold4764/X _13862_/B _13641_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _13642_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10854_ _11049_/A _10854_/B vssd1 vssd1 vccd1 vccd1 _10854_/X sky130_fd_sc_hd__or2_1
XFILLER_0_211_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16361_ _18368_/CLK _16361_/D vssd1 vssd1 vccd1 vccd1 _16361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13573_ hold5521/X _13847_/B _13572_/X _13765_/C1 vssd1 vssd1 vccd1 vccd1 _13573_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ _11655_/A _10785_/B vssd1 vssd1 vccd1 vccd1 _10785_/X sky130_fd_sc_hd__or2_1
XFILLER_0_13_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18100_ _18210_/CLK _18100_/D vssd1 vssd1 vccd1 vccd1 _18100_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15312_ _15480_/A _15312_/B _15312_/C _15312_/D vssd1 vssd1 vccd1 vccd1 _15312_/X
+ sky130_fd_sc_hd__or4_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12524_ hold4474/X _12523_/X _12929_/S vssd1 vssd1 vccd1 vccd1 _12525_/B sky130_fd_sc_hd__mux2_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _18404_/CLK _16292_/D vssd1 vssd1 vccd1 vccd1 _16292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18031_ _18031_/CLK _18031_/D vssd1 vssd1 vccd1 vccd1 _18031_/Q sky130_fd_sc_hd__dfxtp_1
X_15243_ _15490_/A1 _15235_/X _15242_/X _15490_/B1 hold4201/X vssd1 vssd1 vccd1 vccd1
+ _15243_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_87_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12455_ hold71/X _12445_/A _12445_/B _12454_/X _12394_/A vssd1 vssd1 vccd1 vccd1
+ hold72/A sky130_fd_sc_hd__o311a_1
XFILLER_0_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11406_ _12174_/A _11406_/B vssd1 vssd1 vccd1 vccd1 _11406_/X sky130_fd_sc_hd__or2_1
X_15174_ hold6065/X _15165_/B hold1139/X _15042_/A vssd1 vssd1 vccd1 vccd1 _15174_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12386_ _15414_/A hold391/X vssd1 vssd1 vccd1 vccd1 _17286_/D sky130_fd_sc_hd__and2_1
X_14125_ hold1070/X _14142_/B _14124_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _14125_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_239_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11337_ _12210_/A _11337_/B vssd1 vssd1 vccd1 vccd1 _11337_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_150_wb_clk_i clkbuf_6_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18368_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14056_ _14395_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14056_/X sky130_fd_sc_hd__or2_1
X_11268_ _12219_/A _11268_/B vssd1 vssd1 vccd1 vccd1 _11268_/X sky130_fd_sc_hd__or2_1
XFILLER_0_197_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ _14970_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13007_/X sky130_fd_sc_hd__or2_1
X_10219_ hold3899/X _10619_/B _10218_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10219_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11199_ hold3517/X _11127_/A _11198_/X vssd1 vssd1 vccd1 vccd1 _11199_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17815_ _17847_/CLK _17815_/D vssd1 vssd1 vccd1 vccd1 _17815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_234_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17746_ _17746_/CLK _17746_/D vssd1 vssd1 vccd1 vccd1 _17746_/Q sky130_fd_sc_hd__dfxtp_1
X_14958_ _15227_/A hold407/X vssd1 vssd1 vccd1 vccd1 _14958_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13909_ _13909_/A hold972/X vssd1 vssd1 vccd1 vccd1 _17762_/D sky130_fd_sc_hd__and2_1
X_17677_ _17709_/CLK _17677_/D vssd1 vssd1 vccd1 vccd1 _17677_/Q sky130_fd_sc_hd__dfxtp_1
X_14889_ hold2854/X _14880_/B _14888_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14889_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_6_43_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_43_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_212_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16628_ _18166_/CLK _16628_/D vssd1 vssd1 vccd1 vccd1 _16628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16559_ _18213_/CLK _16559_/D vssd1 vssd1 vccd1 vccd1 _16559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09100_ _15541_/A _09102_/B vssd1 vssd1 vccd1 vccd1 _09100_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09031_ _12438_/A hold181/X vssd1 vssd1 vccd1 vccd1 _16132_/D sky130_fd_sc_hd__and2_1
X_18229_ _18229_/CLK _18229_/D vssd1 vssd1 vccd1 vccd1 _18229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_238_wb_clk_i clkbuf_6_60_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18225_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_142_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold301 hold301/A vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold312 hold312/A vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 hold323/A vssd1 vssd1 vccd1 vccd1 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold334 la_data_in[28] vssd1 vssd1 vccd1 vccd1 hold334/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold345 hold345/A vssd1 vssd1 vccd1 vccd1 hold345/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 hold356/A vssd1 vssd1 vccd1 vccd1 hold356/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold367 hold931/X vssd1 vssd1 vccd1 vccd1 hold932/A sky130_fd_sc_hd__buf_6
Xhold378 hold378/A vssd1 vssd1 vccd1 vccd1 hold378/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 hold389/A vssd1 vssd1 vccd1 vccd1 hold389/X sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ _09933_/A _09933_/B vssd1 vssd1 vccd1 vccd1 _09933_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout803 fanout816/X vssd1 vssd1 vccd1 vccd1 _15019_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout814 _15204_/C1 vssd1 vssd1 vccd1 vccd1 _15030_/A sky130_fd_sc_hd__buf_4
XFILLER_0_1_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout825 _14390_/A vssd1 vssd1 vccd1 vccd1 _14542_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout836 fanout843/X vssd1 vssd1 vccd1 vccd1 _14869_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09864_ _09954_/A _09864_/B vssd1 vssd1 vccd1 vccd1 _09864_/X sky130_fd_sc_hd__or2_1
Xfanout847 _17754_/Q vssd1 vssd1 vccd1 vccd1 _13873_/A sky130_fd_sc_hd__buf_8
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout858 _13312_/B1 vssd1 vssd1 vccd1 vccd1 _13296_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_176_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 _14953_/X vssd1 vssd1 vccd1 vccd1 _18263_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout869 _15219_/A vssd1 vssd1 vccd1 vccd1 _15545_/A sky130_fd_sc_hd__buf_12
Xhold1012 _18088_/Q vssd1 vssd1 vccd1 vccd1 hold1012/X sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ _15364_/A _08815_/B vssd1 vssd1 vccd1 vccd1 _16026_/D sky130_fd_sc_hd__and2_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 _14166_/A vssd1 vssd1 vccd1 vccd1 _15511_/A sky130_fd_sc_hd__buf_4
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1034 _14775_/X vssd1 vssd1 vccd1 vccd1 _18178_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ _09987_/A _09795_/B vssd1 vssd1 vccd1 vccd1 _09795_/X sky130_fd_sc_hd__or2_1
Xhold1045 _15839_/Q vssd1 vssd1 vccd1 vccd1 hold1045/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1056 _15686_/Q vssd1 vssd1 vccd1 vccd1 hold1056/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1067 _18021_/Q vssd1 vssd1 vccd1 vccd1 hold1067/X sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ _15284_/A hold871/X vssd1 vssd1 vccd1 vccd1 _15993_/D sky130_fd_sc_hd__and2_1
XFILLER_0_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1078 _13919_/X vssd1 vssd1 vccd1 vccd1 _17767_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 _18218_/Q vssd1 vssd1 vccd1 vccd1 hold1089/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ hold29/X hold323/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08678_/B sky130_fd_sc_hd__mux2_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_240_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10570_ _10603_/A _10570_/B vssd1 vssd1 vccd1 vccd1 _16680_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09229_ hold1708/X _09218_/B _09228_/X _12843_/A vssd1 vssd1 vccd1 vccd1 _09229_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12240_ _12240_/A _12240_/B vssd1 vssd1 vccd1 vccd1 _12240_/X sky130_fd_sc_hd__or2_1
XFILLER_0_224_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12171_ _12267_/A _12171_/B vssd1 vssd1 vccd1 vccd1 _12171_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11122_ hold5095/X _11225_/B _11121_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _11122_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold890 hold890/A vssd1 vssd1 vccd1 vccd1 hold890/X sky130_fd_sc_hd__dlygate4sd3_1
X_15930_ _17520_/CLK _15930_/D vssd1 vssd1 vccd1 vccd1 _15930_/Q sky130_fd_sc_hd__dfxtp_1
X_11053_ hold5026/X _11153_/B _11052_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _11053_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10004_ _16492_/Q _10004_/B _10004_/C vssd1 vssd1 vccd1 vccd1 _10004_/X sky130_fd_sc_hd__and3_1
XTAP_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15861_ _17648_/CLK _15861_/D vssd1 vssd1 vccd1 vccd1 _15861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2280 _14564_/X vssd1 vssd1 vccd1 vccd1 hold2280/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _17728_/CLK _17600_/D vssd1 vssd1 vccd1 vccd1 _17600_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812_ _15205_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14812_/X sky130_fd_sc_hd__or2_1
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2291 _17759_/Q vssd1 vssd1 vccd1 vccd1 hold2291/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15792_ _17689_/CLK _15792_/D vssd1 vssd1 vccd1 vccd1 _15792_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ _17535_/CLK _17531_/D vssd1 vssd1 vccd1 vccd1 _17531_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1590 _15614_/Q vssd1 vssd1 vccd1 vccd1 hold1590/X sky130_fd_sc_hd__dlygate4sd3_1
X_14743_ hold3045/X _14774_/B _14742_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14743_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ _12174_/A _11955_/B vssd1 vssd1 vccd1 vccd1 _11955_/X sky130_fd_sc_hd__or2_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10906_ hold4959/X _11222_/B _10905_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _10906_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17462_ _17462_/CLK _17462_/D vssd1 vssd1 vccd1 vccd1 _17462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14674_ _15229_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14674_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11886_ _12174_/A _11886_/B vssd1 vssd1 vccd1 vccd1 _11886_/X sky130_fd_sc_hd__or2_1
X_16413_ _18384_/CLK _16413_/D vssd1 vssd1 vccd1 vccd1 _16413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13625_ hold2326/X hold4689/X _13817_/C vssd1 vssd1 vccd1 vccd1 _13626_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_7_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17393_ _18453_/CLK _17393_/D vssd1 vssd1 vccd1 vccd1 _17393_/Q sky130_fd_sc_hd__dfxtp_1
X_10837_ hold3820/X _11222_/B _10836_/X _14346_/A vssd1 vssd1 vccd1 vccd1 _10837_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16344_ _18327_/CLK _16344_/D vssd1 vssd1 vccd1 vccd1 _16344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13556_ hold2661/X _17639_/Q _13880_/C vssd1 vssd1 vccd1 vccd1 _13557_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10768_ hold4127/X _11723_/B _10767_/X _14364_/A vssd1 vssd1 vccd1 vccd1 _10768_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12507_ hold44/X _12509_/A2 _08868_/X _12506_/X _09061_/A vssd1 vssd1 vccd1 vccd1
+ hold45/A sky130_fd_sc_hd__o311a_1
XFILLER_0_54_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16275_ _17374_/CLK _16275_/D vssd1 vssd1 vccd1 vccd1 _16275_/Q sky130_fd_sc_hd__dfxtp_1
X_13487_ hold1143/X _17616_/Q _13865_/C vssd1 vssd1 vccd1 vccd1 _13488_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_331_wb_clk_i clkbuf_6_41_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17272_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_207_1416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10699_ hold4853/X _11171_/B _10698_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _10699_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18014_ _18014_/CLK _18014_/D vssd1 vssd1 vccd1 vccd1 _18014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15226_ hold1805/X _15221_/B _15225_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _15226_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12438_ _12438_/A hold95/X vssd1 vssd1 vccd1 vccd1 _17312_/D sky130_fd_sc_hd__and2_1
XFILLER_0_140_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15157_ hold630/X _15157_/B vssd1 vssd1 vccd1 vccd1 hold631/A sky130_fd_sc_hd__or2_1
XFILLER_0_140_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12369_ hold4332/X _13407_/A _12368_/X vssd1 vssd1 vccd1 vccd1 _12369_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3909 _17654_/Q vssd1 vssd1 vccd1 vccd1 hold3909/X sky130_fd_sc_hd__dlygate4sd3_1
X_14108_ _14789_/A _14163_/B vssd1 vssd1 vccd1 vccd1 _14108_/Y sky130_fd_sc_hd__nor2_2
X_15088_ hold6073/X hold341/X hold1466/X _15212_/C1 vssd1 vssd1 vccd1 vccd1 _15088_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14039_ hold2418/X _14038_/B _14038_/Y _13903_/A vssd1 vssd1 vccd1 vccd1 _14039_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08600_ _12416_/A hold723/X vssd1 vssd1 vccd1 vccd1 _15922_/D sky130_fd_sc_hd__and2_1
X_09580_ hold3606/X _10052_/B _09579_/X _15019_/C1 vssd1 vssd1 vccd1 vccd1 _09580_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08531_ _13046_/C _12380_/A vssd1 vssd1 vccd1 vccd1 _08544_/S sky130_fd_sc_hd__or2_2
XFILLER_0_179_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17729_ _17729_/CLK _17729_/D vssd1 vssd1 vccd1 vccd1 _17729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08462_ _14461_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08462_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08393_ _08504_/A hold445/X vssd1 vssd1 vccd1 vccd1 _08393_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_86_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_419_wb_clk_i clkbuf_6_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17093_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09014_ hold679/X hold755/X _09060_/S vssd1 vssd1 vccd1 vccd1 hold756/A sky130_fd_sc_hd__mux2_1
Xhold5801 _17595_/Q vssd1 vssd1 vccd1 vccd1 hold5801/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5812 _09982_/X vssd1 vssd1 vccd1 vccd1 _16484_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5823 _16462_/Q vssd1 vssd1 vccd1 vccd1 hold5823/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5834 _09940_/X vssd1 vssd1 vccd1 vccd1 _16470_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5845 hold6006/X vssd1 vssd1 vccd1 vccd1 _13233_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 hold120/A vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5856 output77/X vssd1 vssd1 vccd1 vccd1 data_out[14] sky130_fd_sc_hd__buf_12
Xhold131 hold38/X vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_143_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5867 hold6015/X vssd1 vssd1 vccd1 vccd1 _13129_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 input21/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__buf_1
XFILLER_0_112_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold153 hold153/A vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5878 output84/X vssd1 vssd1 vccd1 vccd1 data_out[20] sky130_fd_sc_hd__buf_12
Xhold5889 hold6029/X vssd1 vssd1 vccd1 vccd1 _13305_/A sky130_fd_sc_hd__buf_1
XFILLER_0_223_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold164 hold164/A vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 hold175/A vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold186 hold186/A vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 hold197/A vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 _12970_/S vssd1 vssd1 vccd1 vccd1 _12985_/S sky130_fd_sc_hd__clkbuf_8
Xfanout611 _09361_/Y vssd1 vssd1 vccd1 vccd1 _15485_/B1 sky130_fd_sc_hd__buf_8
XFILLER_0_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09916_ hold5827/X _10022_/B _09915_/X _15202_/C1 vssd1 vssd1 vccd1 vccd1 _09916_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout622 _15485_/A2 vssd1 vssd1 vccd1 vccd1 _09365_/B sky130_fd_sc_hd__buf_8
Xfanout633 _08597_/Y vssd1 vssd1 vccd1 vccd1 _12445_/A sky130_fd_sc_hd__buf_6
XFILLER_0_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout644 _12199_/C1 vssd1 vssd1 vccd1 vccd1 _12804_/A sky130_fd_sc_hd__buf_2
Xfanout655 _12597_/A vssd1 vssd1 vccd1 vccd1 _12906_/A sky130_fd_sc_hd__buf_4
Xfanout666 fanout689/X vssd1 vssd1 vccd1 vccd1 _13801_/C1 sky130_fd_sc_hd__buf_2
X_09847_ hold3680/X _10577_/B _09846_/X _15146_/C1 vssd1 vssd1 vccd1 vccd1 _09847_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout677 _15498_/A vssd1 vssd1 vccd1 vccd1 _14147_/C1 sky130_fd_sc_hd__buf_4
Xfanout688 fanout689/X vssd1 vssd1 vccd1 vccd1 _14376_/A sky130_fd_sc_hd__clkbuf_4
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout699 _09440_/B vssd1 vssd1 vccd1 vccd1 _15274_/A sky130_fd_sc_hd__buf_4
XFILLER_0_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09778_ hold3744/X _10046_/B _09777_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09778_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _17519_/Q hold948/X vssd1 vssd1 vccd1 vccd1 _08934_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_198_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _12301_/A _11740_/B vssd1 vssd1 vccd1 vccd1 _17070_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_205_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ hold4939/X _11765_/B _11670_/X _14346_/A vssd1 vssd1 vccd1 vccd1 _11671_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13410_ _13734_/A _13410_/B vssd1 vssd1 vccd1 vccd1 _13410_/X sky130_fd_sc_hd__or2_1
X_10622_ _16698_/Q _10649_/B _10640_/C vssd1 vssd1 vccd1 vccd1 _10622_/X sky130_fd_sc_hd__and3_1
XFILLER_0_187_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14390_ _14390_/A _14390_/B vssd1 vssd1 vccd1 vccd1 _17994_/D sky130_fd_sc_hd__and2_1
XFILLER_0_63_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13341_ _13794_/A _13341_/B vssd1 vssd1 vccd1 vccd1 _13341_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10553_ hold2854/X _16675_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10554_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_165_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16060_ _17291_/CLK _16060_/D vssd1 vssd1 vccd1 vccd1 hold880/A sky130_fd_sc_hd__dfxtp_1
X_13272_ _13265_/X _13271_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17552_/D sky130_fd_sc_hd__o21a_1
X_10484_ hold1313/X _16652_/Q _10625_/C vssd1 vssd1 vccd1 vccd1 _10485_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15011_ hold2081/X hold447/X _15010_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _15011_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12223_ hold4983/X _12317_/B _12222_/X _14211_/C1 vssd1 vssd1 vccd1 vccd1 _12223_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12154_ hold4913/X _12374_/B _12153_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _12154_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_1346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11105_ hold1885/X _16859_/Q _11201_/C vssd1 vssd1 vccd1 vccd1 _11106_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_236_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12085_ hold5078/X _12365_/B _12084_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _12085_/X
+ sky130_fd_sc_hd__o211a_1
X_16962_ _17873_/CLK _16962_/D vssd1 vssd1 vccd1 vccd1 _16962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15913_ _16093_/CLK _15913_/D vssd1 vssd1 vccd1 vccd1 hold620/A sky130_fd_sc_hd__dfxtp_1
X_11036_ hold1348/X _16836_/Q _11168_/C vssd1 vssd1 vccd1 vccd1 _11037_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_235_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16893_ _17968_/CLK _16893_/D vssd1 vssd1 vccd1 vccd1 _16893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_217_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15844_ _17703_/CLK _15844_/D vssd1 vssd1 vccd1 vccd1 _15844_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15775_ _17726_/CLK _15775_/D vssd1 vssd1 vccd1 vccd1 _15775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12987_ _12987_/A _12987_/B vssd1 vssd1 vccd1 vccd1 _17505_/D sky130_fd_sc_hd__and2_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _14726_/A _14730_/B vssd1 vssd1 vccd1 vccd1 _14726_/X sky130_fd_sc_hd__or2_1
X_17514_ _17514_/CLK _17514_/D vssd1 vssd1 vccd1 vccd1 _17514_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11938_ hold3818/X _12353_/B _11937_/X _12289_/C1 vssd1 vssd1 vccd1 vccd1 _11938_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17445_ _17445_/CLK _17445_/D vssd1 vssd1 vccd1 vccd1 _17445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14657_ hold1889/X _14664_/B _14656_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14657_/X
+ sky130_fd_sc_hd__o211a_1
X_11869_ hold5741/X _12350_/B _11868_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _11869_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13608_ _13722_/A _13608_/B vssd1 vssd1 vccd1 vccd1 _13608_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17376_ _17378_/CLK _17376_/D vssd1 vssd1 vccd1 vccd1 _17376_/Q sky130_fd_sc_hd__dfxtp_1
X_14588_ _15197_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14588_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16327_ _18424_/CLK _16327_/D vssd1 vssd1 vccd1 vccd1 _16327_/Q sky130_fd_sc_hd__dfxtp_1
X_13539_ _13734_/A _13539_/B vssd1 vssd1 vccd1 vccd1 _13539_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16258_ _17360_/CLK _16258_/D vssd1 vssd1 vccd1 vccd1 _16258_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5108 _12280_/X vssd1 vssd1 vccd1 vccd1 _17250_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5119 _16850_/Q vssd1 vssd1 vccd1 vccd1 hold5119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15209_ _15209_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15209_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4407 _11782_/Y vssd1 vssd1 vccd1 vccd1 _17084_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16189_ _17882_/CLK _16189_/D vssd1 vssd1 vccd1 vccd1 _16189_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4418 _11739_/Y vssd1 vssd1 vccd1 vccd1 _11740_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4429 _11794_/Y vssd1 vssd1 vccd1 vccd1 _17088_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3706 _16551_/Q vssd1 vssd1 vccd1 vccd1 hold3706/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3717 _09505_/X vssd1 vssd1 vccd1 vccd1 _16325_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3728 _17686_/Q vssd1 vssd1 vccd1 vccd1 hold3728/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3739 _13576_/X vssd1 vssd1 vccd1 vccd1 _17645_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07962_ _15531_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07962_/X sky130_fd_sc_hd__or2_1
XFILLER_0_208_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09701_ hold3099/X _16391_/Q _10004_/C vssd1 vssd1 vccd1 vccd1 _09702_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07893_ hold2697/X _07918_/B _07892_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _07893_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09632_ hold1797/X _16368_/Q _11171_/C vssd1 vssd1 vccd1 vccd1 _09633_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_65_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09563_ hold645/X _13230_/A _10385_/S vssd1 vssd1 vccd1 vccd1 _09564_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_194_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08514_ hold2335/X _08503_/Y _08513_/X _13417_/C1 vssd1 vssd1 vccd1 vccd1 _08514_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09494_ _09494_/A _13055_/C _09494_/C vssd1 vssd1 vccd1 vccd1 _09494_/X sky130_fd_sc_hd__or3_4
XFILLER_0_147_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08445_ _14732_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08445_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_253_wb_clk_i clkbuf_6_59_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18200_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_114_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08376_ hold220/X _15820_/Q hold115/X vssd1 vssd1 vccd1 vccd1 hold221/A sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5620 _17091_/Q vssd1 vssd1 vccd1 vccd1 hold5620/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5631 _16751_/Q vssd1 vssd1 vccd1 vccd1 hold5631/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5642 _12115_/X vssd1 vssd1 vccd1 vccd1 _17195_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5653 _16901_/Q vssd1 vssd1 vccd1 vccd1 hold5653/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5664 _11632_/X vssd1 vssd1 vccd1 vccd1 _17034_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4930 _11104_/X vssd1 vssd1 vccd1 vccd1 _16858_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5675 _17235_/Q vssd1 vssd1 vccd1 vccd1 hold5675/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5686 _11689_/X vssd1 vssd1 vccd1 vccd1 _17053_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4941 _17025_/Q vssd1 vssd1 vccd1 vccd1 hold4941/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4952 _11674_/X vssd1 vssd1 vccd1 vccd1 _17048_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5697 _17129_/Q vssd1 vssd1 vccd1 vccd1 hold5697/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4963 _17592_/Q vssd1 vssd1 vccd1 vccd1 hold4963/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4974 _16402_/Q vssd1 vssd1 vccd1 vccd1 hold4974/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4985 _17607_/Q vssd1 vssd1 vccd1 vccd1 hold4985/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4996 _10753_/X vssd1 vssd1 vccd1 vccd1 _16741_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout430 _13267_/S vssd1 vssd1 vccd1 vccd1 _13307_/S sky130_fd_sc_hd__buf_12
Xfanout441 _13766_/S vssd1 vssd1 vccd1 vccd1 _13829_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout452 fanout485/X vssd1 vssd1 vccd1 vccd1 _11723_/C sky130_fd_sc_hd__clkbuf_4
Xfanout463 _12332_/C vssd1 vssd1 vccd1 vccd1 _13463_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_219_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_217_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout474 _11783_/C vssd1 vssd1 vccd1 vccd1 _12242_/S sky130_fd_sc_hd__clkbuf_8
Xfanout485 _09499_/Y vssd1 vssd1 vccd1 vccd1 fanout485/X sky130_fd_sc_hd__clkbuf_16
Xfanout496 _10964_/S vssd1 vssd1 vccd1 vccd1 _10025_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12910_ hold1690/X hold3334/X _12916_/S vssd1 vssd1 vccd1 vccd1 _12910_/X sky130_fd_sc_hd__mux2_1
X_13890_ _14556_/A hold1119/X _09120_/Y hold1391/X vssd1 vssd1 vccd1 vccd1 _13890_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_216_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12841_ hold1708/X _17458_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12841_/X sky130_fd_sc_hd__mux2_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ hold1643/X _15560_/A2 _15559_/X _12849_/A vssd1 vssd1 vccd1 vccd1 _15560_/X
+ sky130_fd_sc_hd__o211a_1
X_12772_ _16203_/Q hold3530/X _12838_/S vssd1 vssd1 vccd1 vccd1 _12772_/X sky130_fd_sc_hd__mux2_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14511_ _15191_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14511_/X sky130_fd_sc_hd__or2_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11723_ _17065_/Q _11723_/B _11723_/C vssd1 vssd1 vccd1 vccd1 _11723_/X sky130_fd_sc_hd__and3_1
X_15491_ _15491_/A _15491_/B vssd1 vssd1 vccd1 vccd1 _18425_/D sky130_fd_sc_hd__and2_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17900_/CLK _17230_/D vssd1 vssd1 vccd1 vccd1 _17230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ hold3023/X _14433_/B _14441_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _14442_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_232_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11654_ hold2487/X _17042_/Q _11654_/S vssd1 vssd1 vccd1 vccd1 _11655_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10605_ _16532_/Q _10413_/A _10604_/X vssd1 vssd1 vccd1 vccd1 _10605_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17161_ _17161_/CLK _17161_/D vssd1 vssd1 vccd1 vccd1 _17161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14373_ hold384/X hold783/X _14381_/S vssd1 vssd1 vccd1 vccd1 hold784/A sky130_fd_sc_hd__mux2_1
XFILLER_0_52_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11585_ hold2607/X _17019_/Q _12317_/C vssd1 vssd1 vccd1 vccd1 _11586_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16112_ _17335_/CLK _16112_/D vssd1 vssd1 vccd1 vccd1 _16112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13324_ hold5813/X _13808_/B _13323_/X _13417_/C1 vssd1 vssd1 vccd1 vccd1 _13324_/X
+ sky130_fd_sc_hd__o211a_1
X_10536_ _10536_/A _10536_/B vssd1 vssd1 vccd1 vccd1 _10536_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17092_ _17093_/CLK _17092_/D vssd1 vssd1 vccd1 vccd1 _17092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16043_ _18416_/CLK _16043_/D vssd1 vssd1 vccd1 vccd1 hold656/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13255_ _13311_/A1 _13253_/X _13254_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13255_/X
+ sky130_fd_sc_hd__o211a_1
X_10467_ _10476_/A _10467_/B vssd1 vssd1 vccd1 vccd1 _10467_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12206_ hold1664/X hold4811/X _12293_/C vssd1 vssd1 vccd1 vccd1 _12207_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_122_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_57_wb_clk_i clkbuf_6_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17983_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13186_ _17574_/Q _17108_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13186_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_209_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10398_ _10470_/A _10398_/B vssd1 vssd1 vccd1 vccd1 _10398_/X sky130_fd_sc_hd__or2_1
X_12137_ hold1562/X hold5671/X _12242_/S vssd1 vssd1 vccd1 vccd1 _12138_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17994_ _18024_/CLK _17994_/D vssd1 vssd1 vccd1 vccd1 _17994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12068_ hold2691/X hold4695/X _13481_/S vssd1 vssd1 vccd1 vccd1 _12069_/B sky130_fd_sc_hd__mux2_1
X_16945_ _17890_/CLK _16945_/D vssd1 vssd1 vccd1 vccd1 _16945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11019_ _11658_/A _11019_/B vssd1 vssd1 vccd1 vccd1 _11019_/X sky130_fd_sc_hd__or2_1
X_16876_ _17983_/CLK _16876_/D vssd1 vssd1 vccd1 vccd1 _16876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827_ _17738_/CLK _15827_/D vssd1 vssd1 vccd1 vccd1 hold940/A sky130_fd_sc_hd__dfxtp_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_231_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15758_ _17709_/CLK _15758_/D vssd1 vssd1 vccd1 vccd1 _15758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14709_ hold1986/X _14720_/B _14708_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _14709_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15689_ _17236_/CLK _15689_/D vssd1 vssd1 vccd1 vccd1 _15689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08230_ _14395_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08230_/X sky130_fd_sc_hd__or2_1
XFILLER_0_185_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17428_ _17429_/CLK _17428_/D vssd1 vssd1 vccd1 vccd1 _17428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08161_ _08163_/A _08161_/B vssd1 vssd1 vccd1 vccd1 _15718_/D sky130_fd_sc_hd__and2_1
X_17359_ _17380_/CLK _17359_/D vssd1 vssd1 vccd1 vccd1 _17359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08092_ _14330_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08092_/X sky130_fd_sc_hd__or2_1
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4204 _15423_/X vssd1 vssd1 vccd1 vccd1 _15424_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4215 hold5940/X vssd1 vssd1 vccd1 vccd1 hold5941/A sky130_fd_sc_hd__buf_6
Xhold4226 _10629_/Y vssd1 vssd1 vccd1 vccd1 _10630_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4237 _09999_/Y vssd1 vssd1 vccd1 vccd1 _10000_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3503 _16538_/Q vssd1 vssd1 vccd1 vccd1 hold3503/X sky130_fd_sc_hd__buf_1
Xhold4248 _17108_/Q vssd1 vssd1 vccd1 vccd1 hold4248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4259 _16715_/Q vssd1 vssd1 vccd1 vccd1 hold4259/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3514 _11212_/Y vssd1 vssd1 vccd1 vccd1 _16894_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3525 _16491_/Q vssd1 vssd1 vccd1 vccd1 hold3525/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_167_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3536 _16433_/Q vssd1 vssd1 vccd1 vccd1 hold3536/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2802 _18449_/Q vssd1 vssd1 vccd1 vccd1 hold2802/X sky130_fd_sc_hd__dlygate4sd3_1
X_08994_ _12394_/A hold503/X vssd1 vssd1 vccd1 vccd1 _16114_/D sky130_fd_sc_hd__and2_1
Xhold3547 _17586_/Q vssd1 vssd1 vccd1 vccd1 hold3547/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3558 _16590_/Q vssd1 vssd1 vccd1 vccd1 hold3558/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2813 _17967_/Q vssd1 vssd1 vccd1 vccd1 hold2813/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2824 _18097_/Q vssd1 vssd1 vccd1 vccd1 hold2824/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3569 _10516_/X vssd1 vssd1 vccd1 vccd1 _16662_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_167_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2835 _09300_/X vssd1 vssd1 vccd1 vccd1 _16260_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2846 _16266_/Q vssd1 vssd1 vccd1 vccd1 hold2846/X sky130_fd_sc_hd__dlygate4sd3_1
X_07945_ hold3041/X _07978_/B _07944_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _07945_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2857 _15788_/Q vssd1 vssd1 vccd1 vccd1 hold2857/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2868 _14761_/X vssd1 vssd1 vccd1 vccd1 _18171_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_6_2_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
Xhold2879 _18197_/Q vssd1 vssd1 vccd1 vccd1 hold2879/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07876_ hold2714/X _07869_/B _07875_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _07876_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09615_ _11067_/A _09615_/B vssd1 vssd1 vccd1 vccd1 _09615_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_434_wb_clk_i clkbuf_6_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17718_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_214_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09546_ _09912_/A _09546_/B vssd1 vssd1 vccd1 vccd1 _09546_/X sky130_fd_sc_hd__or2_1
XFILLER_0_190_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09477_ _09477_/A _09477_/B _09477_/C vssd1 vssd1 vccd1 vccd1 _09483_/C sky130_fd_sc_hd__and3_1
XFILLER_0_210_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08428_ hold2922/X _08433_/B _08427_/Y _08389_/A vssd1 vssd1 vccd1 vccd1 _08428_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08359_ _12750_/A _08359_/B vssd1 vssd1 vccd1 vccd1 _15811_/D sky130_fd_sc_hd__and2_1
XFILLER_0_151_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11370_ _11658_/A _11370_/B vssd1 vssd1 vccd1 vccd1 _11370_/X sky130_fd_sc_hd__or2_1
XFILLER_0_225_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10321_ hold3345/X _10589_/B _10320_/X _14691_/C1 vssd1 vssd1 vccd1 vccd1 _10321_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5450 _16752_/Q vssd1 vssd1 vccd1 vccd1 hold5450/X sky130_fd_sc_hd__dlygate4sd3_1
X_13040_ input2/X hold899/X hold920/X hold892/X vssd1 vssd1 vccd1 vccd1 hold921/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_123_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10252_ hold4493/X _10628_/B _10251_/X _14697_/C1 vssd1 vssd1 vccd1 vccd1 _10252_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5461 _13588_/X vssd1 vssd1 vccd1 vccd1 _17649_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5472 _17609_/Q vssd1 vssd1 vccd1 vccd1 hold5472/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5483 _13693_/X vssd1 vssd1 vccd1 vccd1 _17684_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5494 _17684_/Q vssd1 vssd1 vccd1 vccd1 hold5494/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4760 _17510_/Q vssd1 vssd1 vccd1 vccd1 hold4760/X sky130_fd_sc_hd__dlygate4sd3_1
X_10183_ hold3664/X _10625_/B _10182_/X _14769_/C1 vssd1 vssd1 vccd1 vccd1 _10183_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4771 _17667_/Q vssd1 vssd1 vccd1 vccd1 hold4771/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4782 _13318_/X vssd1 vssd1 vccd1 vccd1 _17559_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4793 _17191_/Q vssd1 vssd1 vccd1 vccd1 hold4793/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14991_ hold1797/X hold447/X _14990_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _14991_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout260 _11622_/A vssd1 vssd1 vccd1 vccd1 _12210_/A sky130_fd_sc_hd__buf_4
Xfanout271 fanout299/X vssd1 vssd1 vccd1 vccd1 _11556_/A sky130_fd_sc_hd__clkbuf_4
Xfanout282 fanout299/X vssd1 vssd1 vccd1 vccd1 _13599_/A sky130_fd_sc_hd__buf_2
XFILLER_0_156_1226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16730_ _18005_/CLK _16730_/D vssd1 vssd1 vccd1 vccd1 _16730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13942_ _14443_/A hold1613/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13943_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_89_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout293 _11697_/A vssd1 vssd1 vccd1 vccd1 _12240_/A sky130_fd_sc_hd__buf_4
XFILLER_0_96_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16661_ _18227_/CLK _16661_/D vssd1 vssd1 vccd1 vccd1 _16661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13873_ _13873_/A _13873_/B vssd1 vssd1 vccd1 vccd1 _13873_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_175_wb_clk_i clkbuf_6_49_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18383_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18400_ _18400_/CLK _18400_/D vssd1 vssd1 vccd1 vccd1 _18400_/Q sky130_fd_sc_hd__dfxtp_1
X_15612_ _17259_/CLK _15612_/D vssd1 vssd1 vccd1 vccd1 _15612_/Q sky130_fd_sc_hd__dfxtp_1
X_12824_ hold3127/X _12823_/X _12851_/S vssd1 vssd1 vccd1 vccd1 _12824_/X sky130_fd_sc_hd__mux2_1
X_16592_ _18150_/CLK _16592_/D vssd1 vssd1 vccd1 vccd1 _16592_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_104_wb_clk_i clkbuf_6_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17293_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18331_ _18363_/CLK _18331_/D vssd1 vssd1 vccd1 vccd1 _18331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15543_ _15543_/A _15547_/B vssd1 vssd1 vccd1 vccd1 _15543_/Y sky130_fd_sc_hd__nand2_1
X_12755_ hold3394/X _12754_/X _12812_/S vssd1 vssd1 vccd1 vccd1 _12755_/X sky130_fd_sc_hd__mux2_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18262_ _18262_/CLK _18262_/D vssd1 vssd1 vccd1 vccd1 _18262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _12240_/A _11706_/B vssd1 vssd1 vccd1 vccd1 _11706_/X sky130_fd_sc_hd__or2_1
X_15474_ hold602/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15474_/X sky130_fd_sc_hd__or2_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ hold3372/X _12685_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12687_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_154_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14425_ _15539_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14425_/X sky130_fd_sc_hd__or2_1
XFILLER_0_53_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17213_ _17277_/CLK _17213_/D vssd1 vssd1 vccd1 vccd1 _17213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18193_ _18225_/CLK _18193_/D vssd1 vssd1 vccd1 vccd1 _18193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11637_ _11637_/A _11637_/B vssd1 vssd1 vccd1 vccd1 _11637_/X sky130_fd_sc_hd__or2_1
XFILLER_0_155_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17144_ _17144_/CLK _17144_/D vssd1 vssd1 vccd1 vccd1 _17144_/Q sky130_fd_sc_hd__dfxtp_1
X_14356_ _14356_/A _14356_/B vssd1 vssd1 vccd1 vccd1 _17977_/D sky130_fd_sc_hd__and2_1
XFILLER_0_135_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11568_ _11670_/A _11568_/B vssd1 vssd1 vccd1 vccd1 _11568_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold708 hold819/X vssd1 vssd1 vccd1 vccd1 hold820/A sky130_fd_sc_hd__buf_6
X_13307_ _13306_/X hold5988/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13307_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10519_ hold3852/X _10631_/B _10518_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10519_/X
+ sky130_fd_sc_hd__o211a_1
Xhold719 hold719/A vssd1 vssd1 vccd1 vccd1 hold719/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17075_ _17891_/CLK _17075_/D vssd1 vssd1 vccd1 vccd1 _17075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14287_ hold445/X _14502_/B vssd1 vssd1 vccd1 vccd1 _14334_/B sky130_fd_sc_hd__or2_4
X_11499_ _11667_/A _11499_/B vssd1 vssd1 vccd1 vccd1 _11499_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16026_ _16026_/CLK _16026_/D vssd1 vssd1 vccd1 vccd1 hold863/A sky130_fd_sc_hd__dfxtp_1
X_13238_ _13238_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13238_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13169_ _13169_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13169_/X sky130_fd_sc_hd__and2_1
XFILLER_0_237_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2109 _18009_/Q vssd1 vssd1 vccd1 vccd1 hold2109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17977_ _18041_/CLK _17977_/D vssd1 vssd1 vccd1 vccd1 _17977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1408 _14478_/X vssd1 vssd1 vccd1 vccd1 _18036_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1419 _09439_/X vssd1 vssd1 vccd1 vccd1 _16305_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16928_ _17840_/CLK _16928_/D vssd1 vssd1 vccd1 vccd1 _16928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16859_ _18347_/CLK _16859_/D vssd1 vssd1 vccd1 vccd1 _16859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09400_ _09400_/A _09400_/B _09400_/C vssd1 vssd1 vccd1 vccd1 _09401_/S sky130_fd_sc_hd__or3_1
XFILLER_0_149_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09331_ _15173_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09331_/X sky130_fd_sc_hd__or2_1
XFILLER_0_192_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09262_ _12738_/A _09262_/B vssd1 vssd1 vccd1 vccd1 _16242_/D sky130_fd_sc_hd__and2_1
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08213_ _15221_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08213_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09193_ hold2462/X _09214_/B _09192_/X _12798_/A vssd1 vssd1 vccd1 vccd1 _09193_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08144_ _15549_/A hold1329/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08145_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_31_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08075_ hold2783/X _08097_/A2 _08074_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _08075_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4001 _16654_/Q vssd1 vssd1 vccd1 vccd1 hold4001/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4012 _11863_/X vssd1 vssd1 vccd1 vccd1 _17111_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4023 _11806_/X vssd1 vssd1 vccd1 vccd1 _17092_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4034 _16405_/Q vssd1 vssd1 vccd1 vccd1 hold4034/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4045 _12247_/X vssd1 vssd1 vccd1 vccd1 _17239_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3300 _17466_/Q vssd1 vssd1 vccd1 vccd1 hold3300/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3311 _10966_/X vssd1 vssd1 vccd1 vccd1 _16812_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4056 _16762_/Q vssd1 vssd1 vccd1 vccd1 hold4056/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3322 _16575_/Q vssd1 vssd1 vccd1 vccd1 hold3322/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4067 _13423_/X vssd1 vssd1 vccd1 vccd1 _17594_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4078 _13369_/X vssd1 vssd1 vccd1 vccd1 _17576_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3333 _12908_/X vssd1 vssd1 vccd1 vccd1 _12909_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3344 _12647_/X vssd1 vssd1 vccd1 vccd1 _12648_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4089 _16993_/Q vssd1 vssd1 vccd1 vccd1 hold4089/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3355 _17483_/Q vssd1 vssd1 vccd1 vccd1 hold3355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2610 _14201_/X vssd1 vssd1 vccd1 vccd1 _17903_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2621 _14881_/X vssd1 vssd1 vccd1 vccd1 _18229_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3366 _17457_/Q vssd1 vssd1 vccd1 vccd1 hold3366/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ hold373/X hold398/X _08991_/S vssd1 vssd1 vccd1 vccd1 _08978_/B sky130_fd_sc_hd__mux2_1
XTAP_5539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2632 _15110_/X vssd1 vssd1 vccd1 vccd1 _18339_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3377 _17452_/Q vssd1 vssd1 vccd1 vccd1 hold3377/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__buf_2
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2643 _18130_/Q vssd1 vssd1 vccd1 vccd1 hold2643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3388 _09394_/X vssd1 vssd1 vccd1 vccd1 _09395_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3399 _17369_/Q vssd1 vssd1 vccd1 vccd1 hold3399/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2654 _15713_/Q vssd1 vssd1 vccd1 vccd1 hold2654/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1920 _14759_/X vssd1 vssd1 vccd1 vccd1 _18170_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2665 _14801_/X vssd1 vssd1 vccd1 vccd1 _18190_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_6_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18458_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2676 _15228_/X vssd1 vssd1 vccd1 vccd1 _18396_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1931 _16164_/Q vssd1 vssd1 vccd1 vccd1 hold1931/X sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ hold992/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07928_/X sky130_fd_sc_hd__or2_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__buf_6
Xhold1942 _15076_/X vssd1 vssd1 vccd1 vccd1 _18322_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2687 _15753_/Q vssd1 vssd1 vccd1 vccd1 hold2687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1953 _15652_/Q vssd1 vssd1 vccd1 vccd1 hold1953/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2698 _07893_/X vssd1 vssd1 vccd1 vccd1 _15590_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1964 _18016_/Q vssd1 vssd1 vccd1 vccd1 hold1964/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1975 _09111_/X vssd1 vssd1 vccd1 vccd1 _16170_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1986 _18146_/Q vssd1 vssd1 vccd1 vccd1 hold1986/X sky130_fd_sc_hd__dlygate4sd3_1
X_07859_ _15537_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07859_/X sky130_fd_sc_hd__or2_1
XFILLER_0_224_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1997 _09314_/X vssd1 vssd1 vccd1 vccd1 _16267_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10870_ hold5010/X _11153_/B _10869_/X _14552_/C1 vssd1 vssd1 vccd1 vccd1 _10870_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_196_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09529_ hold4591/X _10031_/B _09528_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09529_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _12948_/A _12540_/B vssd1 vssd1 vccd1 vccd1 _17356_/D sky130_fd_sc_hd__and2_1
XFILLER_0_108_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12471_ hold77/X _12445_/A _12445_/B _12470_/X _15254_/A vssd1 vssd1 vccd1 vccd1
+ hold78/A sky130_fd_sc_hd__o311a_1
XFILLER_0_191_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14210_ _15555_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14210_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11422_ hold4050/X _12317_/B _11421_/X _14211_/C1 vssd1 vssd1 vccd1 vccd1 _11422_/X
+ sky130_fd_sc_hd__o211a_1
X_15190_ hold3186/X _15221_/B _15189_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _15190_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14141_ hold1718/X _14142_/B _14140_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _14141_/X
+ sky130_fd_sc_hd__o211a_1
X_11353_ hold5599/X _11744_/B _11352_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _11353_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10304_ hold2302/X _16592_/Q _10634_/C vssd1 vssd1 vccd1 vccd1 _10305_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14072_ _15145_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14072_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11284_ hold5012/X _11195_/B _11283_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _11284_/X
+ sky130_fd_sc_hd__o211a_1
X_13023_ hold937/X hold904/A vssd1 vssd1 vccd1 vccd1 _13025_/B sky130_fd_sc_hd__or2_1
XFILLER_0_120_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17900_ _17900_/CLK _17900_/D vssd1 vssd1 vccd1 vccd1 _17900_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5280 _10825_/X vssd1 vssd1 vccd1 vccd1 _16765_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10235_ hold1732/X _16569_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10236_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5291 _17082_/Q vssd1 vssd1 vccd1 vccd1 hold5291/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4590 _13630_/X vssd1 vssd1 vccd1 vccd1 _17663_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17831_ _17831_/CLK _17831_/D vssd1 vssd1 vccd1 vccd1 _17831_/Q sky130_fd_sc_hd__dfxtp_1
X_10166_ hold2652/X hold4245/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10167_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_233_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_356_wb_clk_i clkbuf_6_41_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17617_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17762_ _17859_/CLK _17762_/D vssd1 vssd1 vccd1 vccd1 hold971/A sky130_fd_sc_hd__dfxtp_1
X_10097_ hold1947/X _16523_/Q _10385_/S vssd1 vssd1 vccd1 vccd1 _10098_/B sky130_fd_sc_hd__mux2_1
X_14974_ _14974_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14974_/X sky130_fd_sc_hd__or2_1
XFILLER_0_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16713_ _18014_/CLK _16713_/D vssd1 vssd1 vccd1 vccd1 _16713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13925_ _13925_/A _13925_/B vssd1 vssd1 vccd1 vccd1 _17770_/D sky130_fd_sc_hd__and2_1
X_17693_ _17725_/CLK _17693_/D vssd1 vssd1 vccd1 vccd1 _17693_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_33_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_33_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_173_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16644_ _18234_/CLK _16644_/D vssd1 vssd1 vccd1 vccd1 _16644_/Q sky130_fd_sc_hd__dfxtp_1
X_13856_ _17739_/Q _13856_/B _13871_/C vssd1 vssd1 vccd1 vccd1 _13856_/X sky130_fd_sc_hd__and3_1
XFILLER_0_202_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12807_ _12810_/A _12807_/B vssd1 vssd1 vccd1 vccd1 _17445_/D sky130_fd_sc_hd__and2_1
XFILLER_0_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16575_ _18197_/CLK _16575_/D vssd1 vssd1 vccd1 vccd1 _16575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13787_ hold1489/X hold5482/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13788_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10999_ hold5070/X _10616_/B _10998_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _10999_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18314_ _18325_/CLK _18314_/D vssd1 vssd1 vccd1 vccd1 hold788/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _12738_/A _12738_/B vssd1 vssd1 vccd1 vccd1 _17422_/D sky130_fd_sc_hd__and2_1
XFILLER_0_45_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15526_ hold3089/X _15547_/B _15525_/X _12849_/A vssd1 vssd1 vccd1 vccd1 _15526_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15457_ hold556/X _09392_/C _09386_/D hold504/X _15456_/X vssd1 vssd1 vccd1 vccd1
+ _15462_/B sky130_fd_sc_hd__a221o_1
X_18245_ _18368_/CLK _18245_/D vssd1 vssd1 vccd1 vccd1 _18245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12669_ _12873_/A _12669_/B vssd1 vssd1 vccd1 vccd1 _17399_/D sky130_fd_sc_hd__and2_1
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14408_ hold2997/X _14446_/A2 _14407_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14408_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15388_ hold868/X _09386_/A _09392_/D hold770/X vssd1 vssd1 vccd1 vccd1 _15388_/X
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_72_wb_clk_i clkbuf_6_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18042_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18176_ _18176_/CLK _18176_/D vssd1 vssd1 vccd1 vccd1 _18176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14339_ hold1159/X _14326_/B _14338_/X _14528_/C1 vssd1 vssd1 vccd1 vccd1 _14339_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17127_ _17127_/CLK _17127_/D vssd1 vssd1 vccd1 vccd1 _17127_/Q sky130_fd_sc_hd__dfxtp_1
Xhold505 hold505/A vssd1 vssd1 vccd1 vccd1 hold505/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold516 hold516/A vssd1 vssd1 vccd1 vccd1 hold516/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 hold527/A vssd1 vssd1 vccd1 vccd1 hold527/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold538 hold538/A vssd1 vssd1 vccd1 vccd1 hold538/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17058_ _17906_/CLK _17058_/D vssd1 vssd1 vccd1 vccd1 _17058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold549 hold578/X vssd1 vssd1 vccd1 vccd1 hold579/A sky130_fd_sc_hd__buf_6
XFILLER_0_110_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16009_ _18416_/CLK _16009_/D vssd1 vssd1 vccd1 vccd1 hold611/A sky130_fd_sc_hd__dfxtp_1
X_08900_ hold180/X hold728/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold729/A sky130_fd_sc_hd__mux2_1
X_09880_ hold4662/X _10070_/B _09879_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _09880_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _15324_/A hold380/X vssd1 vssd1 vccd1 vccd1 _16034_/D sky130_fd_sc_hd__and2_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1205 _15572_/Q vssd1 vssd1 vccd1 vccd1 hold1205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 _08334_/X vssd1 vssd1 vccd1 vccd1 _15800_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08762_ _09440_/B hold700/X vssd1 vssd1 vccd1 vccd1 _16001_/D sky130_fd_sc_hd__and2_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 _15848_/Q vssd1 vssd1 vccd1 vccd1 hold1227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1238 _17780_/Q vssd1 vssd1 vccd1 vccd1 hold1238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 _09203_/X vssd1 vssd1 vccd1 vccd1 _16213_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_164_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_217_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08693_ hold172/X hold832/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08694_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09314_ hold1996/X _09323_/B _09313_/X _14358_/A vssd1 vssd1 vccd1 vccd1 _09314_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09245_ _15521_/A hold2337/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09246_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09176_ _15559_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09176_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08127_ _08135_/A _08127_/B vssd1 vssd1 vccd1 vccd1 _15702_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08058_ _15517_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08058_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3130 _07798_/X vssd1 vssd1 vccd1 vccd1 _07799_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10020_ _13166_/A _09933_/A _10019_/X vssd1 vssd1 vccd1 vccd1 _10020_/Y sky130_fd_sc_hd__a21oi_1
Xhold3141 _17478_/Q vssd1 vssd1 vccd1 vccd1 hold3141/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3152 _17470_/Q vssd1 vssd1 vccd1 vccd1 hold3152/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3163 _18084_/Q vssd1 vssd1 vccd1 vccd1 hold3163/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3174 _12743_/X vssd1 vssd1 vccd1 vccd1 _12744_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3185 _15136_/X vssd1 vssd1 vccd1 vccd1 _18351_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2440 _07868_/X vssd1 vssd1 vccd1 vccd1 _15579_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2451 _15847_/Q vssd1 vssd1 vccd1 vccd1 hold2451/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3196 _10062_/Y vssd1 vssd1 vccd1 vccd1 _10063_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2462 _16208_/Q vssd1 vssd1 vccd1 vccd1 hold2462/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2473 _15546_/X vssd1 vssd1 vccd1 vccd1 _18451_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2484 _14853_/X vssd1 vssd1 vccd1 vccd1 _18215_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1750 _18209_/Q vssd1 vssd1 vccd1 vccd1 hold1750/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2495 _16272_/Q vssd1 vssd1 vccd1 vccd1 hold2495/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1761 _08479_/X vssd1 vssd1 vccd1 vccd1 _15868_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ hold4927/X _12353_/B _11970_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _11971_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1772 _17985_/Q vssd1 vssd1 vccd1 vccd1 hold1772/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1783 _17795_/Q vssd1 vssd1 vccd1 vccd1 hold1783/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1794 _08261_/X vssd1 vssd1 vccd1 vccd1 _15765_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13710_ _13719_/A _13710_/B vssd1 vssd1 vccd1 vccd1 _13710_/X sky130_fd_sc_hd__or2_1
XFILLER_0_233_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10922_ hold2707/X hold4081/X _11210_/C vssd1 vssd1 vccd1 vccd1 _10923_/B sky130_fd_sc_hd__mux2_1
X_14690_ _15191_/A _14730_/B vssd1 vssd1 vccd1 vccd1 _14690_/X sky130_fd_sc_hd__or2_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13641_ _13737_/A _13641_/B vssd1 vssd1 vccd1 vccd1 _13641_/X sky130_fd_sc_hd__or2_1
X_10853_ hold3067/X hold3842/X _11144_/C vssd1 vssd1 vccd1 vccd1 _10854_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_211_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _18373_/CLK _16360_/D vssd1 vssd1 vccd1 vccd1 _16360_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13572_ _13752_/A _13572_/B vssd1 vssd1 vccd1 vccd1 _13572_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10784_ hold1851/X _16752_/Q _11168_/C vssd1 vssd1 vccd1 vccd1 _10785_/B sky130_fd_sc_hd__mux2_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _09418_/B _09362_/A _09392_/B hold807/X _15310_/X vssd1 vssd1 vccd1 vccd1
+ _15312_/D sky130_fd_sc_hd__a221o_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12523_ hold2404/X hold3638/X _12925_/S vssd1 vssd1 vccd1 vccd1 _12523_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16291_ _18408_/CLK _16291_/D vssd1 vssd1 vccd1 vccd1 _16291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15242_ _15489_/A _15242_/B _15242_/C _15242_/D vssd1 vssd1 vccd1 vccd1 _15242_/X
+ sky130_fd_sc_hd__or4_1
X_18030_ _18030_/CLK _18030_/D vssd1 vssd1 vccd1 vccd1 _18030_/Q sky130_fd_sc_hd__dfxtp_1
X_12454_ _17320_/Q _12506_/B vssd1 vssd1 vccd1 vccd1 _12454_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11405_ hold1970/X hold4933/X _12173_/S vssd1 vssd1 vccd1 vccd1 _11406_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_112_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15173_ _15173_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15173_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12385_ hold131/X hold390/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold391/A sky130_fd_sc_hd__mux2_1
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14124_ _14517_/A _14140_/B vssd1 vssd1 vccd1 vccd1 _14124_/X sky130_fd_sc_hd__or2_1
X_11336_ hold3025/X _16936_/Q _12299_/C vssd1 vssd1 vccd1 vccd1 _11337_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14055_ _14735_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14106_/B sky130_fd_sc_hd__or2_4
X_11267_ hold2764/X hold4430/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11268_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13006_ hold1528/X _13003_/Y _13005_/X _12984_/A vssd1 vssd1 vccd1 vccd1 _13006_/X
+ sky130_fd_sc_hd__o211a_1
X_10218_ _10524_/A _10218_/B vssd1 vssd1 vccd1 vccd1 _10218_/X sky130_fd_sc_hd__or2_1
XTAP_6560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11198_ _16890_/Q _11213_/B _11219_/C vssd1 vssd1 vccd1 vccd1 _11198_/X sky130_fd_sc_hd__and3_1
XTAP_6571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_190_wb_clk_i clkbuf_6_52_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18381_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17814_ _17846_/CLK _17814_/D vssd1 vssd1 vccd1 vccd1 _17814_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10149_ _10515_/A _10149_/B vssd1 vssd1 vccd1 vccd1 _10149_/X sky130_fd_sc_hd__or2_1
XFILLER_0_234_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17745_ _17745_/CLK _17745_/D vssd1 vssd1 vccd1 vccd1 _17745_/Q sky130_fd_sc_hd__dfxtp_1
X_14957_ hold1907/X _14952_/B _14956_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _14957_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13908_ _14517_/A hold971/X hold297/X vssd1 vssd1 vccd1 vccd1 hold972/A sky130_fd_sc_hd__mux2_1
X_17676_ _17748_/CLK _17676_/D vssd1 vssd1 vccd1 vccd1 _17676_/Q sky130_fd_sc_hd__dfxtp_1
X_14888_ _15227_/A _14892_/B vssd1 vssd1 vccd1 vccd1 _14888_/X sky130_fd_sc_hd__or2_1
XFILLER_0_77_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16627_ _18223_/CLK _16627_/D vssd1 vssd1 vccd1 vccd1 _16627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13839_ hold4402/X _13773_/A _13838_/X vssd1 vssd1 vccd1 vccd1 _13839_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_230_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16558_ _18154_/CLK _16558_/D vssd1 vssd1 vccd1 vccd1 _16558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15509_ _15509_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15509_/X sky130_fd_sc_hd__or2_1
X_16489_ _18370_/CLK _16489_/D vssd1 vssd1 vccd1 vccd1 _16489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09030_ hold180/X _16132_/Q _09056_/S vssd1 vssd1 vccd1 vccd1 hold181/A sky130_fd_sc_hd__mux2_1
X_18228_ _18228_/CLK _18228_/D vssd1 vssd1 vccd1 vccd1 _18228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18159_ _18215_/CLK _18159_/D vssd1 vssd1 vccd1 vccd1 _18159_/Q sky130_fd_sc_hd__dfxtp_1
Xhold302 hold302/A vssd1 vssd1 vccd1 vccd1 hold302/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 hold34/X vssd1 vssd1 vccd1 vccd1 input23/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold324 hold324/A vssd1 vssd1 vccd1 vccd1 hold324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 hold335/A vssd1 vssd1 vccd1 vccd1 input57/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold346 hold346/A vssd1 vssd1 vccd1 vccd1 hold346/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold357 hold357/A vssd1 vssd1 vccd1 vccd1 hold357/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_278_wb_clk_i clkbuf_6_50_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18176_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09932_ hold1002/X hold4547/X _10028_/C vssd1 vssd1 vccd1 vccd1 _09933_/B sky130_fd_sc_hd__mux2_1
Xhold368 hold368/A vssd1 vssd1 vccd1 vccd1 hold368/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold379 hold379/A vssd1 vssd1 vccd1 vccd1 hold379/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_207_wb_clk_i clkbuf_6_55_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18262_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout804 _15066_/A vssd1 vssd1 vccd1 vccd1 _15048_/A sky130_fd_sc_hd__buf_4
XFILLER_0_102_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout815 fanout816/X vssd1 vssd1 vccd1 vccd1 _15204_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout826 _14863_/C1 vssd1 vssd1 vccd1 vccd1 _14390_/A sky130_fd_sc_hd__clkbuf_4
X_09863_ _18358_/Q hold3612/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09864_/B sky130_fd_sc_hd__mux2_1
Xfanout837 _14691_/C1 vssd1 vssd1 vccd1 vccd1 _14849_/C1 sky130_fd_sc_hd__buf_4
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout848 _17754_/Q vssd1 vssd1 vccd1 vccd1 _13888_/A sky130_fd_sc_hd__buf_8
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout859 hold5970/X vssd1 vssd1 vccd1 vccd1 _13312_/B1 sky130_fd_sc_hd__buf_8
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08814_ hold147/X hold863/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08815_/B sky130_fd_sc_hd__mux2_1
Xhold1002 _18381_/Q vssd1 vssd1 vccd1 vccd1 hold1002/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 _14589_/X vssd1 vssd1 vccd1 vccd1 _18088_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _18335_/Q hold4713/X _09992_/C vssd1 vssd1 vccd1 vccd1 _09795_/B sky130_fd_sc_hd__mux2_1
Xhold1024 _09183_/X vssd1 vssd1 vccd1 vccd1 _16203_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1035 _17832_/Q vssd1 vssd1 vccd1 vccd1 hold1035/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1046 _08418_/X vssd1 vssd1 vccd1 vccd1 _15839_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08745_ hold679/X hold870/X _08779_/S vssd1 vssd1 vccd1 vccd1 hold871/A sky130_fd_sc_hd__mux2_1
Xhold1057 _08093_/X vssd1 vssd1 vccd1 vccd1 _15686_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1068 _14446_/X vssd1 vssd1 vccd1 vccd1 _18021_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 _15714_/Q vssd1 vssd1 vccd1 vccd1 hold1079/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08676_ _12410_/A _08676_/B vssd1 vssd1 vccd1 vccd1 _15959_/D sky130_fd_sc_hd__and2_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09228_ _15557_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09228_/X sky130_fd_sc_hd__or2_1
XFILLER_0_17_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09159_ hold3021/X _09164_/B _09158_/Y _12906_/A vssd1 vssd1 vccd1 vccd1 _09159_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12170_ hold1323/X _17214_/Q _12362_/C vssd1 vssd1 vccd1 vccd1 _12171_/B sky130_fd_sc_hd__mux2_1
X_11121_ _11121_/A _11121_/B vssd1 vssd1 vccd1 vccd1 _11121_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold880 hold880/A vssd1 vssd1 vccd1 vccd1 hold880/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold891 becStatus[2] vssd1 vssd1 vccd1 vccd1 input3/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11052_ _11136_/A _11052_/B vssd1 vssd1 vccd1 vccd1 _11052_/X sky130_fd_sc_hd__or2_1
XTAP_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10003_ _11203_/A _10003_/B vssd1 vssd1 vccd1 vccd1 _10003_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_194_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15860_ _17648_/CLK _15860_/D vssd1 vssd1 vccd1 vccd1 _15860_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2270 input69/X vssd1 vssd1 vccd1 vccd1 hold2270/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14811_ hold2888/X _14826_/B _14810_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14811_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2281 _14565_/X vssd1 vssd1 vccd1 vccd1 _18077_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2292 _17974_/Q vssd1 vssd1 vccd1 vccd1 hold2292/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _17626_/CLK _15791_/D vssd1 vssd1 vccd1 vccd1 _15791_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1580 hold1580/A vssd1 vssd1 vccd1 vccd1 _14974_/A sky130_fd_sc_hd__buf_8
X_17530_ _17533_/CLK _17530_/D vssd1 vssd1 vccd1 vccd1 _17530_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14742_ _15189_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14742_/X sky130_fd_sc_hd__or2_1
Xhold1591 _07943_/X vssd1 vssd1 vccd1 vccd1 _15614_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11954_ hold2293/X _17142_/Q _12173_/S vssd1 vssd1 vccd1 vccd1 _11955_/B sky130_fd_sc_hd__mux2_1
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ _11694_/A _10905_/B vssd1 vssd1 vccd1 vccd1 _10905_/X sky130_fd_sc_hd__or2_1
X_14673_ hold2637/X _14664_/B _14672_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _14673_/X
+ sky130_fd_sc_hd__o211a_1
X_17461_ _17462_/CLK _17461_/D vssd1 vssd1 vccd1 vccd1 _17461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11885_ hold1329/X hold3496/X _13748_/S vssd1 vssd1 vccd1 vccd1 _11886_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16412_ _18357_/CLK _16412_/D vssd1 vssd1 vccd1 vccd1 _16412_/Q sky130_fd_sc_hd__dfxtp_1
X_13624_ hold5777/X _13808_/B _13623_/X _12753_/A vssd1 vssd1 vccd1 vccd1 _13624_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_1395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10836_ _11124_/A _10836_/B vssd1 vssd1 vccd1 vccd1 _10836_/X sky130_fd_sc_hd__or2_1
XFILLER_0_200_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17392_ _18445_/CLK _17392_/D vssd1 vssd1 vccd1 vccd1 _17392_/Q sky130_fd_sc_hd__dfxtp_1
X_16343_ _18392_/CLK _16343_/D vssd1 vssd1 vccd1 vccd1 _16343_/Q sky130_fd_sc_hd__dfxtp_1
X_13555_ hold5610/X _13847_/B _13554_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13555_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10767_ _11043_/A _10767_/B vssd1 vssd1 vccd1 vccd1 _10767_/X sky130_fd_sc_hd__or2_1
XFILLER_0_171_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12506_ _17346_/Q _12506_/B vssd1 vssd1 vccd1 vccd1 _12506_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16274_ _17378_/CLK _16274_/D vssd1 vssd1 vccd1 vccd1 _16274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ hold5351/X _13868_/B _13485_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _13486_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10698_ _11109_/A _10698_/B vssd1 vssd1 vccd1 vccd1 _10698_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15225_ _15225_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15225_/X sky130_fd_sc_hd__or2_1
X_18013_ _18013_/CLK _18013_/D vssd1 vssd1 vccd1 vccd1 _18013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12437_ hold87/X hold94/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__mux2_1
XFILLER_0_207_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15156_ hold2157/X _15167_/B _15155_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _15156_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12368_ _17280_/Q _13886_/B _13886_/C vssd1 vssd1 vccd1 vccd1 _12368_/X sky130_fd_sc_hd__and3_1
XFILLER_0_205_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_238_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_371_wb_clk_i clkbuf_6_32_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17648_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14107_ hold1010/X _14107_/A2 _14106_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _14107_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11319_ _12174_/A _11319_/B vssd1 vssd1 vccd1 vccd1 _11319_/X sky130_fd_sc_hd__or2_1
X_15087_ _15195_/A _15119_/B vssd1 vssd1 vccd1 vccd1 _15087_/X sky130_fd_sc_hd__or2_1
X_12299_ _17257_/Q _12299_/B _12299_/C vssd1 vssd1 vccd1 vccd1 _12299_/X sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_300_wb_clk_i clkbuf_6_38_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17894_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_201_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14038_ _15545_/A _14038_/B vssd1 vssd1 vccd1 vccd1 _14038_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_240_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15989_ _17321_/CLK _15989_/D vssd1 vssd1 vccd1 vccd1 hold823/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08530_ _13056_/C _17520_/Q _08868_/B vssd1 vssd1 vccd1 vccd1 _12380_/A sky130_fd_sc_hd__or3_1
XFILLER_0_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17728_ _17728_/CLK _17728_/D vssd1 vssd1 vccd1 vccd1 _17728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08461_ hold998/X _08488_/B _08460_/X _08367_/A vssd1 vssd1 vccd1 vccd1 hold999/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_216_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17659_ _17689_/CLK _17659_/D vssd1 vssd1 vccd1 vccd1 _17659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08392_ hold444/A hold405/A hold509/A hold337/A vssd1 vssd1 vccd1 vccd1 hold445/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_147_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_459_wb_clk_i clkbuf_6_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17430_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09013_ _09061_/A _09013_/B vssd1 vssd1 vccd1 vccd1 _16123_/D sky130_fd_sc_hd__and2_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5802 _13330_/X vssd1 vssd1 vccd1 vccd1 _17563_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5813 _17593_/Q vssd1 vssd1 vccd1 vccd1 hold5813/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5824 _09820_/X vssd1 vssd1 vccd1 vccd1 _16430_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5835 _16470_/Q vssd1 vssd1 vccd1 vccd1 hold5835/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold110 hold110/A vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 hold4/X vssd1 vssd1 vccd1 vccd1 input17/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5846 output86/X vssd1 vssd1 vccd1 vccd1 data_out[22] sky130_fd_sc_hd__buf_12
Xhold132 hold132/A vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5857 hold6013/X vssd1 vssd1 vccd1 vccd1 _13249_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5868 hold5868/A vssd1 vssd1 vccd1 vccd1 data_out[9] sky130_fd_sc_hd__buf_12
Xhold143 hold17/X vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__clkbuf_4
Xhold5879 hold6024/X vssd1 vssd1 vccd1 vccd1 _13193_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 hold154/A vssd1 vssd1 vccd1 vccd1 hold154/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 hold165/A vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 hold176/A vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_229_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold187 hold187/A vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _12871_/S vssd1 vssd1 vccd1 vccd1 _12970_/S sky130_fd_sc_hd__clkbuf_4
Xfanout612 _09362_/C vssd1 vssd1 vccd1 vccd1 _15486_/B1 sky130_fd_sc_hd__buf_6
Xhold198 hold286/X vssd1 vssd1 vccd1 vccd1 hold287/A sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _09981_/A _09915_/B vssd1 vssd1 vccd1 vccd1 _09915_/X sky130_fd_sc_hd__or2_1
Xfanout623 _09349_/Y vssd1 vssd1 vccd1 vccd1 _15485_/A2 sky130_fd_sc_hd__buf_8
Xfanout634 _12798_/A vssd1 vssd1 vccd1 vccd1 _12786_/A sky130_fd_sc_hd__clkbuf_4
Xfanout645 _12199_/C1 vssd1 vssd1 vccd1 vccd1 _12822_/A sky130_fd_sc_hd__buf_4
Xfanout656 fanout739/X vssd1 vssd1 vccd1 vccd1 _12597_/A sky130_fd_sc_hd__buf_2
XFILLER_0_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09846_ _09954_/A _09846_/B vssd1 vssd1 vccd1 vccd1 _09846_/X sky130_fd_sc_hd__or2_1
Xfanout667 _08171_/A vssd1 vssd1 vccd1 vccd1 _08167_/A sky130_fd_sc_hd__buf_4
Xfanout678 _15498_/A vssd1 vssd1 vccd1 vccd1 _15494_/A sky130_fd_sc_hd__buf_4
Xfanout689 fanout739/X vssd1 vssd1 vccd1 vccd1 fanout689/X sky130_fd_sc_hd__clkbuf_8
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _09978_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09777_/X sky130_fd_sc_hd__or2_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _09061_/A hold524/X vssd1 vssd1 vccd1 vccd1 _15985_/D sky130_fd_sc_hd__and2_1
XFILLER_0_197_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08659_ hold320/X hold868/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08660_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_166_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11670_ _11670_/A _11670_/B vssd1 vssd1 vccd1 vccd1 _11670_/X sky130_fd_sc_hd__or2_1
XFILLER_0_194_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10621_ _10651_/A _10621_/B vssd1 vssd1 vccd1 vccd1 _16697_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_187_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13340_ hold2983/X _17567_/Q _13766_/S vssd1 vssd1 vccd1 vccd1 _13341_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_221_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10552_ hold4632/X _10646_/B _10551_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _10552_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13271_ _13311_/A1 _13269_/X _13270_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13271_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_107_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10483_ hold3862/X _10577_/B _10482_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10483_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_224_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_129_wb_clk_i clkbuf_6_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17318_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15010_ _15225_/A hold510/A vssd1 vssd1 vccd1 vccd1 _15010_/X sky130_fd_sc_hd__or2_1
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12222_ _12285_/A _12222_/B vssd1 vssd1 vccd1 vccd1 _12222_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ _13749_/A _12153_/B vssd1 vssd1 vccd1 vccd1 _12153_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11104_ hold4929/X _11213_/B _11103_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _11104_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12084_ _13749_/A _12084_/B vssd1 vssd1 vccd1 vccd1 _12084_/X sky130_fd_sc_hd__or2_1
X_16961_ _17843_/CLK _16961_/D vssd1 vssd1 vccd1 vccd1 _16961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15912_ _17291_/CLK _15912_/D vssd1 vssd1 vccd1 vccd1 hold666/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11035_ hold4701/X _11765_/B _11034_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _11035_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16892_ _18031_/CLK _16892_/D vssd1 vssd1 vccd1 vccd1 _16892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ _17606_/CLK _15843_/D vssd1 vssd1 vccd1 vccd1 _15843_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ hold3748/X _12985_/X _12986_/S vssd1 vssd1 vccd1 vccd1 _12986_/X sky130_fd_sc_hd__mux2_1
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ _17661_/CLK _15774_/D vssd1 vssd1 vccd1 vccd1 _15774_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ _17513_/CLK _17513_/D vssd1 vssd1 vccd1 vccd1 _17513_/Q sky130_fd_sc_hd__dfxtp_1
X_14725_ hold1766/X _14720_/B _14724_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _14725_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ _13314_/A _11937_/B vssd1 vssd1 vccd1 vccd1 _11937_/X sky130_fd_sc_hd__or2_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _17725_/CLK _17444_/D vssd1 vssd1 vccd1 vccd1 _17444_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14656_ _15103_/A _14672_/B vssd1 vssd1 vccd1 vccd1 _14656_/X sky130_fd_sc_hd__or2_1
X_11868_ _12255_/A _11868_/B vssd1 vssd1 vccd1 vccd1 _11868_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10819_ hold5072/X _11171_/B _10818_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _10819_/X
+ sky130_fd_sc_hd__o211a_1
X_13607_ hold1841/X _17656_/Q _13721_/S vssd1 vssd1 vccd1 vccd1 _13608_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17375_ _17378_/CLK _17375_/D vssd1 vssd1 vccd1 vccd1 _17375_/Q sky130_fd_sc_hd__dfxtp_1
X_14587_ hold3033/X _14610_/B _14586_/X _14853_/C1 vssd1 vssd1 vccd1 vccd1 _14587_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11799_ hold4295/X _12174_/A _11798_/X vssd1 vssd1 vccd1 vccd1 _11799_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16326_ _18411_/CLK _16326_/D vssd1 vssd1 vccd1 vccd1 _16326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13538_ _15818_/Q hold4642/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13539_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16257_ _17360_/CLK _16257_/D vssd1 vssd1 vccd1 vccd1 _16257_/Q sky130_fd_sc_hd__dfxtp_1
X_13469_ hold2451/X hold5341/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13470_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5109 _16843_/Q vssd1 vssd1 vccd1 vccd1 hold5109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15208_ hold1434/X _15219_/B _15207_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _15208_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4408 _17579_/Q vssd1 vssd1 vccd1 vccd1 hold4408/X sky130_fd_sc_hd__dlygate4sd3_1
X_16188_ _17882_/CLK _16188_/D vssd1 vssd1 vccd1 vccd1 _16188_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4419 _16908_/Q vssd1 vssd1 vccd1 vccd1 hold4419/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15139_ _15193_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15139_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3707 _10087_/X vssd1 vssd1 vccd1 vccd1 _16519_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3718 _16891_/Q vssd1 vssd1 vccd1 vccd1 hold3718/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_107_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3729 _13603_/X vssd1 vssd1 vccd1 vccd1 _17654_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07961_ hold2859/X _07991_/A2 _07960_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _07961_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09700_ hold4713/X _09992_/B _09699_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _09700_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07892_ _14850_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07892_/X sky130_fd_sc_hd__or2_1
X_09631_ hold3734/X _10004_/B _09630_/X _15048_/A vssd1 vssd1 vccd1 vccd1 _09631_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09562_ hold3622/X _10052_/B _09561_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _09562_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08513_ _15517_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08513_/X sky130_fd_sc_hd__or2_1
XFILLER_0_195_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09493_ _09494_/A _13055_/C _09494_/C vssd1 vssd1 vccd1 vccd1 wire337/A sky130_fd_sc_hd__nor3_4
XFILLER_0_148_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08444_ hold1207/X _08433_/B _08443_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _08444_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08375_ _09272_/A hold614/X vssd1 vssd1 vccd1 vccd1 _15819_/D sky130_fd_sc_hd__and2_1
XFILLER_0_135_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_293_wb_clk_i clkbuf_6_39_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18053_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_222_wb_clk_i clkbuf_6_61_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18191_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5610 _17670_/Q vssd1 vssd1 vccd1 vccd1 hold5610/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5621 _11707_/X vssd1 vssd1 vccd1 vccd1 _17059_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5632 _10687_/X vssd1 vssd1 vccd1 vccd1 _16719_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5643 _17639_/Q vssd1 vssd1 vccd1 vccd1 hold5643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5654 _11713_/X vssd1 vssd1 vccd1 vccd1 _17061_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4920 _09658_/X vssd1 vssd1 vccd1 vccd1 _16376_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5665 _16989_/Q vssd1 vssd1 vccd1 vccd1 hold5665/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4931 _17126_/Q vssd1 vssd1 vccd1 vccd1 hold4931/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5676 _12139_/X vssd1 vssd1 vccd1 vccd1 _17203_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5687 _17193_/Q vssd1 vssd1 vccd1 vccd1 hold5687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4942 _11509_/X vssd1 vssd1 vccd1 vccd1 _16993_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5698 _11821_/X vssd1 vssd1 vccd1 vccd1 _17097_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4953 _17057_/Q vssd1 vssd1 vccd1 vccd1 hold4953/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4964 _13321_/X vssd1 vssd1 vccd1 vccd1 _17560_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_1394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4975 _09640_/X vssd1 vssd1 vccd1 vccd1 _16370_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4986 _13366_/X vssd1 vssd1 vccd1 vccd1 _17575_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout420 _14054_/Y vssd1 vssd1 vccd1 vccd1 _14107_/A2 sky130_fd_sc_hd__buf_6
Xfanout431 _13054_/X vssd1 vssd1 vccd1 vccd1 _13181_/S sky130_fd_sc_hd__clkbuf_16
Xhold4997 _16849_/Q vssd1 vssd1 vccd1 vccd1 hold4997/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout442 _13766_/S vssd1 vssd1 vccd1 vccd1 _13862_/C sky130_fd_sc_hd__clkbuf_8
Xfanout453 _11741_/C vssd1 vssd1 vccd1 vccd1 _12317_/C sky130_fd_sc_hd__clkbuf_8
Xfanout464 _13868_/C vssd1 vssd1 vccd1 vccd1 _12332_/C sky130_fd_sc_hd__buf_4
Xfanout475 fanout485/X vssd1 vssd1 vccd1 vccd1 _11783_/C sky130_fd_sc_hd__clkbuf_4
Xfanout486 _11144_/C vssd1 vssd1 vccd1 vccd1 _11153_/C sky130_fd_sc_hd__clkbuf_8
X_09829_ hold3566/X _10046_/B _09828_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _09829_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout497 _09499_/Y vssd1 vssd1 vccd1 vccd1 _10964_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_225_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ _12843_/A _12840_/B vssd1 vssd1 vccd1 vccd1 _17456_/D sky130_fd_sc_hd__and2_1
XFILLER_0_198_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_232_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12771_ _12777_/A _12771_/B vssd1 vssd1 vccd1 vccd1 _17433_/D sky130_fd_sc_hd__and2_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11722_ _12301_/A _11722_/B vssd1 vssd1 vccd1 vccd1 _17064_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_90_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14510_ hold2129/X _14537_/B _14509_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _14510_/X
+ sky130_fd_sc_hd__o211a_1
X_15490_ _15490_/A1 _15483_/X _15489_/X _15490_/B1 hold5974/A vssd1 vssd1 vccd1 vccd1
+ _15490_/X sky130_fd_sc_hd__a32o_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ hold5657/X _12323_/B _11652_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _11653_/X
+ sky130_fd_sc_hd__o211a_1
X_14441_ _15229_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14441_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10604_ _10604_/A _10604_/B _10604_/C vssd1 vssd1 vccd1 vccd1 _10604_/X sky130_fd_sc_hd__and3_1
XFILLER_0_181_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14372_ _14372_/A _14372_/B vssd1 vssd1 vccd1 vccd1 _17985_/D sky130_fd_sc_hd__and2_1
XFILLER_0_36_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17160_ _17628_/CLK _17160_/D vssd1 vssd1 vccd1 vccd1 _17160_/Q sky130_fd_sc_hd__dfxtp_1
X_11584_ hold5161/X _11771_/B _11583_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _11584_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16111_ _17314_/CLK _16111_/D vssd1 vssd1 vccd1 vccd1 hold858/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13323_ _13719_/A _13323_/B vssd1 vssd1 vccd1 vccd1 _13323_/X sky130_fd_sc_hd__or2_1
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10535_ hold1863/X hold3830/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10536_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17091_ _17907_/CLK _17091_/D vssd1 vssd1 vccd1 vccd1 _17091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16042_ _16098_/CLK _16042_/D vssd1 vssd1 vccd1 vccd1 hold633/A sky130_fd_sc_hd__dfxtp_1
X_13254_ _13254_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13254_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10466_ hold1064/X hold3720/X _10571_/C vssd1 vssd1 vccd1 vccd1 _10467_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_122_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12205_ hold5689/X _12299_/B _12204_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _12205_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13185_ _13185_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13185_/X sky130_fd_sc_hd__and2_1
X_10397_ hold2906/X _16623_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10398_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12136_ hold5803/X _12332_/B _12135_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _12136_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17993_ _18208_/CLK _17993_/D vssd1 vssd1 vccd1 vccd1 _17993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12067_ hold4815/X _12353_/B _12066_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _12067_/X
+ sky130_fd_sc_hd__o211a_1
X_16944_ _17888_/CLK _16944_/D vssd1 vssd1 vccd1 vccd1 _16944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_97_wb_clk_i clkbuf_6_22_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16082_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11018_ hold1523/X hold4147/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11019_/B sky130_fd_sc_hd__mux2_1
X_16875_ _18072_/CLK _16875_/D vssd1 vssd1 vccd1 vccd1 _16875_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_26_wb_clk_i clkbuf_6_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17378_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_189_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15826_ _17737_/CLK _15826_/D vssd1 vssd1 vccd1 vccd1 _15826_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15757_ _17748_/CLK _15757_/D vssd1 vssd1 vccd1 vccd1 _15757_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12969_ _12978_/A _12969_/B vssd1 vssd1 vccd1 vccd1 _17499_/D sky130_fd_sc_hd__and2_1
XFILLER_0_73_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14708_ _15209_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14708_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15688_ _17262_/CLK _15688_/D vssd1 vssd1 vccd1 vccd1 _15688_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17427_ _17427_/CLK _17427_/D vssd1 vssd1 vccd1 vccd1 _17427_/Q sky130_fd_sc_hd__dfxtp_1
X_14639_ hold2739/X _14666_/B _14638_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _14639_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08160_ _14166_/A hold1451/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08160_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_172_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17358_ _17360_/CLK _17358_/D vssd1 vssd1 vccd1 vccd1 _17358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16309_ _18408_/CLK _16309_/D vssd1 vssd1 vccd1 vccd1 _16309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08091_ hold1513/X _08088_/B _08090_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _08091_/X
+ sky130_fd_sc_hd__o211a_1
X_17289_ _17335_/CLK _17289_/D vssd1 vssd1 vccd1 vccd1 _17289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4205 hold5966/X vssd1 vssd1 vccd1 vccd1 hold5967/A sky130_fd_sc_hd__buf_6
XFILLER_0_80_1322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4216 _09385_/X vssd1 vssd1 vccd1 vccd1 _16281_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4227 _16545_/Q vssd1 vssd1 vccd1 vccd1 hold4227/X sky130_fd_sc_hd__buf_1
Xhold4238 hold6115/X vssd1 vssd1 vccd1 vccd1 hold4238/X sky130_fd_sc_hd__buf_1
Xhold3504 _10623_/Y vssd1 vssd1 vccd1 vccd1 _10624_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4249 _12333_/Y vssd1 vssd1 vccd1 vccd1 _12334_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3515 _16536_/Q vssd1 vssd1 vccd1 vccd1 hold3515/X sky130_fd_sc_hd__buf_1
Xhold3526 _09907_/X vssd1 vssd1 vccd1 vccd1 _16459_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08993_ hold495/X hold502/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold503/A sky130_fd_sc_hd__mux2_1
Xhold3537 _09733_/X vssd1 vssd1 vccd1 vccd1 _16401_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3548 _13878_/Y vssd1 vssd1 vccd1 vccd1 _13879_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2803 _15542_/X vssd1 vssd1 vccd1 vccd1 _18449_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3559 _10204_/X vssd1 vssd1 vccd1 vccd1 _16558_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2814 _14335_/X vssd1 vssd1 vccd1 vccd1 _17967_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2825 _14607_/X vssd1 vssd1 vccd1 vccd1 _18097_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07944_ _15513_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07944_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2836 _18168_/Q vssd1 vssd1 vccd1 vccd1 hold2836/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2847 _09312_/X vssd1 vssd1 vccd1 vccd1 _16266_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2858 _08310_/X vssd1 vssd1 vccd1 vccd1 _15788_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2869 _18234_/Q vssd1 vssd1 vccd1 vccd1 hold2869/X sky130_fd_sc_hd__dlygate4sd3_1
X_07875_ _14726_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07875_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09614_ _18275_/Q _16362_/Q _11162_/C vssd1 vssd1 vccd1 vccd1 _09615_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_223_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ hold3100/X _13182_/A _10025_/C vssd1 vssd1 vccd1 vccd1 _09546_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_214_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09476_ _09477_/B _09477_/C _09477_/A vssd1 vssd1 vccd1 vccd1 _09478_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08427_ _15215_/A _08433_/B vssd1 vssd1 vccd1 vccd1 _08427_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_403_wb_clk_i clkbuf_6_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18019_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_164_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08358_ hold951/X hold1051/X hold115/X vssd1 vssd1 vccd1 vccd1 _08359_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_47_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08289_ _15513_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08289_/X sky130_fd_sc_hd__or2_1
XFILLER_0_190_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6130 data_in[8] vssd1 vssd1 vccd1 vccd1 hold449/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10320_ _10470_/A _10320_/B vssd1 vssd1 vccd1 vccd1 _10320_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5440 _17034_/Q vssd1 vssd1 vccd1 vccd1 hold5440/X sky130_fd_sc_hd__dlygate4sd3_1
X_10251_ _10515_/A _10251_/B vssd1 vssd1 vccd1 vccd1 _10251_/X sky130_fd_sc_hd__or2_1
Xhold5451 _10690_/X vssd1 vssd1 vccd1 vccd1 _16720_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5462 _17141_/Q vssd1 vssd1 vccd1 vccd1 hold5462/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5473 _13372_/X vssd1 vssd1 vccd1 vccd1 _17577_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5484 _17002_/Q vssd1 vssd1 vccd1 vccd1 hold5484/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5495 _13597_/X vssd1 vssd1 vccd1 vccd1 _17652_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4750 _12070_/X vssd1 vssd1 vccd1 vccd1 _17180_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10182_ _10530_/A _10182_/B vssd1 vssd1 vccd1 vccd1 _10182_/X sky130_fd_sc_hd__or2_1
Xhold4761 _13001_/X vssd1 vssd1 vccd1 vccd1 _13002_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4772 _13546_/X vssd1 vssd1 vccd1 vccd1 _17635_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4783 _16984_/Q vssd1 vssd1 vccd1 vccd1 hold4783/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4794 _12007_/X vssd1 vssd1 vccd1 vccd1 _17159_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_218_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14990_ _15205_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14990_/X sky130_fd_sc_hd__or2_1
XFILLER_0_121_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout250 _13800_/A vssd1 vssd1 vccd1 vccd1 _13716_/A sky130_fd_sc_hd__buf_4
Xfanout261 _11622_/A vssd1 vssd1 vccd1 vccd1 _12093_/A sky130_fd_sc_hd__buf_4
Xfanout272 _13581_/A vssd1 vssd1 vccd1 vccd1 _13773_/A sky130_fd_sc_hd__buf_4
Xfanout283 _12273_/A vssd1 vssd1 vccd1 vccd1 _13749_/A sky130_fd_sc_hd__buf_4
X_13941_ _13941_/A _13941_/B vssd1 vssd1 vccd1 vccd1 _17778_/D sky130_fd_sc_hd__and2_1
XFILLER_0_233_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout294 fanout299/X vssd1 vssd1 vccd1 vccd1 _11697_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_195_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_23_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_23_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_16660_ _18220_/CLK _16660_/D vssd1 vssd1 vccd1 vccd1 _16660_/Q sky130_fd_sc_hd__dfxtp_1
X_13872_ hold4367/X _13773_/A _13871_/X vssd1 vssd1 vccd1 vccd1 _13872_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_236_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15611_ _18430_/CLK _15611_/D vssd1 vssd1 vccd1 vccd1 _15611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12823_ hold2571/X _17452_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _12823_/X sky130_fd_sc_hd__mux2_1
X_16591_ _18149_/CLK _16591_/D vssd1 vssd1 vccd1 vccd1 _16591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18330_ _18394_/CLK _18330_/D vssd1 vssd1 vccd1 vccd1 _18330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15542_ hold2802/X _15547_/B _15541_/Y _12873_/A vssd1 vssd1 vccd1 vccd1 _15542_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_201_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12754_ _16249_/Q hold3226/X _12766_/S vssd1 vssd1 vccd1 vccd1 _12754_/X sky130_fd_sc_hd__mux2_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18261_ _18389_/CLK hold997/X vssd1 vssd1 vccd1 vccd1 hold996/A sky130_fd_sc_hd__dfxtp_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ hold3035/X hold4093/X _12335_/C vssd1 vssd1 vccd1 vccd1 _11706_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_84_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15473_ _15473_/A _15473_/B vssd1 vssd1 vccd1 vccd1 _18423_/D sky130_fd_sc_hd__and2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ hold1738/X hold3362/X _12844_/S vssd1 vssd1 vccd1 vccd1 _12685_/X sky130_fd_sc_hd__mux2_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_144_wb_clk_i clkbuf_6_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18374_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_1312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17212_ _17244_/CLK _17212_/D vssd1 vssd1 vccd1 vccd1 _17212_/Q sky130_fd_sc_hd__dfxtp_1
X_14424_ hold1843/X _14433_/B _14423_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _14424_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11636_ _17884_/Q _17036_/Q _11732_/C vssd1 vssd1 vccd1 vccd1 _11637_/B sky130_fd_sc_hd__mux2_1
X_18192_ _18192_/CLK _18192_/D vssd1 vssd1 vccd1 vccd1 _18192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17143_ _17281_/CLK _17143_/D vssd1 vssd1 vccd1 vccd1 _17143_/Q sky130_fd_sc_hd__dfxtp_1
X_14355_ hold933/A hold1281/X _14381_/S vssd1 vssd1 vccd1 vccd1 _14355_/X sky130_fd_sc_hd__mux2_1
X_11567_ hold1849/X hold4989/X _11765_/C vssd1 vssd1 vccd1 vccd1 _11568_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10518_ _10536_/A _10518_/B vssd1 vssd1 vccd1 vccd1 _10518_/X sky130_fd_sc_hd__or2_1
X_13306_ _17589_/Q _17123_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13306_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_150_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold709 hold709/A vssd1 vssd1 vccd1 vccd1 hold709/X sky130_fd_sc_hd__dlygate4sd3_1
X_17074_ _17859_/CLK _17074_/D vssd1 vssd1 vccd1 vccd1 _17074_/Q sky130_fd_sc_hd__dfxtp_1
X_14286_ hold445/X _14502_/B vssd1 vssd1 vccd1 vccd1 _14286_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_40_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11498_ hold1233/X hold5347/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11499_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16025_ _16026_/CLK _16025_/D vssd1 vssd1 vccd1 vccd1 hold845/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13237_ _13236_/X hold3503/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13237_/X sky130_fd_sc_hd__mux2_1
X_10449_ _10551_/A _10449_/B vssd1 vssd1 vccd1 vccd1 _10449_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13168_ _13161_/X _13167_/X _13296_/B1 vssd1 vssd1 vccd1 vccd1 _17539_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_6_62_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_62_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_12119_ hold1817/X hold5062/X _13481_/S vssd1 vssd1 vccd1 vccd1 _12120_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17976_ _17976_/CLK _17976_/D vssd1 vssd1 vccd1 vccd1 _17976_/Q sky130_fd_sc_hd__dfxtp_1
X_13099_ _13098_/X hold6003/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13099_/X sky130_fd_sc_hd__mux2_1
Xhold1409 _17827_/Q vssd1 vssd1 vccd1 vccd1 hold1409/X sky130_fd_sc_hd__dlygate4sd3_1
X_16927_ _17799_/CLK _16927_/D vssd1 vssd1 vccd1 vccd1 _16927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16858_ _18066_/CLK _16858_/D vssd1 vssd1 vccd1 vccd1 _16858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15809_ _17624_/CLK _15809_/D vssd1 vssd1 vccd1 vccd1 _15809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16789_ _18024_/CLK _16789_/D vssd1 vssd1 vccd1 vccd1 _16789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ hold1696/X _09325_/B _09329_/X _12597_/A vssd1 vssd1 vccd1 vccd1 _09330_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09261_ _15537_/A hold1237/X hold271/X vssd1 vssd1 vccd1 vccd1 _09262_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_47_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18459_ _18462_/CLK _18459_/D vssd1 vssd1 vccd1 vccd1 _18459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08212_ hold1425/X _08213_/B _08211_/Y _08389_/A vssd1 vssd1 vccd1 vccd1 _08212_/X
+ sky130_fd_sc_hd__o211a_1
X_09192_ _15521_/A _09206_/B vssd1 vssd1 vccd1 vccd1 _09192_/X sky130_fd_sc_hd__or2_1
XFILLER_0_172_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08143_ _08143_/A hold109/X vssd1 vssd1 vccd1 vccd1 hold110/A sky130_fd_sc_hd__and2_1
XFILLER_0_71_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08074_ _15533_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08074_/X sky130_fd_sc_hd__or2_1
Xhold4002 _10396_/X vssd1 vssd1 vccd1 vccd1 _16622_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4013 _16586_/Q vssd1 vssd1 vccd1 vccd1 hold4013/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4024 _16621_/Q vssd1 vssd1 vccd1 vccd1 hold4024/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4035 _09649_/X vssd1 vssd1 vccd1 vccd1 _16373_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3301 _16633_/Q vssd1 vssd1 vccd1 vccd1 hold3301/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4046 _17184_/Q vssd1 vssd1 vccd1 vccd1 hold4046/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4057 _10720_/X vssd1 vssd1 vccd1 vccd1 _16730_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3312 _17482_/Q vssd1 vssd1 vccd1 vccd1 hold3312/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3323 _10159_/X vssd1 vssd1 vccd1 vccd1 _16543_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4068 _16774_/Q vssd1 vssd1 vccd1 vccd1 hold4068/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3334 _17481_/Q vssd1 vssd1 vccd1 vccd1 hold3334/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4079 _16710_/Q vssd1 vssd1 vccd1 vccd1 hold4079/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3345 _16629_/Q vssd1 vssd1 vccd1 vccd1 hold3345/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2600 _07921_/X vssd1 vssd1 vccd1 vccd1 _15604_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2611 _16166_/Q vssd1 vssd1 vccd1 vccd1 hold2611/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3356 _17393_/Q vssd1 vssd1 vccd1 vccd1 hold3356/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__clkbuf_2
XTAP_5529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3367 _12842_/X vssd1 vssd1 vccd1 vccd1 _12843_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2622 _15703_/Q vssd1 vssd1 vccd1 vccd1 hold2622/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08976_ _15254_/A _08976_/B vssd1 vssd1 vccd1 vccd1 _16105_/D sky130_fd_sc_hd__and2_1
Xhold3378 _12827_/X vssd1 vssd1 vccd1 vccd1 _12828_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2633 _16198_/Q vssd1 vssd1 vccd1 vccd1 hold2633/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2644 _14675_/X vssd1 vssd1 vccd1 vccd1 _18130_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3389 _17370_/Q vssd1 vssd1 vccd1 vccd1 hold3389/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1910 _09149_/X vssd1 vssd1 vccd1 vccd1 _16187_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__buf_2
Xhold2655 _15675_/Q vssd1 vssd1 vccd1 vccd1 hold2655/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2666 _18034_/Q vssd1 vssd1 vccd1 vccd1 hold2666/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1921 _16225_/Q vssd1 vssd1 vccd1 vccd1 hold1921/X sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ hold1945/X _07924_/B _07926_/X _12199_/C1 vssd1 vssd1 vccd1 vccd1 _07927_/X
+ sky130_fd_sc_hd__o211a_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2677 _18156_/Q vssd1 vssd1 vccd1 vccd1 hold2677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1932 _09099_/X vssd1 vssd1 vccd1 vccd1 _16164_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2688 _08237_/X vssd1 vssd1 vccd1 vccd1 _15753_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1943 _17755_/Q vssd1 vssd1 vccd1 vccd1 hold1943/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2699 _18292_/Q vssd1 vssd1 vccd1 vccd1 hold2699/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1954 _08022_/X vssd1 vssd1 vccd1 vccd1 _15652_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1965 _14436_/X vssd1 vssd1 vccd1 vccd1 _18016_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07858_ hold1762/X _07869_/B _07857_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _07858_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1976 _18095_/Q vssd1 vssd1 vccd1 vccd1 hold1976/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1987 _14709_/X vssd1 vssd1 vccd1 vccd1 _18146_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1998 _18185_/Q vssd1 vssd1 vccd1 vccd1 hold1998/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07789_ _07789_/A vssd1 vssd1 vccd1 vccd1 _09342_/A sky130_fd_sc_hd__inv_2
XFILLER_0_151_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09528_ _09948_/A _09528_/B vssd1 vssd1 vccd1 vccd1 _09528_/X sky130_fd_sc_hd__or2_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _09463_/C _09463_/D _09458_/Y vssd1 vssd1 vccd1 vccd1 _16313_/D sky130_fd_sc_hd__o21a_1
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_213_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12470_ _17328_/Q _12506_/B vssd1 vssd1 vccd1 vccd1 _12470_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11421_ _11553_/A _11421_/B vssd1 vssd1 vccd1 vccd1 _11421_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14140_ _14604_/A _14140_/B vssd1 vssd1 vccd1 vccd1 _14140_/X sky130_fd_sc_hd__or2_1
X_11352_ _11649_/A _11352_/B vssd1 vssd1 vccd1 vccd1 _11352_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10303_ hold3339/X _10649_/B _10302_/X _14691_/C1 vssd1 vssd1 vccd1 vccd1 _10303_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14071_ hold1511/X _14107_/A2 _14070_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _14071_/X
+ sky130_fd_sc_hd__o211a_1
X_11283_ _11661_/A _11283_/B vssd1 vssd1 vccd1 vccd1 _11283_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13022_ _09494_/A hold904/A _11203_/A vssd1 vssd1 vccd1 vccd1 hold905/A sky130_fd_sc_hd__a21oi_1
Xhold5270 _11518_/X vssd1 vssd1 vccd1 vccd1 _16996_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10234_ hold5092/X _10616_/B _10233_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _10234_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5281 _17700_/Q vssd1 vssd1 vccd1 vccd1 hold5281/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5292 _11680_/X vssd1 vssd1 vccd1 vccd1 _17050_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_1250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4580 _10546_/X vssd1 vssd1 vccd1 vccd1 _16672_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17830_ _18060_/CLK _17830_/D vssd1 vssd1 vccd1 vccd1 _17830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4591 _16365_/Q vssd1 vssd1 vccd1 vccd1 hold4591/X sky130_fd_sc_hd__dlygate4sd3_1
X_10165_ hold4600/X _10646_/B _10164_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10165_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3890 _16671_/Q vssd1 vssd1 vccd1 vccd1 hold3890/X sky130_fd_sc_hd__dlygate4sd3_1
X_17761_ _17838_/CLK _17761_/D vssd1 vssd1 vccd1 vccd1 _17761_/Q sky130_fd_sc_hd__dfxtp_1
X_14973_ hold1609/X _15004_/B _14972_/X _15482_/A vssd1 vssd1 vccd1 vccd1 _14973_/X
+ sky130_fd_sc_hd__o211a_1
X_10096_ hold5146/X _11186_/B _10095_/X _15160_/C1 vssd1 vssd1 vccd1 vccd1 _10096_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16712_ _18043_/CLK _16712_/D vssd1 vssd1 vccd1 vccd1 _16712_/Q sky130_fd_sc_hd__dfxtp_1
X_13924_ _14604_/A hold1505/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13925_/B sky130_fd_sc_hd__mux2_1
X_17692_ _17724_/CLK _17692_/D vssd1 vssd1 vccd1 vccd1 _17692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_396_wb_clk_i clkbuf_6_36_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17887_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_236_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16643_ _18224_/CLK _16643_/D vssd1 vssd1 vccd1 vccd1 _16643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13855_ _13888_/A _13855_/B vssd1 vssd1 vccd1 vccd1 _13855_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_325_wb_clk_i clkbuf_6_46_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17779_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ hold3210/X _12805_/X _12839_/S vssd1 vssd1 vccd1 vccd1 _12806_/X sky130_fd_sc_hd__mux2_1
X_16574_ _18210_/CLK _16574_/D vssd1 vssd1 vccd1 vccd1 _16574_/Q sky130_fd_sc_hd__dfxtp_1
X_10998_ _11121_/A _10998_/B vssd1 vssd1 vccd1 vccd1 _10998_/X sky130_fd_sc_hd__or2_1
XFILLER_0_128_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13786_ hold5464/X _13880_/B _13785_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13786_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18313_ _18347_/CLK _18313_/D vssd1 vssd1 vccd1 vccd1 hold654/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15525_ _15525_/A _15549_/B vssd1 vssd1 vccd1 vccd1 _15525_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ hold3161/X _12736_/X _12749_/S vssd1 vssd1 vccd1 vccd1 _12737_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _18372_/CLK _18244_/D vssd1 vssd1 vccd1 vccd1 _18244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15456_ hold854/X _09365_/B _09392_/B hold588/X vssd1 vssd1 vccd1 vccd1 _15456_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12668_ hold3145/X _12667_/X _12851_/S vssd1 vssd1 vccd1 vccd1 _12669_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_170_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14407_ _14980_/A _14443_/B vssd1 vssd1 vccd1 vccd1 _14407_/X sky130_fd_sc_hd__or2_1
XFILLER_0_115_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18175_ _18205_/CLK _18175_/D vssd1 vssd1 vccd1 vccd1 _18175_/Q sky130_fd_sc_hd__dfxtp_1
X_11619_ _12093_/A _11619_/B vssd1 vssd1 vccd1 vccd1 _11619_/X sky130_fd_sc_hd__or2_1
X_15387_ hold459/X _09357_/A _09386_/D _15896_/Q _15386_/X vssd1 vssd1 vccd1 vccd1
+ _15392_/B sky130_fd_sc_hd__a221o_2
XFILLER_0_163_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12599_ hold3294/X _12598_/X _12923_/S vssd1 vssd1 vccd1 vccd1 _12600_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_80_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17126_ _17190_/CLK _17126_/D vssd1 vssd1 vccd1 vccd1 _17126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14338_ _14732_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14338_/X sky130_fd_sc_hd__or2_1
Xhold506 hold506/A vssd1 vssd1 vccd1 vccd1 hold506/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold517 hold517/A vssd1 vssd1 vccd1 vccd1 hold517/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold528 hold528/A vssd1 vssd1 vccd1 vccd1 hold528/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 hold539/A vssd1 vssd1 vccd1 vccd1 hold539/X sky130_fd_sc_hd__dlygate4sd3_1
X_17057_ _17843_/CLK _17057_/D vssd1 vssd1 vccd1 vccd1 _17057_/Q sky130_fd_sc_hd__dfxtp_1
X_14269_ hold2347/X _14268_/B _14268_/Y _15028_/A vssd1 vssd1 vccd1 vccd1 _14269_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16008_ _18416_/CLK _16008_/D vssd1 vssd1 vccd1 vccd1 hold477/A sky130_fd_sc_hd__dfxtp_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_wb_clk_i clkbuf_6_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17877_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ hold169/X hold379/X _08860_/S vssd1 vssd1 vccd1 vccd1 hold380/A sky130_fd_sc_hd__mux2_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 _07854_/X vssd1 vssd1 vccd1 vccd1 _15572_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ hold180/X hold699/X _08779_/S vssd1 vssd1 vccd1 vccd1 hold700/A sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 _15712_/Q vssd1 vssd1 vccd1 vccd1 hold1217/X sky130_fd_sc_hd__dlygate4sd3_1
X_17959_ _17964_/CLK _17959_/D vssd1 vssd1 vccd1 vccd1 _17959_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 _08436_/X vssd1 vssd1 vccd1 vccd1 _15848_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1239 _17792_/Q vssd1 vssd1 vccd1 vccd1 hold1239/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_240_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08692_ _15414_/A hold609/X vssd1 vssd1 vccd1 vccd1 _15967_/D sky130_fd_sc_hd__and2_1
XFILLER_0_212_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09313_ _09313_/A _09315_/B vssd1 vssd1 vccd1 vccd1 _09313_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09244_ _12786_/A hold918/X vssd1 vssd1 vccd1 vccd1 _16233_/D sky130_fd_sc_hd__and2_1
XFILLER_0_75_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09175_ hold1334/X _09177_/A2 _09174_/X _12924_/A vssd1 vssd1 vccd1 vccd1 _09175_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08126_ _15531_/A _15702_/Q hold108/X vssd1 vssd1 vccd1 vccd1 _08126_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08057_ hold2877/X _08097_/A2 _08056_/X _08363_/A vssd1 vssd1 vccd1 vccd1 _08057_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3120 _17467_/Q vssd1 vssd1 vccd1 vccd1 hold3120/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3131 _17372_/Q vssd1 vssd1 vccd1 vccd1 hold3131/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3142 _12905_/X vssd1 vssd1 vccd1 vccd1 _12906_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3153 _12881_/X vssd1 vssd1 vccd1 vccd1 _12882_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3164 _14581_/X vssd1 vssd1 vccd1 vccd1 _18084_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2430 _14325_/X vssd1 vssd1 vccd1 vccd1 _17962_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3175 _17426_/Q vssd1 vssd1 vccd1 vccd1 hold3175/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2441 _18086_/Q vssd1 vssd1 vccd1 vccd1 hold2441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3186 _18377_/Q vssd1 vssd1 vccd1 vccd1 hold3186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3197 _16343_/Q vssd1 vssd1 vccd1 vccd1 _13214_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2452 _08434_/X vssd1 vssd1 vccd1 vccd1 _15847_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08959_ hold77/X _16097_/Q _08991_/S vssd1 vssd1 vccd1 vccd1 hold250/A sky130_fd_sc_hd__mux2_1
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2463 _09193_/X vssd1 vssd1 vccd1 vccd1 _16208_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_1393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2474 _15605_/Q vssd1 vssd1 vccd1 vccd1 hold2474/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2485 _18163_/Q vssd1 vssd1 vccd1 vccd1 hold2485/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1740 _15575_/Q vssd1 vssd1 vccd1 vccd1 hold1740/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1751 _14839_/X vssd1 vssd1 vccd1 vccd1 _18209_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2496 _09324_/X vssd1 vssd1 vccd1 vccd1 _16272_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _13314_/A _11970_/B vssd1 vssd1 vccd1 vccd1 _11970_/X sky130_fd_sc_hd__or2_1
Xhold1762 _15574_/Q vssd1 vssd1 vccd1 vccd1 hold1762/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1773 _15777_/Q vssd1 vssd1 vccd1 vccd1 hold1773/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1784 _13977_/X vssd1 vssd1 vccd1 vccd1 _17795_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1795 _15763_/Q vssd1 vssd1 vccd1 vccd1 hold1795/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10921_ hold5154/X _11789_/B _10920_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _10921_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_233_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10852_ hold5327/X _11732_/B _10851_/X _13895_/A vssd1 vssd1 vccd1 vccd1 _10852_/X
+ sky130_fd_sc_hd__o211a_1
X_13640_ hold1215/X _17667_/Q _13862_/C vssd1 vssd1 vccd1 vccd1 _13641_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ hold5647/X _11071_/A2 _10782_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _10783_/X
+ sky130_fd_sc_hd__o211a_1
X_13571_ hold1773/X _17644_/Q _13841_/C vssd1 vssd1 vccd1 vccd1 _13572_/B sky130_fd_sc_hd__mux2_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15310_ hold763/X _09367_/A _15446_/B1 hold880/X vssd1 vssd1 vccd1 vccd1 _15310_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12522_ _12984_/A _12522_/B vssd1 vssd1 vccd1 vccd1 _17350_/D sky130_fd_sc_hd__and2_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _18408_/CLK _16290_/D vssd1 vssd1 vccd1 vccd1 _16290_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15241_ _09404_/B _15477_/A2 _15487_/B1 hold466/X _15240_/X vssd1 vssd1 vccd1 vccd1
+ _15242_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_240_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12453_ hold684/X _12509_/A2 _12501_/A3 _12452_/X _12426_/A vssd1 vssd1 vccd1 vccd1
+ hold159/A sky130_fd_sc_hd__o311a_1
XFILLER_0_23_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11404_ hold5347/X _12329_/B _11403_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11404_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12384_ _12438_/A hold809/X vssd1 vssd1 vccd1 vccd1 _17285_/D sky130_fd_sc_hd__and2_1
X_15172_ hold6052/X _15167_/B hold842/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 hold843/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_1348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_240_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14123_ hold3068/X _14142_/B _14122_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _14123_/X
+ sky130_fd_sc_hd__o211a_1
X_11335_ hold5659/X _12299_/B _11334_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _11335_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_239_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11266_ hold4018/X _12317_/B _11265_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11266_/X
+ sky130_fd_sc_hd__o211a_1
X_14054_ _14735_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14054_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_197_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10217_ hold1889/X hold3840/X _10601_/C vssd1 vssd1 vccd1 vccd1 _10218_/B sky130_fd_sc_hd__mux2_1
X_13005_ hold927/X _13017_/B vssd1 vssd1 vccd1 vccd1 _13005_/X sky130_fd_sc_hd__or2_1
XTAP_6550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11197_ _12331_/A _11197_/B vssd1 vssd1 vccd1 vccd1 _11197_/Y sky130_fd_sc_hd__nor2_1
XTAP_6561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17813_ _17877_/CLK _17813_/D vssd1 vssd1 vccd1 vccd1 _17813_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10148_ hold2300/X hold4225/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10149_/B sky130_fd_sc_hd__mux2_1
XTAP_6594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17744_ _17744_/CLK _17744_/D vssd1 vssd1 vccd1 vccd1 _17744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10079_ _18075_/Q _16517_/Q _10571_/C vssd1 vssd1 vccd1 vccd1 _10080_/B sky130_fd_sc_hd__mux2_1
X_14956_ _15225_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14956_/X sky130_fd_sc_hd__or2_1
XFILLER_0_238_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13907_ _13929_/A _13907_/B vssd1 vssd1 vccd1 vccd1 _17761_/D sky130_fd_sc_hd__and2_1
XFILLER_0_203_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17675_ _17707_/CLK _17675_/D vssd1 vssd1 vccd1 vccd1 _17675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14887_ hold1801/X hold332/X _14886_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _14887_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16626_ _18170_/CLK _16626_/D vssd1 vssd1 vccd1 vccd1 _16626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13838_ _17733_/Q _13856_/B _13871_/C vssd1 vssd1 vccd1 vccd1 _13838_/X sky130_fd_sc_hd__and3_1
XFILLER_0_43_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16557_ _18087_/CLK _16557_/D vssd1 vssd1 vccd1 vccd1 _16557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13769_ hold1680/X hold4048/X _13865_/C vssd1 vssd1 vccd1 vccd1 _13770_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15508_ hold445/X hold363/X vssd1 vssd1 vccd1 vccd1 _15549_/B sky130_fd_sc_hd__or2_2
XFILLER_0_116_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16488_ _18373_/CLK _16488_/D vssd1 vssd1 vccd1 vccd1 _16488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18227_ _18227_/CLK _18227_/D vssd1 vssd1 vccd1 vccd1 _18227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15439_ hold718/X _09386_/A _15437_/X vssd1 vssd1 vccd1 vccd1 _15442_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18158_ _18226_/CLK _18158_/D vssd1 vssd1 vccd1 vccd1 _18158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold303 hold303/A vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold314 input23/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dlygate4sd3_1
X_17109_ _17269_/CLK _17109_/D vssd1 vssd1 vccd1 vccd1 _17109_/Q sky130_fd_sc_hd__dfxtp_1
Xhold325 hold325/A vssd1 vssd1 vccd1 vccd1 hold325/X sky130_fd_sc_hd__dlygate4sd3_1
X_18089_ _18177_/CLK _18089_/D vssd1 vssd1 vccd1 vccd1 _18089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold336 input57/X vssd1 vssd1 vccd1 vccd1 hold336/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 hold347/A vssd1 vssd1 vccd1 vccd1 hold347/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold358 hold358/A vssd1 vssd1 vccd1 vccd1 hold358/X sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ hold4610/X _10025_/B _09930_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09931_/X
+ sky130_fd_sc_hd__o211a_1
Xhold369 hold369/A vssd1 vssd1 vccd1 vccd1 hold369/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout805 _15066_/A vssd1 vssd1 vccd1 vccd1 _15064_/A sky130_fd_sc_hd__buf_4
Xfanout816 fanout843/X vssd1 vssd1 vccd1 vccd1 fanout816/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout827 _14863_/C1 vssd1 vssd1 vccd1 vccd1 _14887_/C1 sky130_fd_sc_hd__buf_4
X_09862_ hold4158/X _10052_/B _09861_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _16444_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout838 _14691_/C1 vssd1 vssd1 vccd1 vccd1 _14889_/C1 sky130_fd_sc_hd__buf_4
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout849 _17754_/Q vssd1 vssd1 vccd1 vccd1 _12331_/A sky130_fd_sc_hd__buf_8
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08813_ _15364_/A _08813_/B vssd1 vssd1 vccd1 vccd1 _16025_/D sky130_fd_sc_hd__and2_1
Xhold1003 _15198_/X vssd1 vssd1 vccd1 vccd1 _18381_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ hold4640/X _10031_/B _09792_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09793_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1014 _17995_/Q vssd1 vssd1 vccd1 vccd1 hold1014/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_247_wb_clk_i clkbuf_6_59_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18220_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1025 _15566_/Q vssd1 vssd1 vccd1 vccd1 hold1025/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1036 _14053_/X vssd1 vssd1 vccd1 vccd1 _17832_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1047 _17925_/Q vssd1 vssd1 vccd1 vccd1 hold1047/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ _12410_/A _08744_/B vssd1 vssd1 vccd1 vccd1 _15992_/D sky130_fd_sc_hd__and2_1
Xhold1058 _18152_/Q vssd1 vssd1 vccd1 vccd1 hold1058/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1069 _16239_/Q vssd1 vssd1 vccd1 vccd1 hold1069/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ hold147/X hold732/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08676_/B sky130_fd_sc_hd__mux2_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09227_ hold1921/X _09218_/B _09226_/X _12843_/A vssd1 vssd1 vccd1 vccd1 _09227_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09158_ _15541_/A _09164_/B vssd1 vssd1 vccd1 vccd1 _09158_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08109_ _08137_/A _08109_/B vssd1 vssd1 vccd1 vccd1 _15693_/D sky130_fd_sc_hd__and2_1
XFILLER_0_47_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09089_ hold2769/X _09102_/B _09088_/X _14358_/A vssd1 vssd1 vccd1 vccd1 _09089_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11120_ hold2353/X hold5074/X _11216_/C vssd1 vssd1 vccd1 vccd1 _11121_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold870 hold870/A vssd1 vssd1 vccd1 vccd1 hold870/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 hold881/A vssd1 vssd1 vccd1 vccd1 hold881/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 input3/X vssd1 vssd1 vccd1 vccd1 hold892/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11051_ hold1517/X _16841_/Q _11153_/C vssd1 vssd1 vccd1 vccd1 _11052_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_219_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10002_ _13118_/A _09912_/A _10001_/X vssd1 vssd1 vccd1 vccd1 _10002_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2260 _15146_/X vssd1 vssd1 vccd1 vccd1 _18356_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ _14988_/A _14830_/B vssd1 vssd1 vccd1 vccd1 _14810_/X sky130_fd_sc_hd__or2_1
XTAP_5178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2271 _12512_/X vssd1 vssd1 vccd1 vccd1 hold2271/X sky130_fd_sc_hd__buf_1
Xhold2282 _18089_/Q vssd1 vssd1 vccd1 vccd1 hold2282/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15790_ _17722_/CLK _15790_/D vssd1 vssd1 vccd1 vccd1 _15790_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2293 _15682_/Q vssd1 vssd1 vccd1 vccd1 hold2293/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1570 _17873_/Q vssd1 vssd1 vccd1 vccd1 hold1570/X sky130_fd_sc_hd__dlygate4sd3_1
X_14741_ hold2135/X _14772_/B _14740_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14741_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1581 _14170_/X vssd1 vssd1 vccd1 vccd1 hold1581/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1592 _17965_/Q vssd1 vssd1 vccd1 vccd1 hold1592/X sky130_fd_sc_hd__dlygate4sd3_1
X_11953_ hold5575/X _12335_/B _11952_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11953_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10904_ hold1014/X _16792_/Q _11789_/C vssd1 vssd1 vccd1 vccd1 _10905_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17460_ _17462_/CLK _17460_/D vssd1 vssd1 vccd1 vccd1 _17460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14672_ _14726_/A _14672_/B vssd1 vssd1 vccd1 vccd1 _14672_/X sky130_fd_sc_hd__or2_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11884_ hold5773/X _12362_/B _11883_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _11884_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16411_ _18324_/CLK _16411_/D vssd1 vssd1 vccd1 vccd1 _16411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13623_ _13719_/A _13623_/B vssd1 vssd1 vccd1 vccd1 _13623_/X sky130_fd_sc_hd__or2_1
XFILLER_0_95_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17391_ _18443_/CLK _17391_/D vssd1 vssd1 vccd1 vccd1 _17391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10835_ _17972_/Q _16769_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _10836_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16342_ _18327_/CLK _16342_/D vssd1 vssd1 vccd1 vccd1 _16342_/Q sky130_fd_sc_hd__dfxtp_1
X_13554_ _13752_/A _13554_/B vssd1 vssd1 vccd1 vccd1 _13554_/X sky130_fd_sc_hd__or2_1
X_10766_ hold537/X _16746_/Q _11723_/C vssd1 vssd1 vccd1 vccd1 _10767_/B sky130_fd_sc_hd__mux2_1
X_12505_ hold56/X _08597_/Y _08868_/X _12504_/X _09003_/A vssd1 vssd1 vccd1 vccd1
+ hold57/A sky130_fd_sc_hd__o311a_1
XFILLER_0_165_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16273_ _17374_/CLK hold962/X vssd1 vssd1 vccd1 vccd1 hold961/A sky130_fd_sc_hd__dfxtp_1
X_10697_ hold3104/X hold4341/X _11204_/C vssd1 vssd1 vccd1 vccd1 _10698_/B sky130_fd_sc_hd__mux2_1
X_13485_ _13581_/A _13485_/B vssd1 vssd1 vccd1 vccd1 _13485_/X sky130_fd_sc_hd__or2_1
X_18012_ _18461_/CLK _18012_/D vssd1 vssd1 vccd1 vccd1 _18012_/Q sky130_fd_sc_hd__dfxtp_1
X_15224_ hold6063/X _15219_/B hold485/X _15024_/A vssd1 vssd1 vccd1 vccd1 hold486/A
+ sky130_fd_sc_hd__o211a_1
X_12436_ _15374_/A hold119/X vssd1 vssd1 vccd1 vccd1 _17311_/D sky130_fd_sc_hd__and2_1
XFILLER_0_120_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15155_ _15209_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15155_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12367_ _13888_/A _12367_/B vssd1 vssd1 vccd1 vccd1 _12367_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_23_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14106_ _14732_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14106_/X sky130_fd_sc_hd__or2_1
XFILLER_0_239_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_238_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ hold1093/X hold4295/X _12173_/S vssd1 vssd1 vccd1 vccd1 _11319_/B sky130_fd_sc_hd__mux2_1
X_15086_ hold1031/X hold340/X _15085_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _15086_/X
+ sky130_fd_sc_hd__o211a_1
X_12298_ _13819_/A _12298_/B vssd1 vssd1 vccd1 vccd1 _12298_/Y sky130_fd_sc_hd__nor2_1
X_14037_ hold2526/X _14040_/B _14036_/Y _13905_/A vssd1 vssd1 vccd1 vccd1 _14037_/X
+ sky130_fd_sc_hd__o211a_1
X_11249_ hold1943/X hold4345/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11250_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_340_wb_clk_i clkbuf_6_43_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17749_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15988_ _18308_/CLK _15988_/D vssd1 vssd1 vccd1 vccd1 _15988_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17727_ _17729_/CLK _17727_/D vssd1 vssd1 vccd1 vccd1 _17727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14939_ hold1211/X _14946_/B _14938_/X _15204_/C1 vssd1 vssd1 vccd1 vccd1 _14939_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08460_ _15085_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08460_/X sky130_fd_sc_hd__or2_1
X_17658_ _17690_/CLK _17658_/D vssd1 vssd1 vccd1 vccd1 _17658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16609_ _18218_/CLK _16609_/D vssd1 vssd1 vccd1 vccd1 _16609_/Q sky130_fd_sc_hd__dfxtp_1
X_08391_ _08391_/A _08391_/B vssd1 vssd1 vccd1 vccd1 _15827_/D sky130_fd_sc_hd__and2_1
XFILLER_0_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17589_ _17735_/CLK _17589_/D vssd1 vssd1 vccd1 vccd1 _17589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09012_ hold29/X hold327/X _09060_/S vssd1 vssd1 vccd1 vccd1 _09013_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5803 _17234_/Q vssd1 vssd1 vccd1 vccd1 hold5803/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold100 hold100/A vssd1 vssd1 vccd1 vccd1 hold100/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5814 _13324_/X vssd1 vssd1 vccd1 vccd1 _17561_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5825 _16366_/Q vssd1 vssd1 vccd1 vccd1 hold5825/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5836 _09844_/X vssd1 vssd1 vccd1 vccd1 _16438_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold111 hold506/X vssd1 vssd1 vccd1 vccd1 hold507/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5847 hold6009/X vssd1 vssd1 vccd1 vccd1 _13241_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 input17/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__buf_1
Xhold5858 output88/X vssd1 vssd1 vccd1 vccd1 data_out[24] sky130_fd_sc_hd__buf_12
Xhold133 hold615/X vssd1 vssd1 vccd1 vccd1 hold616/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold144 hold144/A vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5869 hold6017/X vssd1 vssd1 vccd1 vccd1 _13145_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 hold155/A vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold166 hold166/A vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 hold177/A vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 hold188/A vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_428_wb_clk_i clkbuf_6_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _15856_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09914_ hold2213/X hold5823/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09915_/B sky130_fd_sc_hd__mux2_1
Xfanout602 _12513_/X vssd1 vssd1 vccd1 vccd1 _12871_/S sky130_fd_sc_hd__buf_8
XFILLER_0_10_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold199 hold288/X vssd1 vssd1 vccd1 vccd1 hold289/A sky130_fd_sc_hd__buf_6
Xfanout613 _09360_/Y vssd1 vssd1 vccd1 vccd1 _09362_/C sky130_fd_sc_hd__buf_6
Xfanout624 _15484_/A2 vssd1 vssd1 vccd1 vccd1 _09386_/A sky130_fd_sc_hd__buf_6
XFILLER_0_42_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout635 _12798_/A vssd1 vssd1 vccd1 vccd1 _12777_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_186_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout646 _12199_/C1 vssd1 vssd1 vccd1 vccd1 _08363_/A sky130_fd_sc_hd__buf_4
X_09845_ hold2412/X hold3276/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09846_/B sky130_fd_sc_hd__mux2_1
Xfanout657 _12588_/A vssd1 vssd1 vccd1 vccd1 _15502_/A sky130_fd_sc_hd__buf_4
Xfanout668 _08171_/A vssd1 vssd1 vccd1 vccd1 _08163_/A sky130_fd_sc_hd__buf_4
Xfanout679 fanout689/X vssd1 vssd1 vccd1 vccd1 _15498_/A sky130_fd_sc_hd__clkbuf_4
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09776_ hold1110/X _16416_/Q _10067_/C vssd1 vssd1 vccd1 vccd1 _09777_/B sky130_fd_sc_hd__mux2_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ hold278/X hold523/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold524/A sky130_fd_sc_hd__mux2_1
XFILLER_0_198_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_240_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08658_ _12418_/A hold669/X vssd1 vssd1 vccd1 vccd1 _15951_/D sky130_fd_sc_hd__and2_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _12416_/A hold474/X vssd1 vssd1 vccd1 vccd1 _15918_/D sky130_fd_sc_hd__and2_1
XFILLER_0_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10620_ hold3200/X _10524_/A _10619_/X vssd1 vssd1 vccd1 vccd1 _10620_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10551_ _10551_/A _10551_/B vssd1 vssd1 vccd1 vccd1 _10551_/X sky130_fd_sc_hd__or2_1
XFILLER_0_146_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10482_ _10482_/A _10482_/B vssd1 vssd1 vccd1 vccd1 _10482_/X sky130_fd_sc_hd__or2_1
X_13270_ _13270_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13270_/X sky130_fd_sc_hd__or2_1
XFILLER_0_228_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12221_ hold2912/X hold4968/X _12317_/C vssd1 vssd1 vccd1 vccd1 _12222_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_241_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12152_ hold978/X _17208_/Q _13748_/S vssd1 vssd1 vccd1 vccd1 _12153_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_241_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_169_wb_clk_i clkbuf_6_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18345_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11103_ _11103_/A _11103_/B vssd1 vssd1 vccd1 vccd1 _11103_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12083_ hold3095/X _17185_/Q _13748_/S vssd1 vssd1 vccd1 vccd1 _12084_/B sky130_fd_sc_hd__mux2_1
X_16960_ _17840_/CLK _16960_/D vssd1 vssd1 vccd1 vccd1 _16960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15911_ _17309_/CLK _15911_/D vssd1 vssd1 vccd1 vccd1 _15911_/Q sky130_fd_sc_hd__dfxtp_1
X_11034_ _11670_/A _11034_/B vssd1 vssd1 vccd1 vccd1 _11034_/X sky130_fd_sc_hd__or2_1
X_16891_ _18347_/CLK _16891_/D vssd1 vssd1 vccd1 vccd1 _16891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15842_ _17739_/CLK _15842_/D vssd1 vssd1 vccd1 vccd1 _15842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2090 _17833_/Q vssd1 vssd1 vccd1 vccd1 hold2090/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_232_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _17724_/CLK _15773_/D vssd1 vssd1 vccd1 vccd1 _15773_/Q sky130_fd_sc_hd__dfxtp_1
X_12985_ hold1748/X _17506_/Q _12985_/S vssd1 vssd1 vccd1 vccd1 _12985_/X sky130_fd_sc_hd__mux2_1
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ _17512_/CLK _17512_/D vssd1 vssd1 vccd1 vccd1 _17512_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_231_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14724_ _15225_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14724_/X sky130_fd_sc_hd__or2_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ hold1317/X _17136_/Q _12227_/S vssd1 vssd1 vccd1 vccd1 _11937_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_59_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17443_ _17725_/CLK _17443_/D vssd1 vssd1 vccd1 vccd1 _17443_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14655_ hold2047/X _14666_/B _14654_/X _14895_/C1 vssd1 vssd1 vccd1 vccd1 _14655_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11867_ hold1129/X hold5705/X _13463_/S vssd1 vssd1 vccd1 vccd1 _11868_/B sky130_fd_sc_hd__mux2_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13606_ hold4943/X _13814_/B _13605_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _13606_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10818_ _11010_/A _10818_/B vssd1 vssd1 vccd1 vccd1 _10818_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17374_ _17374_/CLK _17374_/D vssd1 vssd1 vccd1 vccd1 _17374_/Q sky130_fd_sc_hd__dfxtp_1
X_14586_ _14980_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14586_/X sky130_fd_sc_hd__or2_1
XFILLER_0_144_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11798_ _17090_/Q _11798_/B _12173_/S vssd1 vssd1 vccd1 vccd1 _11798_/X sky130_fd_sc_hd__and3_1
XFILLER_0_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16325_ _18398_/CLK _16325_/D vssd1 vssd1 vccd1 vccd1 _16325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13537_ hold4683/X _13862_/B _13536_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _13537_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10749_ _11655_/A _10749_/B vssd1 vssd1 vccd1 vccd1 _10749_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16256_ _17486_/CLK _16256_/D vssd1 vssd1 vccd1 vccd1 _16256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13468_ hold5533/X _13880_/B _13467_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13468_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15207_ _15207_/A _15227_/B vssd1 vssd1 vccd1 vccd1 _15207_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12419_ hold215/X hold518/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12420_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_211_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16187_ _18448_/CLK _16187_/D vssd1 vssd1 vccd1 vccd1 _16187_/Q sky130_fd_sc_hd__dfxtp_1
X_13399_ hold4123/X _13877_/B _13398_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _13399_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4409 _13857_/Y vssd1 vssd1 vccd1 vccd1 _13858_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15138_ hold2412/X _15167_/B _15137_/X _15146_/C1 vssd1 vssd1 vccd1 vccd1 _15138_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3708 _16410_/Q vssd1 vssd1 vccd1 vccd1 hold3708/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3719 _11107_/X vssd1 vssd1 vccd1 vccd1 _16859_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15069_ hold289/X _18320_/Q _15069_/S vssd1 vssd1 vccd1 vccd1 hold290/A sky130_fd_sc_hd__mux2_1
X_07960_ _15529_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07960_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07891_ hold2203/X _07918_/B _07890_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _07891_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09630_ _09984_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09630_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09561_ _09957_/A _09561_/B vssd1 vssd1 vccd1 vccd1 _09561_/X sky130_fd_sc_hd__or2_1
XFILLER_0_210_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08512_ hold2333/X _08503_/Y _08511_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _08512_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09492_ hold935/X _12380_/B vssd1 vssd1 vccd1 vccd1 _09494_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_33_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08443_ _14443_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08443_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08374_ hold597/X hold613/X hold115/X vssd1 vssd1 vccd1 vccd1 hold614/A sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_225_1315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5600 _11353_/X vssd1 vssd1 vccd1 vccd1 _16941_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5611 _13555_/X vssd1 vssd1 vccd1 vccd1 _17638_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5622 _17072_/Q vssd1 vssd1 vccd1 vccd1 hold5622/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5633 _16948_/Q vssd1 vssd1 vccd1 vccd1 hold5633/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5644 _13462_/X vssd1 vssd1 vccd1 vccd1 _17607_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4910 _10708_/X vssd1 vssd1 vccd1 vccd1 _16726_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5655 _17021_/Q vssd1 vssd1 vccd1 vccd1 hold5655/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4921 _17280_/Q vssd1 vssd1 vccd1 vccd1 hold4921/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5666 _11401_/X vssd1 vssd1 vccd1 vccd1 _16957_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4932 _11812_/X vssd1 vssd1 vccd1 vccd1 _17094_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5677 _17053_/Q vssd1 vssd1 vccd1 vccd1 hold5677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4943 _17687_/Q vssd1 vssd1 vccd1 vccd1 hold4943/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_262_wb_clk_i clkbuf_6_56_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18194_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5688 _12013_/X vssd1 vssd1 vccd1 vccd1 _17161_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5699 _17139_/Q vssd1 vssd1 vccd1 vccd1 hold5699/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4954 _11605_/X vssd1 vssd1 vccd1 vccd1 _17025_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4965 _17509_/Q vssd1 vssd1 vccd1 vccd1 hold4965/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_217_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4976 _17147_/Q vssd1 vssd1 vccd1 vccd1 hold4976/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout410 _14232_/Y vssd1 vssd1 vccd1 vccd1 _14268_/B sky130_fd_sc_hd__buf_8
XFILLER_0_22_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4987 _17272_/Q vssd1 vssd1 vccd1 vccd1 hold4987/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout421 _14052_/B vssd1 vssd1 vccd1 vccd1 _14042_/B sky130_fd_sc_hd__buf_6
Xfanout432 _13054_/X vssd1 vssd1 vccd1 vccd1 _13309_/S sky130_fd_sc_hd__clkbuf_16
Xhold4998 _10981_/X vssd1 vssd1 vccd1 vccd1 _16817_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout443 fanout485/X vssd1 vssd1 vccd1 vccd1 _13766_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_217_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout454 _11741_/C vssd1 vssd1 vccd1 vccd1 _12323_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_214_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout465 fanout485/X vssd1 vssd1 vccd1 vccd1 _13868_/C sky130_fd_sc_hd__buf_4
Xfanout476 _11210_/C vssd1 vssd1 vccd1 vccd1 _11753_/C sky130_fd_sc_hd__clkbuf_8
X_09828_ _09978_/A _09828_/B vssd1 vssd1 vccd1 vccd1 _09828_/X sky130_fd_sc_hd__or2_1
Xfanout487 _10964_/S vssd1 vssd1 vccd1 vccd1 _11144_/C sky130_fd_sc_hd__buf_6
Xfanout498 _10985_/S vssd1 vssd1 vccd1 vccd1 _11204_/C sky130_fd_sc_hd__buf_6
Xclkbuf_6_13_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_13_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_225_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09759_ _09978_/A _09759_/B vssd1 vssd1 vccd1 vccd1 _09759_/X sky130_fd_sc_hd__or2_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12770_ hold3570/X _12769_/X _12839_/S vssd1 vssd1 vccd1 vccd1 _12770_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ hold4674/X _12210_/A _11720_/X vssd1 vssd1 vccd1 vccd1 _11721_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_230_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ hold2646/X _14433_/B _14439_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _14440_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _12219_/A _11652_/B vssd1 vssd1 vccd1 vccd1 _11652_/X sky130_fd_sc_hd__or2_1
XFILLER_0_194_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10603_ _10603_/A _10603_/B vssd1 vssd1 vccd1 vccd1 _16691_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_147_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14371_ _15539_/A hold1772/X _14381_/S vssd1 vssd1 vccd1 vccd1 _14372_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_80_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11583_ _12243_/A _11583_/B vssd1 vssd1 vccd1 vccd1 _11583_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16110_ _17339_/CLK _16110_/D vssd1 vssd1 vccd1 vccd1 hold569/A sky130_fd_sc_hd__dfxtp_1
X_13322_ hold2333/X hold4300/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13323_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10534_ hold5422/X _11213_/B _10533_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10534_/X
+ sky130_fd_sc_hd__o211a_1
X_17090_ _17906_/CLK _17090_/D vssd1 vssd1 vccd1 vccd1 _17090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16041_ _17297_/CLK _16041_/D vssd1 vssd1 vccd1 vccd1 hold153/A sky130_fd_sc_hd__dfxtp_1
X_10465_ hold3243/X _10571_/B _10464_/X _14893_/C1 vssd1 vssd1 vccd1 vccd1 _10465_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13253_ _13252_/X hold4225/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13253_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12204_ _12210_/A _12204_/B vssd1 vssd1 vccd1 vccd1 _12204_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13184_ _13177_/X _13183_/X _13296_/B1 vssd1 vssd1 vccd1 vccd1 _17541_/D sky130_fd_sc_hd__o21a_1
X_10396_ hold4001/X _10649_/B _10395_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10396_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_6_52_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_52_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_209_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12135_ _12159_/A _12135_/B vssd1 vssd1 vccd1 vccd1 _12135_/X sky130_fd_sc_hd__or2_1
X_17992_ _18024_/CLK _17992_/D vssd1 vssd1 vccd1 vccd1 _17992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16943_ _17889_/CLK _16943_/D vssd1 vssd1 vccd1 vccd1 _16943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_236_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12066_ _13314_/A _12066_/B vssd1 vssd1 vccd1 vccd1 _12066_/X sky130_fd_sc_hd__or2_1
XFILLER_0_198_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11017_ hold5366/X _11789_/B _11016_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _11017_/X
+ sky130_fd_sc_hd__o211a_1
X_16874_ _18045_/CLK _16874_/D vssd1 vssd1 vccd1 vccd1 _16874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15825_ _17672_/CLK _15825_/D vssd1 vssd1 vccd1 vccd1 _15825_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15756_ _17707_/CLK _15756_/D vssd1 vssd1 vccd1 vccd1 _15756_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12968_ hold3242/X _12967_/X _12971_/S vssd1 vssd1 vccd1 vccd1 _12969_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_66_wb_clk_i clkbuf_6_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17314_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14707_ hold2679/X _14718_/B _14706_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14707_/X
+ sky130_fd_sc_hd__o211a_1
X_11919_ _12198_/A _11919_/B vssd1 vssd1 vccd1 vccd1 _11919_/X sky130_fd_sc_hd__or2_1
XFILLER_0_185_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15687_ _17741_/CLK _15687_/D vssd1 vssd1 vccd1 vccd1 _15687_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12899_ hold3354/X _12898_/X _12923_/S vssd1 vssd1 vccd1 vccd1 _12900_/B sky130_fd_sc_hd__mux2_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _17426_/CLK _17426_/D vssd1 vssd1 vccd1 vccd1 _17426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14638_ _15193_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14638_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17357_ _17486_/CLK _17357_/D vssd1 vssd1 vccd1 vccd1 _17357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14569_ _15193_/A _14557_/Y hold2242/X _15218_/C1 vssd1 vssd1 vccd1 vccd1 _14569_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16308_ _16315_/CLK _16308_/D vssd1 vssd1 vccd1 vccd1 _16308_/Q sky130_fd_sc_hd__dfxtp_1
X_08090_ _15549_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08090_/X sky130_fd_sc_hd__or2_1
X_17288_ _17288_/CLK _17288_/D vssd1 vssd1 vccd1 vccd1 hold805/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16239_ _17427_/CLK _16239_/D vssd1 vssd1 vccd1 vccd1 _16239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4206 _15413_/X vssd1 vssd1 vccd1 vccd1 _15414_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4217 _16006_/Q vssd1 vssd1 vccd1 vccd1 _15365_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4228 _10644_/Y vssd1 vssd1 vccd1 vccd1 _10645_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4239 _17570_/Q vssd1 vssd1 vccd1 vccd1 hold4239/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3505 _17121_/Q vssd1 vssd1 vccd1 vccd1 hold3505/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3516 _10617_/Y vssd1 vssd1 vccd1 vccd1 _10618_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3527 _17576_/Q vssd1 vssd1 vccd1 vccd1 hold3527/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08992_ _09057_/A hold101/X vssd1 vssd1 vccd1 vccd1 _16113_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3538 _16905_/Q vssd1 vssd1 vccd1 vccd1 hold3538/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2804 _17982_/Q vssd1 vssd1 vccd1 vccd1 hold2804/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3549 _13879_/Y vssd1 vssd1 vccd1 vccd1 _17746_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2815 _18155_/Q vssd1 vssd1 vccd1 vccd1 hold2815/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2826 _15857_/Q vssd1 vssd1 vccd1 vccd1 hold2826/X sky130_fd_sc_hd__dlygate4sd3_1
X_07943_ hold1590/X _07991_/A2 _07942_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _07943_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2837 _14755_/X vssd1 vssd1 vccd1 vccd1 _18168_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2848 _15759_/Q vssd1 vssd1 vccd1 vccd1 hold2848/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2859 _15623_/Q vssd1 vssd1 vccd1 vccd1 hold2859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07874_ hold1325/X _07869_/B _07873_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _07874_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09613_ hold3694/X _10028_/B _09612_/X _15042_/A vssd1 vssd1 vccd1 vccd1 _09613_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09544_ hold5831/X _10022_/B _09543_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09544_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09475_ _09477_/B _09477_/C _09474_/Y vssd1 vssd1 vccd1 vccd1 _16319_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08426_ hold1791/X _08433_/B _08425_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08426_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08357_ _12738_/A _08357_/B vssd1 vssd1 vccd1 vccd1 _15810_/D sky130_fd_sc_hd__and2_1
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08288_ hold1773/X _08336_/A2 _08287_/X _13765_/C1 vssd1 vssd1 vccd1 vccd1 _08288_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6120 _15854_/Q vssd1 vssd1 vccd1 vccd1 hold6120/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6131 _16314_/Q vssd1 vssd1 vccd1 vccd1 hold6131/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_443_wb_clk_i clkbuf_6_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17222_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5430 _17201_/Q vssd1 vssd1 vccd1 vccd1 hold5430/X sky130_fd_sc_hd__dlygate4sd3_1
X_10250_ hold1029/X _16574_/Q _10628_/C vssd1 vssd1 vccd1 vccd1 _10251_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5441 _11536_/X vssd1 vssd1 vccd1 vccd1 _17002_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5452 _17642_/Q vssd1 vssd1 vccd1 vccd1 hold5452/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5463 _11857_/X vssd1 vssd1 vccd1 vccd1 _17109_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5474 _17006_/Q vssd1 vssd1 vccd1 vccd1 hold5474/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4740 _12160_/X vssd1 vssd1 vccd1 vccd1 _17210_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5485 _11440_/X vssd1 vssd1 vccd1 vccd1 _16970_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10181_ hold1734/X _16551_/Q _10625_/C vssd1 vssd1 vccd1 vccd1 _10182_/B sky130_fd_sc_hd__mux2_1
Xhold5496 _17708_/Q vssd1 vssd1 vccd1 vccd1 hold5496/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4751 _16915_/Q vssd1 vssd1 vccd1 vccd1 hold4751/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4762 _17097_/Q vssd1 vssd1 vccd1 vccd1 hold4762/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4773 _16488_/Q vssd1 vssd1 vccd1 vccd1 hold4773/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4784 _11386_/X vssd1 vssd1 vccd1 vccd1 _16952_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4795 _17254_/Q vssd1 vssd1 vccd1 vccd1 hold4795/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout240 _10634_/B vssd1 vssd1 vccd1 vccd1 _10067_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_206_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout251 _13800_/A vssd1 vssd1 vccd1 vccd1 _12198_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout262 fanout299/X vssd1 vssd1 vccd1 vccd1 _11622_/A sky130_fd_sc_hd__clkbuf_4
Xfanout273 _13581_/A vssd1 vssd1 vccd1 vccd1 _13776_/A sky130_fd_sc_hd__buf_2
X_13940_ _14960_/A hold1093/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13940_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_227_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout284 _12273_/A vssd1 vssd1 vccd1 vccd1 _13407_/A sky130_fd_sc_hd__buf_4
XFILLER_0_191_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout295 _11127_/A vssd1 vssd1 vccd1 vccd1 _11694_/A sky130_fd_sc_hd__buf_4
XFILLER_0_199_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13871_ _17744_/Q _13871_/B _13871_/C vssd1 vssd1 vccd1 vccd1 _13871_/X sky130_fd_sc_hd__and3_1
XFILLER_0_96_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15610_ _18445_/CLK _15610_/D vssd1 vssd1 vccd1 vccd1 _15610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12822_ _12822_/A _12822_/B vssd1 vssd1 vccd1 vccd1 _17450_/D sky130_fd_sc_hd__and2_1
X_16590_ _18154_/CLK _16590_/D vssd1 vssd1 vccd1 vccd1 _16590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_232_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15541_ _15541_/A _15547_/B vssd1 vssd1 vccd1 vccd1 _15541_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_96_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12753_ _12753_/A _12753_/B vssd1 vssd1 vccd1 vccd1 _17427_/D sky130_fd_sc_hd__and2_1
XFILLER_0_84_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18260_ _18346_/CLK _18260_/D vssd1 vssd1 vccd1 vccd1 _18260_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ hold5016/X _11798_/B _11703_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _11704_/X
+ sky130_fd_sc_hd__o211a_1
X_15472_ _15481_/A1 _15465_/X _15471_/X _15490_/B1 _18423_/Q vssd1 vssd1 vccd1 vccd1
+ _15472_/X sky130_fd_sc_hd__a32o_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _12843_/A _12684_/B vssd1 vssd1 vccd1 vccd1 _17404_/D sky130_fd_sc_hd__and2_1
XFILLER_0_166_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17590_/CLK _17211_/D vssd1 vssd1 vccd1 vccd1 _17211_/Q sky130_fd_sc_hd__dfxtp_1
X_14423_ _15103_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14423_/X sky130_fd_sc_hd__or2_1
X_18191_ _18191_/CLK _18191_/D vssd1 vssd1 vccd1 vccd1 _18191_/Q sky130_fd_sc_hd__dfxtp_1
X_11635_ hold5197/X _11732_/B _11634_/X _13895_/A vssd1 vssd1 vccd1 vccd1 _11635_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17142_ _17906_/CLK _17142_/D vssd1 vssd1 vccd1 vccd1 _17142_/Q sky130_fd_sc_hd__dfxtp_1
X_14354_ _14354_/A _14354_/B vssd1 vssd1 vccd1 vccd1 _17976_/D sky130_fd_sc_hd__and2_1
XFILLER_0_141_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11566_ hold5321/X _11195_/B _11565_/X _14462_/C1 vssd1 vssd1 vccd1 vccd1 _11566_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_184_wb_clk_i clkbuf_6_54_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16480_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13305_ _13305_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13305_/X sky130_fd_sc_hd__and2_1
XFILLER_0_208_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10517_ hold2940/X hold3298/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10518_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17073_ _17838_/CLK _17073_/D vssd1 vssd1 vccd1 vccd1 _17073_/Q sky130_fd_sc_hd__dfxtp_1
X_14285_ hold583/X _14268_/B _14284_/X _14376_/A vssd1 vssd1 vccd1 vccd1 hold584/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11497_ hold5655/X _12329_/B _11496_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _11497_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_113_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17520_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16024_ _17338_/CLK _16024_/D vssd1 vssd1 vccd1 vccd1 hold827/A sky130_fd_sc_hd__dfxtp_1
X_13236_ hold3517/X _13235_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13236_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_0_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10448_ hold2027/X _16640_/Q _10604_/C vssd1 vssd1 vccd1 vccd1 _10449_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13167_ _13311_/A1 _13165_/X _13166_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13167_/X
+ sky130_fd_sc_hd__o211a_1
X_10379_ hold1461/X _16617_/Q _10571_/C vssd1 vssd1 vccd1 vccd1 _10380_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_236_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12118_ hold3870/X _12308_/B _12117_/X _08167_/A vssd1 vssd1 vccd1 vccd1 _12118_/X
+ sky130_fd_sc_hd__o211a_1
X_17975_ _18039_/CLK hold419/X vssd1 vssd1 vccd1 vccd1 _17975_/Q sky130_fd_sc_hd__dfxtp_1
X_13098_ _17563_/Q _17097_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13098_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12049_ hold5607/X _12335_/B _12048_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _17173_/D
+ sky130_fd_sc_hd__o211a_1
X_16926_ _17774_/CLK _16926_/D vssd1 vssd1 vccd1 vccd1 _16926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_237_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16857_ _18060_/CLK _16857_/D vssd1 vssd1 vccd1 vccd1 _16857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15808_ _17720_/CLK _15808_/D vssd1 vssd1 vccd1 vccd1 _15808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16788_ _18023_/CLK _16788_/D vssd1 vssd1 vccd1 vccd1 _16788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15739_ _17742_/CLK _15739_/D vssd1 vssd1 vccd1 vccd1 _15739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09260_ _12753_/A _09260_/B vssd1 vssd1 vccd1 vccd1 _16241_/D sky130_fd_sc_hd__and2_1
XFILLER_0_146_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18458_ _18458_/CLK _18458_/D vssd1 vssd1 vccd1 vccd1 _18458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08211_ _15219_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08211_/Y sky130_fd_sc_hd__nand2_1
X_17409_ _17434_/CLK _17409_/D vssd1 vssd1 vccd1 vccd1 _17409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09191_ hold982/X _09214_/B _09190_/X _12837_/A vssd1 vssd1 vccd1 vccd1 hold983/A
+ sky130_fd_sc_hd__o211a_1
X_18389_ _18389_/CLK _18389_/D vssd1 vssd1 vccd1 vccd1 _18389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08142_ hold97/X _15710_/Q hold108/X vssd1 vssd1 vccd1 vccd1 hold109/A sky130_fd_sc_hd__mux2_1
XFILLER_0_43_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08073_ hold1317/X _08097_/A2 _08072_/X _12289_/C1 vssd1 vssd1 vccd1 vccd1 _08073_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4003 _17678_/Q vssd1 vssd1 vccd1 vccd1 hold4003/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4014 _10192_/X vssd1 vssd1 vccd1 vccd1 _16554_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4025 _10297_/X vssd1 vssd1 vccd1 vccd1 _16589_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4036 _17437_/Q vssd1 vssd1 vccd1 vccd1 hold4036/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3302 _10333_/X vssd1 vssd1 vccd1 vccd1 _16601_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4047 _11986_/X vssd1 vssd1 vccd1 vccd1 _17152_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4058 _17419_/Q vssd1 vssd1 vccd1 vccd1 hold4058/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3313 _12917_/X vssd1 vssd1 vccd1 vccd1 _12918_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3324 _16780_/Q vssd1 vssd1 vccd1 vccd1 hold3324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4069 _10756_/X vssd1 vssd1 vccd1 vccd1 _16742_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3335 _17471_/Q vssd1 vssd1 vccd1 vccd1 hold3335/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3346 _10321_/X vssd1 vssd1 vccd1 vccd1 _16597_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2601 _18027_/Q vssd1 vssd1 vccd1 vccd1 hold2601/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2612 _09103_/X vssd1 vssd1 vccd1 vccd1 _16166_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08975_ hold5/X hold541/X _08991_/S vssd1 vssd1 vccd1 vccd1 _08976_/B sky130_fd_sc_hd__mux2_1
Xhold3357 _17388_/Q vssd1 vssd1 vccd1 vccd1 hold3357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2623 _17930_/Q vssd1 vssd1 vccd1 vccd1 hold2623/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3368 _17458_/Q vssd1 vssd1 vccd1 vccd1 hold3368/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__clkbuf_1
Xhold3379 _17403_/Q vssd1 vssd1 vccd1 vccd1 hold3379/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2634 _09171_/X vssd1 vssd1 vccd1 vccd1 _16198_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1900 _14793_/X vssd1 vssd1 vccd1 vccd1 _18186_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2645 _15723_/Q vssd1 vssd1 vccd1 vccd1 hold2645/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07926_ _15549_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07926_/X sky130_fd_sc_hd__or2_1
Xhold2656 _08071_/X vssd1 vssd1 vccd1 vccd1 _15675_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1911 _17818_/Q vssd1 vssd1 vccd1 vccd1 hold1911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2667 _14474_/X vssd1 vssd1 vccd1 vccd1 _18034_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1922 _09227_/X vssd1 vssd1 vccd1 vccd1 _16225_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_199_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1933 _18011_/Q vssd1 vssd1 vccd1 vccd1 hold1933/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2678 _14729_/X vssd1 vssd1 vccd1 vccd1 _18156_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2689 _18125_/Q vssd1 vssd1 vccd1 vccd1 hold2689/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1944 _13894_/X vssd1 vssd1 vccd1 vccd1 _13895_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1955 _17991_/Q vssd1 vssd1 vccd1 vccd1 hold1955/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1966 _15641_/Q vssd1 vssd1 vccd1 vccd1 hold1966/X sky130_fd_sc_hd__dlygate4sd3_1
X_07857_ _14529_/A _07871_/B vssd1 vssd1 vccd1 vccd1 _07857_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1977 _14603_/X vssd1 vssd1 vccd1 vccd1 _18095_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1988 _18257_/Q vssd1 vssd1 vccd1 vccd1 hold1988/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1999 _14791_/X vssd1 vssd1 vccd1 vccd1 _18185_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07788_ _07788_/A vssd1 vssd1 vccd1 vccd1 _07788_/Y sky130_fd_sc_hd__inv_2
X_09527_ hold1853/X _13134_/A _10031_/C vssd1 vssd1 vccd1 vccd1 _09528_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_210_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_213_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ _09463_/C _09463_/D _09478_/B vssd1 vssd1 vccd1 vccd1 _09458_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_149_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08409_ hold933/X _08439_/B vssd1 vssd1 vccd1 vccd1 _08409_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09389_ _07805_/A _09362_/A _09362_/D vssd1 vssd1 vccd1 vccd1 _09389_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_191_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11420_ hold1167/X _16964_/Q _11741_/C vssd1 vssd1 vccd1 vccd1 _11421_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11351_ hold3059/X _16941_/Q _11738_/C vssd1 vssd1 vccd1 vccd1 _11352_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10302_ _10470_/A _10302_/B vssd1 vssd1 vccd1 vccd1 _10302_/X sky130_fd_sc_hd__or2_1
X_14070_ _14517_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14070_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_240_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11282_ hold1196/X hold4393/X _11660_/S vssd1 vssd1 vccd1 vccd1 _11283_/B sky130_fd_sc_hd__mux2_1
Xhold5260 _11665_/X vssd1 vssd1 vccd1 vccd1 _17045_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13021_ _13048_/A hold894/X hold704/X vssd1 vssd1 vccd1 vccd1 hold903/A sky130_fd_sc_hd__a21o_1
XFILLER_0_120_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10233_ _11088_/A _10233_/B vssd1 vssd1 vccd1 vccd1 _10233_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5271 _17018_/Q vssd1 vssd1 vccd1 vccd1 hold5271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5282 _13645_/X vssd1 vssd1 vccd1 vccd1 _17668_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5293 _16940_/Q vssd1 vssd1 vccd1 vccd1 hold5293/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4570 _13639_/X vssd1 vssd1 vccd1 vccd1 _17666_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4581 _16436_/Q vssd1 vssd1 vccd1 vccd1 hold4581/X sky130_fd_sc_hd__dlygate4sd3_1
X_10164_ _10551_/A _10164_/B vssd1 vssd1 vccd1 vccd1 _10164_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4592 _09529_/X vssd1 vssd1 vccd1 vccd1 _16333_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_234_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_238_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3880 _16472_/Q vssd1 vssd1 vccd1 vccd1 hold3880/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3891 _10447_/X vssd1 vssd1 vccd1 vccd1 _16639_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14972_ _14972_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14972_/X sky130_fd_sc_hd__or2_1
X_10095_ _11109_/A _10095_/B vssd1 vssd1 vccd1 vccd1 _10095_/X sky130_fd_sc_hd__or2_1
X_17760_ _17867_/CLK _17760_/D vssd1 vssd1 vccd1 vccd1 hold957/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_215_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16711_ _18010_/CLK _16711_/D vssd1 vssd1 vccd1 vccd1 _16711_/Q sky130_fd_sc_hd__dfxtp_1
X_13923_ _13923_/A _13923_/B vssd1 vssd1 vccd1 vccd1 _17769_/D sky130_fd_sc_hd__and2_1
X_17691_ _17723_/CLK _17691_/D vssd1 vssd1 vccd1 vccd1 _17691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16642_ _18200_/CLK _16642_/D vssd1 vssd1 vccd1 vccd1 _16642_/Q sky130_fd_sc_hd__dfxtp_1
X_13854_ hold4421/X _13758_/A _13853_/X vssd1 vssd1 vccd1 vccd1 _13854_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_236_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12805_ hold2673/X _17446_/Q _12811_/S vssd1 vssd1 vccd1 vccd1 _12805_/X sky130_fd_sc_hd__mux2_1
X_16573_ _18099_/CLK _16573_/D vssd1 vssd1 vccd1 vccd1 _16573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13785_ _13791_/A _13785_/B vssd1 vssd1 vccd1 vccd1 _13785_/X sky130_fd_sc_hd__or2_1
XFILLER_0_230_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10997_ hold2328/X hold4993/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10998_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18312_ _18375_/CLK _18312_/D vssd1 vssd1 vccd1 vccd1 hold833/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15524_ hold1414/X _15560_/A2 _15523_/X _12849_/A vssd1 vssd1 vccd1 vccd1 _15524_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ hold1668/X _17423_/Q _12811_/S vssd1 vssd1 vccd1 vccd1 _12736_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_365_wb_clk_i clkbuf_6_34_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17672_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18243_ _18271_/CLK _18243_/D vssd1 vssd1 vccd1 vccd1 _18243_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15455_ hold565/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15455_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ hold2472/X hold3122/X _12850_/S vssd1 vssd1 vccd1 vccd1 _12667_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_154_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14406_ hold2707/X _14446_/A2 _14405_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _14406_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18174_ _18174_/CLK _18174_/D vssd1 vssd1 vccd1 vccd1 _18174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11618_ hold2460/X hold4119/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11619_/B sky130_fd_sc_hd__mux2_1
X_15386_ _17342_/Q _15486_/B1 _09362_/D hold175/X vssd1 vssd1 vccd1 vccd1 _15386_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12598_ hold1696/X hold3286/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12598_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17125_ _17157_/CLK _17125_/D vssd1 vssd1 vccd1 vccd1 _17125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14337_ hold1583/X _14326_/B _14336_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14337_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11549_ hold2489/X _17007_/Q _11741_/C vssd1 vssd1 vccd1 vccd1 _11550_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold507 hold507/A vssd1 vssd1 vccd1 vccd1 input58/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 hold518/A vssd1 vssd1 vccd1 vccd1 hold518/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold529 hold529/A vssd1 vssd1 vccd1 vccd1 hold529/X sky130_fd_sc_hd__dlygate4sd3_1
X_17056_ _17904_/CLK _17056_/D vssd1 vssd1 vccd1 vccd1 _17056_/Q sky130_fd_sc_hd__dfxtp_1
X_14268_ _15163_/A _14268_/B vssd1 vssd1 vccd1 vccd1 _14268_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_204_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16007_ _18418_/CLK _16007_/D vssd1 vssd1 vccd1 vccd1 hold400/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13219_ _13218_/X hold5998/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13219_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_209_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ hold2308/X _14198_/B _14198_/Y _13933_/A vssd1 vssd1 vccd1 vccd1 _14199_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1207 _15852_/Q vssd1 vssd1 vccd1 vccd1 hold1207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08760_ _15274_/A _08760_/B vssd1 vssd1 vccd1 vccd1 _16000_/D sky130_fd_sc_hd__and2_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17958_ _17967_/CLK _17958_/D vssd1 vssd1 vccd1 vccd1 _17958_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1218 _15796_/Q vssd1 vssd1 vccd1 vccd1 hold1218/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_81_wb_clk_i clkbuf_6_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17486_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1229 _15648_/Q vssd1 vssd1 vccd1 vccd1 hold1229/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_240_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16909_ _17885_/CLK _16909_/D vssd1 vssd1 vccd1 vccd1 _16909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08691_ hold169/X hold608/X _08721_/S vssd1 vssd1 vccd1 vccd1 hold609/A sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_240_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_10_wb_clk_i clkbuf_6_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17194_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17889_ _17889_/CLK _17889_/D vssd1 vssd1 vccd1 vccd1 _17889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09312_ hold2846/X _09323_/B _09311_/X _14358_/A vssd1 vssd1 vccd1 vccd1 _09312_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09243_ _15519_/A hold917/X _09283_/S vssd1 vssd1 vccd1 vccd1 hold918/A sky130_fd_sc_hd__mux2_1
XFILLER_0_63_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09174_ _15557_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09174_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08125_ _08125_/A _08125_/B vssd1 vssd1 vccd1 vccd1 _15701_/D sky130_fd_sc_hd__and2_1
XFILLER_0_181_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08056_ _15515_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08056_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3110 _18030_/Q vssd1 vssd1 vccd1 vccd1 hold3110/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3121 _12872_/X vssd1 vssd1 vccd1 vccd1 _12873_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3132 _12587_/X vssd1 vssd1 vccd1 vccd1 _12588_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3143 _17395_/Q vssd1 vssd1 vccd1 vccd1 hold3143/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3154 _17402_/Q vssd1 vssd1 vccd1 vccd1 hold3154/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2420 _15769_/Q vssd1 vssd1 vccd1 vccd1 hold2420/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3165 _17420_/Q vssd1 vssd1 vccd1 vccd1 hold3165/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3176 _12749_/X vssd1 vssd1 vccd1 vccd1 _12750_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2431 _15591_/Q vssd1 vssd1 vccd1 vccd1 hold2431/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08958_ _15473_/A hold164/X vssd1 vssd1 vccd1 vccd1 _16096_/D sky130_fd_sc_hd__and2_1
XFILLER_0_208_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2442 _14585_/X vssd1 vssd1 vccd1 vccd1 _18086_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3187 _15190_/X vssd1 vssd1 vccd1 vccd1 _18377_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3198 _10038_/Y vssd1 vssd1 vccd1 vccd1 _10039_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2453 _15635_/Q vssd1 vssd1 vccd1 vccd1 hold2453/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2464 _16195_/Q vssd1 vssd1 vccd1 vccd1 hold2464/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1730 _18082_/Q vssd1 vssd1 vccd1 vccd1 hold1730/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2475 _07923_/X vssd1 vssd1 vccd1 vccd1 _15605_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2486 _14745_/X vssd1 vssd1 vccd1 vccd1 _18163_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1741 _07860_/X vssd1 vssd1 vccd1 vccd1 _15575_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07909_ hold1323/X _07918_/B _07908_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _07909_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1752 _15628_/Q vssd1 vssd1 vccd1 vccd1 hold1752/X sky130_fd_sc_hd__dlygate4sd3_1
X_08889_ _12416_/A hold826/X vssd1 vssd1 vccd1 vccd1 _16062_/D sky130_fd_sc_hd__and2_1
Xhold2497 _18243_/Q vssd1 vssd1 vccd1 vccd1 hold2497/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_224_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1763 _07858_/X vssd1 vssd1 vccd1 vccd1 _15574_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1774 _08288_/X vssd1 vssd1 vccd1 vccd1 _15777_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1785 _18173_/Q vssd1 vssd1 vccd1 vccd1 hold1785/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10920_ _11694_/A _10920_/B vssd1 vssd1 vccd1 vccd1 _10920_/X sky130_fd_sc_hd__or2_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1796 _08257_/X vssd1 vssd1 vccd1 vccd1 _15763_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10851_ _11637_/A _10851_/B vssd1 vssd1 vccd1 vccd1 _10851_/X sky130_fd_sc_hd__or2_1
XFILLER_0_233_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13570_ hold5476/X _13847_/B _13569_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13570_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _11655_/A _10782_/B vssd1 vssd1 vccd1 vccd1 _10782_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12521_ hold4511/X _12520_/X _12929_/S vssd1 vssd1 vccd1 vccd1 _12522_/B sky130_fd_sc_hd__mux2_1
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ hold582/X _15448_/A2 _15446_/B1 hold647/X vssd1 vssd1 vccd1 vccd1 _15240_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ _17319_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12452_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11403_ _12234_/A _11403_/B vssd1 vssd1 vccd1 vccd1 _11403_/X sky130_fd_sc_hd__or2_1
X_15171_ hold991/A _15179_/B vssd1 vssd1 vccd1 vccd1 hold842/A sky130_fd_sc_hd__or2_1
XFILLER_0_152_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12383_ hold618/X hold808/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold809/A sky130_fd_sc_hd__mux2_1
XFILLER_0_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14122_ _14461_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14122_/X sky130_fd_sc_hd__or2_1
X_11334_ _12210_/A _11334_/B vssd1 vssd1 vccd1 vccd1 _11334_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14053_ hold1035/X _14040_/B _14052_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _14053_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11265_ _12285_/A _11265_/B vssd1 vssd1 vccd1 vccd1 _11265_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5090 _17221_/Q vssd1 vssd1 vccd1 vccd1 hold5090/X sky130_fd_sc_hd__dlygate4sd3_1
X_13004_ _14897_/A hold363/X vssd1 vssd1 vccd1 vccd1 _13017_/B sky130_fd_sc_hd__or2_2
X_10216_ hold3670/X _10598_/B _10215_/X _14895_/C1 vssd1 vssd1 vccd1 vccd1 _10216_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11196_ hold3590/X _11100_/A _11195_/X vssd1 vssd1 vccd1 vccd1 _11196_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17812_ _17856_/CLK _17812_/D vssd1 vssd1 vccd1 vccd1 _17812_/Q sky130_fd_sc_hd__dfxtp_1
X_10147_ hold3700/X _10589_/B _10146_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _10147_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14955_ hold6080/X _14946_/B hold240/X _15030_/A vssd1 vssd1 vccd1 vccd1 hold241/A
+ sky130_fd_sc_hd__o211a_1
XTAP_5883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17743_ _17743_/CLK _17743_/D vssd1 vssd1 vccd1 vccd1 _17743_/Q sky130_fd_sc_hd__dfxtp_1
X_10078_ hold3595/X _10598_/B _10077_/X _15218_/C1 vssd1 vssd1 vccd1 vccd1 _10078_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_216_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13906_ _14461_/A hold2764/X hold297/X vssd1 vssd1 vccd1 vccd1 _13907_/B sky130_fd_sc_hd__mux2_1
X_14886_ _15225_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14886_/X sky130_fd_sc_hd__or2_1
X_17674_ _17738_/CLK _17674_/D vssd1 vssd1 vccd1 vccd1 _17674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16625_ _18197_/CLK _16625_/D vssd1 vssd1 vccd1 vccd1 _16625_/Q sky130_fd_sc_hd__dfxtp_1
X_13837_ _13873_/A _13837_/B vssd1 vssd1 vccd1 vccd1 _13837_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_230_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16556_ _18212_/CLK _16556_/D vssd1 vssd1 vccd1 vccd1 _16556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13768_ _13862_/A _13795_/A2 _13767_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13768_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12719_ hold3783/X _12718_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12719_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15507_ hold445/X hold363/X vssd1 vssd1 vccd1 vccd1 _15507_/Y sky130_fd_sc_hd__nor2_1
X_16487_ _18240_/CLK _16487_/D vssd1 vssd1 vccd1 vccd1 _16487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13699_ hold4658/X _13795_/A2 _13698_/X _13795_/C1 vssd1 vssd1 vccd1 vccd1 _13699_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15438_ hold777/X _09367_/A _09362_/C _17347_/Q vssd1 vssd1 vccd1 vccd1 _15438_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_216_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18226_ _18226_/CLK _18226_/D vssd1 vssd1 vccd1 vccd1 _18226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18157_ _18221_/CLK _18157_/D vssd1 vssd1 vccd1 vccd1 _18157_/Q sky130_fd_sc_hd__dfxtp_1
X_15369_ hold174/X _15485_/A2 _15488_/A2 hold153/X _15368_/X vssd1 vssd1 vccd1 vccd1
+ _15372_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_14_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold304 hold441/X vssd1 vssd1 vccd1 vccd1 hold442/A sky130_fd_sc_hd__dlygate4sd3_1
X_17108_ _17270_/CLK _17108_/D vssd1 vssd1 vccd1 vccd1 _17108_/Q sky130_fd_sc_hd__dfxtp_1
Xhold315 hold35/X vssd1 vssd1 vccd1 vccd1 hold315/X sky130_fd_sc_hd__clkbuf_4
X_18088_ _18106_/CLK _18088_/D vssd1 vssd1 vccd1 vccd1 _18088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold326 hold326/A vssd1 vssd1 vccd1 vccd1 hold326/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold337 hold337/A vssd1 vssd1 vccd1 vccd1 hold337/X sky130_fd_sc_hd__clkbuf_4
Xhold348 hold348/A vssd1 vssd1 vccd1 vccd1 hold348/X sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ _09948_/A _09930_/B vssd1 vssd1 vccd1 vccd1 _09930_/X sky130_fd_sc_hd__or2_1
XFILLER_0_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17039_ _17887_/CLK _17039_/D vssd1 vssd1 vccd1 vccd1 _17039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold359 hold359/A vssd1 vssd1 vccd1 vccd1 input61/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout806 fanout816/X vssd1 vssd1 vccd1 vccd1 _15066_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09861_ _09957_/A _09861_/B vssd1 vssd1 vccd1 vccd1 _09861_/X sky130_fd_sc_hd__or2_1
Xfanout817 _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14867_/C1 sky130_fd_sc_hd__buf_4
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout828 _14863_/C1 vssd1 vssd1 vccd1 vccd1 _14883_/C1 sky130_fd_sc_hd__clkbuf_8
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout839 fanout843/X vssd1 vssd1 vccd1 vccd1 _14691_/C1 sky130_fd_sc_hd__clkbuf_4
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ hold71/X hold845/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08813_/B sky130_fd_sc_hd__mux2_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _09912_/A _09792_/B vssd1 vssd1 vccd1 vccd1 _09792_/X sky130_fd_sc_hd__or2_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1004 la_data_in[11] vssd1 vssd1 vccd1 vccd1 hold519/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 _15696_/Q vssd1 vssd1 vccd1 vccd1 hold1015/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 _07842_/X vssd1 vssd1 vccd1 vccd1 _15566_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08743_ hold29/X hold544/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08744_/B sky130_fd_sc_hd__mux2_1
Xhold1037 _15783_/Q vssd1 vssd1 vccd1 vccd1 hold1037/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1048 _14249_/X vssd1 vssd1 vccd1 vccd1 _17925_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1059 _14721_/X vssd1 vssd1 vccd1 vccd1 _18152_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08674_ _15491_/A hold260/X vssd1 vssd1 vccd1 vccd1 _15958_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_287_wb_clk_i clkbuf_6_48_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17967_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_216_wb_clk_i clkbuf_6_60_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18115_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09226_ _15555_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09226_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09157_ hold2181/X _09164_/B _09156_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _09157_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08108_ _15513_/A hold2966/X hold108/X vssd1 vssd1 vccd1 vccd1 _08109_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09088_ _14988_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _09088_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08039_ _14726_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08039_/X sky130_fd_sc_hd__or2_1
XFILLER_0_101_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold860 hold860/A vssd1 vssd1 vccd1 vccd1 hold860/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 hold871/A vssd1 vssd1 vccd1 vccd1 hold871/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 hold882/A vssd1 vssd1 vccd1 vccd1 hold882/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 hold900/X vssd1 vssd1 vccd1 vccd1 hold901/A sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ hold3791/X _11144_/B _11049_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _11050_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10001_ _16491_/Q _10025_/B _10025_/C vssd1 vssd1 vccd1 vccd1 _10001_/X sky130_fd_sc_hd__and3_1
XFILLER_0_219_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2250 becStatus[3] vssd1 vssd1 vccd1 vccd1 hold919/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2261 _18219_/Q vssd1 vssd1 vccd1 vccd1 hold2261/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2272 _12626_/S vssd1 vssd1 vccd1 vccd1 hold2272/X sky130_fd_sc_hd__buf_2
Xhold2283 _14591_/X vssd1 vssd1 vccd1 vccd1 _18089_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2294 _08085_/X vssd1 vssd1 vccd1 vccd1 _15682_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1560 _17883_/Q vssd1 vssd1 vccd1 vccd1 hold1560/X sky130_fd_sc_hd__dlygate4sd3_1
X_14740_ _15187_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14740_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1571 _14139_/X vssd1 vssd1 vccd1 vccd1 _17873_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11952_ _12240_/A _11952_/B vssd1 vssd1 vccd1 vccd1 _11952_/X sky130_fd_sc_hd__or2_1
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1582 _14171_/X vssd1 vssd1 vccd1 vccd1 _17888_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1593 _14331_/X vssd1 vssd1 vccd1 vccd1 _17965_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10903_ hold4993/X _10616_/B _10902_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _10903_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14671_ hold2073/X _14664_/B _14670_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14671_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _12267_/A _11883_/B vssd1 vssd1 vccd1 vccd1 _11883_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16410_ _18323_/CLK _16410_/D vssd1 vssd1 vccd1 vccd1 _16410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13622_ hold2357/X hold5767/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13623_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_233_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10834_ hold5353/X _11225_/B _10833_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _10834_/X
+ sky130_fd_sc_hd__o211a_1
X_17390_ _18453_/CLK _17390_/D vssd1 vssd1 vccd1 vccd1 _17390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16341_ _18356_/CLK _16341_/D vssd1 vssd1 vccd1 vccd1 _16341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13553_ hold1226/X hold5597/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13554_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_211_1372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10765_ hold3985/X _11144_/B _10764_/X _14354_/A vssd1 vssd1 vccd1 vccd1 _10765_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12504_ _17345_/Q _12506_/B vssd1 vssd1 vccd1 vccd1 _12504_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16272_ _17374_/CLK _16272_/D vssd1 vssd1 vccd1 vccd1 _16272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13484_ hold1207/X _17615_/Q _13841_/C vssd1 vssd1 vccd1 vccd1 _13485_/B sky130_fd_sc_hd__mux2_1
X_10696_ hold4016/X _11753_/B _10695_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _10696_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15223_ hold484/X _15227_/B vssd1 vssd1 vccd1 vccd1 hold485/A sky130_fd_sc_hd__or2_1
XFILLER_0_180_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18011_ _18043_/CLK _18011_/D vssd1 vssd1 vccd1 vccd1 _18011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12435_ hold82/X hold118/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold119/A sky130_fd_sc_hd__mux2_1
XFILLER_0_81_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15154_ hold6082/X _15165_/B _15153_/X _15212_/C1 vssd1 vssd1 vccd1 vccd1 _15154_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12366_ hold3496/X _13749_/A _12365_/X vssd1 vssd1 vccd1 vccd1 _12366_/Y sky130_fd_sc_hd__a21oi_1
X_14105_ hold1393/X _14094_/B _14104_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _14105_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11317_ hold5585/X _12335_/B _11316_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11317_/X
+ sky130_fd_sc_hd__o211a_1
X_15085_ _15085_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15085_/X sky130_fd_sc_hd__or2_1
XFILLER_0_61_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12297_ hold4323/X _13716_/A _12296_/X vssd1 vssd1 vccd1 vccd1 _12297_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_238_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14036_ _15543_/A _14038_/B vssd1 vssd1 vccd1 vccd1 _14036_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_226_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11248_ hold5434/X _11726_/B _11247_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _11248_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11179_ _11206_/A _11179_/B vssd1 vssd1 vccd1 vccd1 _16883_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_101_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15987_ _16098_/CLK _15987_/D vssd1 vssd1 vccd1 vccd1 hold854/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17726_ _17726_/CLK _17726_/D vssd1 vssd1 vccd1 vccd1 _17726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14938_ _15207_/A hold407/X vssd1 vssd1 vccd1 vccd1 _14938_/X sky130_fd_sc_hd__or2_1
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_380_wb_clk_i clkbuf_6_33_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17244_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17657_ _17722_/CLK _17657_/D vssd1 vssd1 vccd1 vccd1 _17657_/Q sky130_fd_sc_hd__dfxtp_1
X_14869_ hold2958/X _14880_/B _14868_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14869_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16608_ _18231_/CLK _16608_/D vssd1 vssd1 vccd1 vccd1 _16608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08390_ _14732_/A hold940/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08391_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_175_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17588_ _17620_/CLK _17588_/D vssd1 vssd1 vccd1 vccd1 _17588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16539_ _18115_/CLK _16539_/D vssd1 vssd1 vccd1 vccd1 _16539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09011_ _12420_/A _09011_/B vssd1 vssd1 vccd1 vccd1 _16122_/D sky130_fd_sc_hd__and2_1
XFILLER_0_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18209_ _18217_/CLK _18209_/D vssd1 vssd1 vccd1 vccd1 _18209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5804 _12136_/X vssd1 vssd1 vccd1 vccd1 _17202_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5815 _17594_/Q vssd1 vssd1 vccd1 vccd1 hold5815/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold101 hold101/A vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5826 _09532_/X vssd1 vssd1 vccd1 vccd1 _16334_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold112 hold508/X vssd1 vssd1 vccd1 vccd1 hold509/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_227_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold123 hold123/A vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5837 _16368_/Q vssd1 vssd1 vccd1 vccd1 hold5837/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5848 output87/X vssd1 vssd1 vccd1 vccd1 data_out[23] sky130_fd_sc_hd__buf_12
Xhold5859 hold6012/X vssd1 vssd1 vccd1 vccd1 _13185_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 hold617/X vssd1 vssd1 vccd1 vccd1 hold618/A sky130_fd_sc_hd__buf_1
XFILLER_0_130_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold145 hold145/A vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold156 hold156/A vssd1 vssd1 vccd1 vccd1 hold156/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold167 hold58/X vssd1 vssd1 vccd1 vccd1 input9/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 hold10/X vssd1 vssd1 vccd1 vccd1 input11/A sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ hold3580/X _10025_/B _09912_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09913_/X
+ sky130_fd_sc_hd__o211a_1
Xhold189 hold189/A vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _09484_/B vssd1 vssd1 vccd1 vccd1 _09478_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout614 _09358_/Y vssd1 vssd1 vccd1 vccd1 _15487_/B1 sky130_fd_sc_hd__buf_6
XFILLER_0_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout625 _09347_/Y vssd1 vssd1 vccd1 vccd1 _15484_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout636 _12798_/A vssd1 vssd1 vccd1 vccd1 _12810_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09844_ hold5835/X _10022_/B _09843_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09844_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout647 _12199_/C1 vssd1 vssd1 vccd1 vccd1 _12103_/C1 sky130_fd_sc_hd__buf_2
Xfanout658 _12588_/A vssd1 vssd1 vccd1 vccd1 _12660_/A sky130_fd_sc_hd__buf_4
Xfanout669 fanout689/X vssd1 vssd1 vccd1 vccd1 _08171_/A sky130_fd_sc_hd__clkbuf_4
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ hold3604/X _10049_/B _09774_/X _15212_/C1 vssd1 vssd1 vccd1 vccd1 _09775_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08726_ _15434_/A _08726_/B vssd1 vssd1 vccd1 vccd1 _15984_/D sky130_fd_sc_hd__and2_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ hold495/X hold668/X _08657_/S vssd1 vssd1 vccd1 vccd1 hold669/A sky130_fd_sc_hd__mux2_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ hold87/X hold473/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold474/A sky130_fd_sc_hd__mux2_1
XFILLER_0_165_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10550_ hold1801/X hold4602/X _10646_/C vssd1 vssd1 vccd1 vccd1 _10551_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09209_ hold1666/X _09214_/B _09208_/X _12822_/A vssd1 vssd1 vccd1 vccd1 _09209_/X
+ sky130_fd_sc_hd__o211a_1
X_10481_ hold1750/X hold3282/X _10601_/C vssd1 vssd1 vccd1 vccd1 _10482_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12220_ hold5458/X _12323_/B _12219_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _12220_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_6_42_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_42_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12151_ hold4037/X _12365_/B _12150_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _12151_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11102_ hold1684/X _16858_/Q _11213_/C vssd1 vssd1 vccd1 vccd1 _11103_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_208_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12082_ hold5137/X _13886_/B _12081_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _17184_/D
+ sky130_fd_sc_hd__o211a_1
Xhold690 hold690/A vssd1 vssd1 vccd1 vccd1 hold690/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_229_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15910_ _18401_/CLK _15910_/D vssd1 vssd1 vccd1 vccd1 hold639/A sky130_fd_sc_hd__dfxtp_1
X_11033_ hold2693/X hold3927/X _11765_/C vssd1 vssd1 vccd1 vccd1 _11034_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16890_ _18005_/CLK _16890_/D vssd1 vssd1 vccd1 vccd1 _16890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _17648_/CLK _15841_/D vssd1 vssd1 vccd1 vccd1 _15841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2080 _14083_/X vssd1 vssd1 vccd1 vccd1 _17846_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_138_wb_clk_i clkbuf_6_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16124_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2091 _14057_/X vssd1 vssd1 vccd1 vccd1 _17833_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ _12984_/A _12984_/B vssd1 vssd1 vccd1 vccd1 _17504_/D sky130_fd_sc_hd__and2_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ _17723_/CLK _15772_/D vssd1 vssd1 vccd1 vccd1 _15772_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1390 input2/X vssd1 vssd1 vccd1 vccd1 _13019_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17511_ _17512_/CLK _17511_/D vssd1 vssd1 vccd1 vccd1 _17511_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14723_ hold1994/X _14718_/B _14722_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14723_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11935_ hold5129/X _12317_/B _11934_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _11935_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14654_ _15209_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14654_/X sky130_fd_sc_hd__or2_1
X_17442_ _17445_/CLK _17442_/D vssd1 vssd1 vccd1 vccd1 _17442_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11866_ hold3976/X _12374_/B _11865_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _11866_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13605_ _13722_/A _13605_/B vssd1 vssd1 vccd1 vccd1 _13605_/X sky130_fd_sc_hd__or2_1
XFILLER_0_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10817_ hold1448/X hold3844/X _11171_/C vssd1 vssd1 vccd1 vccd1 _10818_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14585_ hold2441/X _14612_/B _14584_/X _15218_/C1 vssd1 vssd1 vccd1 vccd1 _14585_/X
+ sky130_fd_sc_hd__o211a_1
X_17373_ _17374_/CLK _17373_/D vssd1 vssd1 vccd1 vccd1 _17373_/Q sky130_fd_sc_hd__dfxtp_1
X_11797_ _12337_/A _11797_/B vssd1 vssd1 vccd1 vccd1 _11797_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_184_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16324_ _18399_/CLK _16324_/D vssd1 vssd1 vccd1 vccd1 _16324_/Q sky130_fd_sc_hd__dfxtp_1
X_13536_ _13737_/A _13536_/B vssd1 vssd1 vccd1 vccd1 _13536_/X sky130_fd_sc_hd__or2_1
X_10748_ hold583/X hold3978/X _11168_/C vssd1 vssd1 vccd1 vccd1 _10749_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16255_ _17517_/CLK _16255_/D vssd1 vssd1 vccd1 vccd1 _16255_/Q sky130_fd_sc_hd__dfxtp_1
X_13467_ _13791_/A _13467_/B vssd1 vssd1 vccd1 vccd1 _13467_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10679_ hold1939/X hold4281/X _11162_/C vssd1 vssd1 vccd1 vccd1 _10680_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15206_ hold1821/X _15221_/B _15205_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _15206_/X
+ sky130_fd_sc_hd__o211a_1
X_12418_ _12418_/A _12418_/B vssd1 vssd1 vccd1 vccd1 _17302_/D sky130_fd_sc_hd__and2_1
XFILLER_0_3_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16186_ _18448_/CLK _16186_/D vssd1 vssd1 vccd1 vccd1 _16186_/Q sky130_fd_sc_hd__dfxtp_1
X_13398_ _13791_/A _13398_/B vssd1 vssd1 vccd1 vccd1 _13398_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15137_ _15191_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15137_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12349_ _13873_/A _12349_/B vssd1 vssd1 vccd1 vccd1 _12349_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_239_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3709 _09664_/X vssd1 vssd1 vccd1 vccd1 _16378_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15068_ _15068_/A _15068_/B vssd1 vssd1 vccd1 vccd1 _18319_/D sky130_fd_sc_hd__and2_1
XFILLER_0_103_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14019_ hold3114/X _14038_/B _14018_/X _12588_/A vssd1 vssd1 vccd1 vccd1 _14019_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07890_ hold911/X _07936_/B vssd1 vssd1 vccd1 vccd1 _07890_/X sky130_fd_sc_hd__or2_1
XFILLER_0_235_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218_1334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09560_ hold1988/X _13222_/A _10040_/C vssd1 vssd1 vccd1 vccd1 _09561_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08511_ _15515_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08511_/X sky130_fd_sc_hd__or2_1
XFILLER_0_218_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17709_ _17709_/CLK _17709_/D vssd1 vssd1 vccd1 vccd1 _17709_/Q sky130_fd_sc_hd__dfxtp_1
X_09491_ _17520_/Q _13034_/D vssd1 vssd1 vccd1 vccd1 _13056_/D sky130_fd_sc_hd__nand2_2
XFILLER_0_72_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08442_ hold1564/X _08442_/A2 _08441_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _08442_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_1400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08373_ _08373_/A hold230/X vssd1 vssd1 vccd1 vccd1 hold231/A sky130_fd_sc_hd__and2_1
XFILLER_0_191_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_1327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5601 _17188_/Q vssd1 vssd1 vccd1 vccd1 hold5601/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5612 _17163_/Q vssd1 vssd1 vccd1 vccd1 hold5612/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5623 _11650_/X vssd1 vssd1 vccd1 vccd1 _17040_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5634 _11278_/X vssd1 vssd1 vccd1 vccd1 _16916_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4900 _10669_/X vssd1 vssd1 vccd1 vccd1 _16713_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5645 _16947_/Q vssd1 vssd1 vccd1 vccd1 hold5645/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4911 _16822_/Q vssd1 vssd1 vccd1 vccd1 hold4911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5656 _11497_/X vssd1 vssd1 vccd1 vccd1 _16989_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4922 _12274_/X vssd1 vssd1 vccd1 vccd1 _17248_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5667 _17075_/Q vssd1 vssd1 vccd1 vccd1 hold5667/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5678 _11593_/X vssd1 vssd1 vccd1 vccd1 _17021_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4933 _16959_/Q vssd1 vssd1 vccd1 vccd1 hold4933/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4944 _13606_/X vssd1 vssd1 vccd1 vccd1 _17655_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5689 _17257_/Q vssd1 vssd1 vccd1 vccd1 hold5689/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4955 _16828_/Q vssd1 vssd1 vccd1 vccd1 hold4955/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout400 _14447_/Y vssd1 vssd1 vccd1 vccd1 _14481_/B sky130_fd_sc_hd__buf_6
Xhold4966 _17155_/Q vssd1 vssd1 vccd1 vccd1 hold4966/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4977 _11875_/X vssd1 vssd1 vccd1 vccd1 _17115_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout411 _14232_/Y vssd1 vssd1 vccd1 vccd1 _14272_/B sky130_fd_sc_hd__clkbuf_8
Xhold4988 _12250_/X vssd1 vssd1 vccd1 vccd1 _17240_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout422 _14040_/B vssd1 vssd1 vccd1 vccd1 _14038_/B sky130_fd_sc_hd__buf_6
Xhold4999 _17364_/Q vssd1 vssd1 vccd1 vccd1 hold4999/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout433 _13311_/A1 vssd1 vssd1 vccd1 vccd1 _13199_/A1 sky130_fd_sc_hd__buf_8
Xfanout444 _12227_/S vssd1 vssd1 vccd1 vccd1 _13409_/S sky130_fd_sc_hd__clkbuf_8
Xfanout455 fanout485/X vssd1 vssd1 vccd1 vccd1 _11741_/C sky130_fd_sc_hd__buf_4
Xfanout466 _13877_/C vssd1 vssd1 vccd1 vccd1 _13883_/C sky130_fd_sc_hd__buf_6
X_09827_ _18346_/Q hold3536/X _10067_/C vssd1 vssd1 vccd1 vccd1 _09828_/B sky130_fd_sc_hd__mux2_1
Xfanout477 _11210_/C vssd1 vssd1 vccd1 vccd1 _11660_/S sky130_fd_sc_hd__buf_6
XFILLER_0_214_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout488 _11201_/C vssd1 vssd1 vccd1 vccd1 _11162_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_241_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_213_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout499 _10985_/S vssd1 vssd1 vccd1 vccd1 _11186_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_216_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_231_wb_clk_i clkbuf_6_62_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18181_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09758_ hold1509/X _16410_/Q _10067_/C vssd1 vssd1 vccd1 vccd1 _09759_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08709_ hold53/X hold799/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08710_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ hold2297/X _16387_/Q _10601_/C vssd1 vssd1 vccd1 vccd1 _09690_/B sky130_fd_sc_hd__mux2_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _17064_/Q _12299_/B _12299_/C vssd1 vssd1 vccd1 vccd1 _11720_/X sky130_fd_sc_hd__and3_1
XFILLER_0_139_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11651_ hold2505/X hold5253/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11652_/B sky130_fd_sc_hd__mux2_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10602_ _16531_/Q _10482_/A _10601_/X vssd1 vssd1 vccd1 vccd1 _10602_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_194_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14370_ _15044_/A _14370_/B vssd1 vssd1 vccd1 vccd1 _17984_/D sky130_fd_sc_hd__and2_1
XFILLER_0_25_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11582_ hold1070/X _17018_/Q _12242_/S vssd1 vssd1 vccd1 vccd1 _11583_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13321_ hold4963/X _13814_/B _13320_/X _13417_/C1 vssd1 vssd1 vccd1 vccd1 _13321_/X
+ sky130_fd_sc_hd__o211a_1
X_10533_ _11103_/A _10533_/B vssd1 vssd1 vccd1 vccd1 _10533_/X sky130_fd_sc_hd__or2_1
XFILLER_0_88_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16040_ _18425_/CLK _16040_/D vssd1 vssd1 vccd1 vccd1 hold601/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13252_ hold4326/X _13251_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13252_/X sky130_fd_sc_hd__mux2_2
X_10464_ _10560_/A _10464_/B vssd1 vssd1 vccd1 vccd1 _10464_/X sky130_fd_sc_hd__or2_1
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12203_ hold3027/X hold5681/X _12299_/C vssd1 vssd1 vccd1 vccd1 _12204_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_122_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13183_ _13199_/A1 _13181_/X _13182_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13183_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10395_ _10554_/A _10395_/B vssd1 vssd1 vccd1 vccd1 _10395_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12134_ hold1103/X _17202_/Q _12362_/C vssd1 vssd1 vccd1 vccd1 _12135_/B sky130_fd_sc_hd__mux2_1
X_17991_ _18023_/CLK _17991_/D vssd1 vssd1 vccd1 vccd1 _17991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_319_wb_clk_i clkbuf_6_47_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17861_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12065_ hold3041/X _17179_/Q _13409_/S vssd1 vssd1 vccd1 vccd1 _12066_/B sky130_fd_sc_hd__mux2_1
X_16942_ _17886_/CLK _16942_/D vssd1 vssd1 vccd1 vccd1 _16942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11016_ _11694_/A _11016_/B vssd1 vssd1 vccd1 vccd1 _11016_/X sky130_fd_sc_hd__or2_1
XFILLER_0_223_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16873_ _18014_/CLK _16873_/D vssd1 vssd1 vccd1 vccd1 _16873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15824_ _17639_/CLK _15824_/D vssd1 vssd1 vccd1 vccd1 _15824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ hold1702/X hold3222/X _12970_/S vssd1 vssd1 vccd1 vccd1 _12967_/X sky130_fd_sc_hd__mux2_1
X_15755_ _17740_/CLK _15755_/D vssd1 vssd1 vccd1 vccd1 _15755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ _15099_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14706_/X sky130_fd_sc_hd__or2_1
X_11918_ hold1277/X _17130_/Q _12293_/C vssd1 vssd1 vccd1 vccd1 _11919_/B sky130_fd_sc_hd__mux2_1
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15686_ _17608_/CLK _15686_/D vssd1 vssd1 vccd1 vccd1 _15686_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12898_ hold2562/X hold3305/X _12916_/S vssd1 vssd1 vccd1 vccd1 _12898_/X sky130_fd_sc_hd__mux2_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ _17425_/CLK _17425_/D vssd1 vssd1 vccd1 vccd1 _17425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14637_ hold2516/X _14664_/B _14636_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _14637_/X
+ sky130_fd_sc_hd__o211a_1
X_11849_ hold3124/X hold4722/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11850_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14568_ _15492_/A _14573_/B hold2241/X vssd1 vssd1 vccd1 vccd1 _14568_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17356_ _17486_/CLK _17356_/D vssd1 vssd1 vccd1 vccd1 _17356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_wb_clk_i clkbuf_6_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17882_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_144_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16307_ _16315_/CLK _16307_/D vssd1 vssd1 vccd1 vccd1 _16307_/Q sky130_fd_sc_hd__dfxtp_1
X_13519_ hold3967/X _13808_/B _13518_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _13519_/X
+ sky130_fd_sc_hd__o211a_1
X_17287_ _18410_/CLK _17287_/D vssd1 vssd1 vccd1 vccd1 hold847/A sky130_fd_sc_hd__dfxtp_1
X_14499_ hold579/X _14499_/B vssd1 vssd1 vccd1 vccd1 _14499_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16238_ _17427_/CLK _16238_/D vssd1 vssd1 vccd1 vccd1 _16238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4207 _16016_/Q vssd1 vssd1 vccd1 vccd1 _15465_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4218 _15373_/X vssd1 vssd1 vccd1 vccd1 _15374_/B sky130_fd_sc_hd__dlygate4sd3_1
X_16169_ _17506_/CLK _16169_/D vssd1 vssd1 vccd1 vccd1 _16169_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4229 _10645_/Y vssd1 vssd1 vccd1 vccd1 _16705_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3506 _12372_/Y vssd1 vssd1 vccd1 vccd1 _12373_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08991_ hold87/X hold100/X _08991_/S vssd1 vssd1 vccd1 vccd1 hold101/A sky130_fd_sc_hd__mux2_1
Xhold3517 _16730_/Q vssd1 vssd1 vccd1 vccd1 hold3517/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3528 _13848_/Y vssd1 vssd1 vccd1 vccd1 _13849_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3539 _11724_/Y vssd1 vssd1 vccd1 vccd1 _11725_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2805 _18006_/Q vssd1 vssd1 vccd1 vccd1 hold2805/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2816 _14727_/X vssd1 vssd1 vccd1 vccd1 _18155_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07942_ hold915/X _07986_/B vssd1 vssd1 vccd1 vccd1 _07942_/X sky130_fd_sc_hd__or2_1
Xhold2827 _08457_/X vssd1 vssd1 vccd1 vccd1 _15857_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2838 _18266_/Q vssd1 vssd1 vccd1 vccd1 hold2838/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2849 _08249_/X vssd1 vssd1 vccd1 vccd1 _15759_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07873_ _14330_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07873_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09612_ _09933_/A _09612_/B vssd1 vssd1 vccd1 vccd1 _09612_/X sky130_fd_sc_hd__or2_1
XFILLER_0_190_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_222_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_218_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09543_ _09981_/A _09543_/B vssd1 vssd1 vccd1 vccd1 _09543_/X sky130_fd_sc_hd__or2_1
XFILLER_0_116_1416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09474_ _09477_/B _09477_/C _09478_/B vssd1 vssd1 vccd1 vccd1 _09474_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_231_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08425_ _14604_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08425_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08356_ _15525_/A hold3016/X hold115/X vssd1 vssd1 vccd1 vccd1 _08357_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08287_ hold915/X _08335_/B vssd1 vssd1 vccd1 vccd1 _08287_/X sky130_fd_sc_hd__or2_1
XFILLER_0_190_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6110 la_data_in[15] vssd1 vssd1 vccd1 vccd1 hold6110/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6121 la_data_in[5] vssd1 vssd1 vccd1 vccd1 hold420/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6132 _16517_/Q vssd1 vssd1 vccd1 vccd1 hold6132/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5420 _16664_/Q vssd1 vssd1 vccd1 vccd1 hold5420/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5431 _12037_/X vssd1 vssd1 vccd1 vccd1 _17169_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5442 _17259_/Q vssd1 vssd1 vccd1 vccd1 hold5442/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5453 _13471_/X vssd1 vssd1 vccd1 vccd1 _17610_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5464 _17747_/Q vssd1 vssd1 vccd1 vccd1 hold5464/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4730 _11065_/X vssd1 vssd1 vccd1 vccd1 _16845_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5475 _11452_/X vssd1 vssd1 vccd1 vccd1 _16974_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4741 _16441_/Q vssd1 vssd1 vccd1 vccd1 hold4741/X sky130_fd_sc_hd__dlygate4sd3_1
X_10180_ hold3876/X _10598_/B _10179_/X _10564_/C1 vssd1 vssd1 vccd1 vccd1 _10180_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5486 _17736_/Q vssd1 vssd1 vccd1 vccd1 hold5486/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5497 _13669_/X vssd1 vssd1 vccd1 vccd1 _17676_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4752 _11754_/Y vssd1 vssd1 vccd1 vccd1 _11755_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4763 _12300_/Y vssd1 vssd1 vccd1 vccd1 _12301_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4774 _09898_/X vssd1 vssd1 vccd1 vccd1 _16456_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_412_wb_clk_i clkbuf_6_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17908_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4785 _17623_/Q vssd1 vssd1 vccd1 vccd1 hold4785/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout230 _10634_/B vssd1 vssd1 vccd1 vccd1 _10616_/B sky130_fd_sc_hd__buf_4
Xhold4796 _12196_/X vssd1 vssd1 vccd1 vccd1 _17222_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout241 _10589_/B vssd1 vssd1 vccd1 vccd1 _10625_/B sky130_fd_sc_hd__buf_4
Xfanout252 _13800_/A vssd1 vssd1 vccd1 vccd1 _13797_/A sky130_fd_sc_hd__buf_4
Xfanout263 _11043_/A vssd1 vssd1 vccd1 vccd1 _11631_/A sky130_fd_sc_hd__buf_4
Xfanout274 _13581_/A vssd1 vssd1 vccd1 vccd1 _13752_/A sky130_fd_sc_hd__buf_4
Xfanout285 fanout299/X vssd1 vssd1 vccd1 vccd1 _12273_/A sky130_fd_sc_hd__buf_4
XFILLER_0_227_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout296 _11127_/A vssd1 vssd1 vccd1 vccd1 _11670_/A sky130_fd_sc_hd__buf_4
XFILLER_0_214_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13870_ _13873_/A _13870_/B vssd1 vssd1 vccd1 vccd1 _13870_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12821_ hold3136/X _12820_/X _12851_/S vssd1 vssd1 vccd1 vccd1 _12822_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_202_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ hold4039/X _12751_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12753_/B sky130_fd_sc_hd__mux2_1
X_15540_ hold2201/X _15547_/B _15539_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _15540_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_189_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11703_ _12174_/A _11703_/B vssd1 vssd1 vccd1 vccd1 _11703_/X sky130_fd_sc_hd__or2_1
X_15471_ _15480_/A _15471_/B _15471_/C _15471_/D vssd1 vssd1 vccd1 vccd1 _15471_/X
+ sky130_fd_sc_hd__or4_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ hold3376/X _12682_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12684_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14422_ hold2109/X _14433_/B _14421_/X _13895_/A vssd1 vssd1 vccd1 vccd1 _14422_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _17242_/CLK _17210_/D vssd1 vssd1 vccd1 vccd1 _17210_/Q sky130_fd_sc_hd__dfxtp_1
X_11634_ _11637_/A _11634_/B vssd1 vssd1 vccd1 vccd1 _11634_/X sky130_fd_sc_hd__or2_1
X_18190_ _18222_/CLK _18190_/D vssd1 vssd1 vccd1 vccd1 _18190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14353_ _14980_/A hold2901/X _14381_/S vssd1 vssd1 vccd1 vccd1 _14354_/B sky130_fd_sc_hd__mux2_1
X_17141_ _17779_/CLK _17141_/D vssd1 vssd1 vccd1 vccd1 _17141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11565_ _11661_/A _11565_/B vssd1 vssd1 vccd1 vccd1 _11565_/X sky130_fd_sc_hd__or2_1
X_13304_ _13297_/X _13303_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17556_/D sky130_fd_sc_hd__o21a_1
X_10516_ _10610_/A _10628_/B _10515_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10516_/X
+ sky130_fd_sc_hd__o211a_1
X_17072_ _17885_/CLK _17072_/D vssd1 vssd1 vccd1 vccd1 _17072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14284_ hold579/X _14284_/B vssd1 vssd1 vccd1 vccd1 _14284_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11496_ _12234_/A _11496_/B vssd1 vssd1 vccd1 vccd1 _11496_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16023_ _17325_/CLK _16023_/D vssd1 vssd1 vccd1 vccd1 hold136/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13235_ _13234_/X _16922_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13235_/X sky130_fd_sc_hd__mux2_1
X_10447_ hold3890/X _10631_/B _10446_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _10447_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13166_ _13166_/A _13294_/B vssd1 vssd1 vccd1 vccd1 _13166_/X sky130_fd_sc_hd__or2_1
X_10378_ hold3897/X _10568_/B _10377_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _10378_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_237_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_153_wb_clk_i clkbuf_6_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18424_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12117_ _13797_/A _12117_/B vssd1 vssd1 vccd1 vccd1 _12117_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13097_ _13097_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13097_/X sky130_fd_sc_hd__and2_1
X_17974_ _18036_/CLK _17974_/D vssd1 vssd1 vccd1 vccd1 _17974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_236_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12048_ _12240_/A _12048_/B vssd1 vssd1 vccd1 vccd1 _12048_/X sky130_fd_sc_hd__or2_1
X_16925_ _17894_/CLK _16925_/D vssd1 vssd1 vccd1 vccd1 _16925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16856_ _18059_/CLK _16856_/D vssd1 vssd1 vccd1 vccd1 _16856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15807_ _15856_/CLK _15807_/D vssd1 vssd1 vccd1 vccd1 hold963/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16787_ _18054_/CLK _16787_/D vssd1 vssd1 vccd1 vccd1 _16787_/Q sky130_fd_sc_hd__dfxtp_1
X_13999_ hold1085/X _13986_/B _13998_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _13999_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15738_ _17709_/CLK _15738_/D vssd1 vssd1 vccd1 vccd1 _15738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_1281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_213_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18457_ _18457_/CLK _18457_/D vssd1 vssd1 vccd1 vccd1 _18457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15669_ _17161_/CLK _15669_/D vssd1 vssd1 vccd1 vccd1 _15669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08210_ hold2304/X _08209_/B _08209_/Y _13777_/C1 vssd1 vssd1 vccd1 vccd1 _08210_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17408_ _17437_/CLK _17408_/D vssd1 vssd1 vccd1 vccd1 _17408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09190_ _15519_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09190_/X sky130_fd_sc_hd__or2_1
X_18388_ _18388_/CLK hold378/X vssd1 vssd1 vccd1 vccd1 _18388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08141_ _08143_/A hold356/X vssd1 vssd1 vccd1 vccd1 _15709_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17339_ _17339_/CLK hold66/X vssd1 vssd1 vccd1 vccd1 _17339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08072_ _15531_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08072_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4004 _13579_/X vssd1 vssd1 vccd1 vccd1 _17646_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4015 _17493_/Q vssd1 vssd1 vccd1 vccd1 hold4015/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4026 _17165_/Q vssd1 vssd1 vccd1 vccd1 hold4026/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4037 _17239_/Q vssd1 vssd1 vccd1 vccd1 hold4037/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3303 _16681_/Q vssd1 vssd1 vccd1 vccd1 _10571_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4048 _17710_/Q vssd1 vssd1 vccd1 vccd1 hold4048/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3314 _17484_/Q vssd1 vssd1 vccd1 vccd1 hold3314/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4059 _16786_/Q vssd1 vssd1 vccd1 vccd1 hold4059/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3325 _10774_/X vssd1 vssd1 vccd1 vccd1 _16748_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3336 _12884_/X vssd1 vssd1 vccd1 vccd1 _12885_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08974_ _12438_/A hold216/X vssd1 vssd1 vccd1 vccd1 _16104_/D sky130_fd_sc_hd__and2_1
Xhold3347 _16707_/Q vssd1 vssd1 vccd1 vccd1 hold3347/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2602 _14460_/X vssd1 vssd1 vccd1 vccd1 _18027_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2613 _18015_/Q vssd1 vssd1 vccd1 vccd1 hold2613/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3358 _12635_/X vssd1 vssd1 vccd1 vccd1 _12636_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2624 _14259_/X vssd1 vssd1 vccd1 vccd1 _17930_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3369 _12845_/X vssd1 vssd1 vccd1 vccd1 _12846_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2635 _17922_/Q vssd1 vssd1 vccd1 vccd1 hold2635/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1901 _18035_/Q vssd1 vssd1 vccd1 vccd1 hold1901/X sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ hold2512/X _07924_/B _07924_/Y _08167_/A vssd1 vssd1 vccd1 vccd1 _07925_/X
+ sky130_fd_sc_hd__o211a_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__buf_1
Xhold2646 _18018_/Q vssd1 vssd1 vccd1 vccd1 hold2646/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2657 _16182_/Q vssd1 vssd1 vccd1 vccd1 hold2657/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1912 _14025_/X vssd1 vssd1 vccd1 vccd1 _17818_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2668 _18301_/Q vssd1 vssd1 vccd1 vccd1 hold2668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1923 _16222_/Q vssd1 vssd1 vccd1 vccd1 hold1923/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2679 _18145_/Q vssd1 vssd1 vccd1 vccd1 hold2679/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1934 _14426_/X vssd1 vssd1 vccd1 vccd1 _18011_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1945 _15607_/Q vssd1 vssd1 vccd1 vccd1 hold1945/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1956 _18043_/Q vssd1 vssd1 vccd1 vccd1 hold1956/X sky130_fd_sc_hd__dlygate4sd3_1
X_07856_ hold2616/X _07865_/B _07855_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _07856_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1967 _08000_/X vssd1 vssd1 vccd1 vccd1 _15641_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1978 _18191_/Q vssd1 vssd1 vccd1 vccd1 hold1978/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1989 _14941_/X vssd1 vssd1 vccd1 vccd1 _18257_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07787_ _10603_/A vssd1 vssd1 vccd1 vccd1 _07787_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_190_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09526_ hold4484/X _10028_/B _09525_/X _15048_/A vssd1 vssd1 vccd1 vccd1 _09526_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_213_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09457_ _09463_/D _09478_/B _09457_/C vssd1 vssd1 vccd1 vccd1 _16312_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_78_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ hold2650/X _08442_/A2 _08407_/X _12738_/A vssd1 vssd1 vccd1 vccd1 _08408_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09388_ hold5937/A _09342_/B _09342_/Y _09387_/X _12412_/A vssd1 vssd1 vccd1 vccd1
+ _09388_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_108_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08339_ _08504_/A hold113/X vssd1 vssd1 vccd1 vccd1 hold114/A sky130_fd_sc_hd__or2_1
XFILLER_0_85_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11350_ hold5505/X _11732_/B _11349_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _11350_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10301_ hold1871/X hold3320/X _10649_/C vssd1 vssd1 vccd1 vccd1 _10302_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11281_ hold4961/X _11765_/B _11280_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _11281_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13020_ _09489_/B hold901/X vssd1 vssd1 vccd1 vccd1 hold902/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_24_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5250 _13387_/X vssd1 vssd1 vccd1 vccd1 _17582_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10232_ hold2351/X _16568_/Q _11213_/C vssd1 vssd1 vccd1 vccd1 _10233_/B sky130_fd_sc_hd__mux2_1
Xhold5261 _16979_/Q vssd1 vssd1 vccd1 vccd1 hold5261/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5272 _11488_/X vssd1 vssd1 vccd1 vccd1 _16986_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5283 _17674_/Q vssd1 vssd1 vccd1 vccd1 hold5283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5294 _11254_/X vssd1 vssd1 vccd1 vccd1 _16908_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4560 _13447_/X vssd1 vssd1 vccd1 vccd1 _17602_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4571 _16705_/Q vssd1 vssd1 vccd1 vccd1 hold4571/X sky130_fd_sc_hd__dlygate4sd3_1
X_10163_ hold2585/X hold4227/X _10646_/C vssd1 vssd1 vccd1 vccd1 _10164_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4582 _09742_/X vssd1 vssd1 vccd1 vccd1 _16404_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4593 _17361_/Q vssd1 vssd1 vccd1 vccd1 hold4593/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3870 _17228_/Q vssd1 vssd1 vccd1 vccd1 hold3870/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_234_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14971_ hold2185/X hold447/X _14970_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _14971_/X
+ sky130_fd_sc_hd__o211a_1
X_10094_ hold2238/X hold4330/X _11204_/C vssd1 vssd1 vccd1 vccd1 _10095_/B sky130_fd_sc_hd__mux2_1
Xhold3881 _09850_/X vssd1 vssd1 vccd1 vccd1 _16440_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3892 _17413_/Q vssd1 vssd1 vccd1 vccd1 hold3892/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16710_ _17913_/CLK _16710_/D vssd1 vssd1 vccd1 vccd1 _16710_/Q sky130_fd_sc_hd__dfxtp_1
X_13922_ _14477_/A hold2070/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13923_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_96_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17690_ _17690_/CLK _17690_/D vssd1 vssd1 vccd1 vccd1 _17690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16641_ _18218_/CLK _16641_/D vssd1 vssd1 vccd1 vccd1 _16641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13853_ _17738_/Q _13874_/B _13874_/C vssd1 vssd1 vccd1 vccd1 _13853_/X sky130_fd_sc_hd__and3_1
XFILLER_0_230_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_230_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12804_ _12804_/A _12804_/B vssd1 vssd1 vccd1 vccd1 _17444_/D sky130_fd_sc_hd__and2_1
X_16572_ _18162_/CLK _16572_/D vssd1 vssd1 vccd1 vccd1 _16572_/Q sky130_fd_sc_hd__dfxtp_1
X_10996_ hold5058/X _11186_/B _10995_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _10996_/X
+ sky130_fd_sc_hd__o211a_1
X_13784_ hold1438/X hold5412/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13785_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18311_ _18357_/CLK _18311_/D vssd1 vssd1 vccd1 vccd1 _18311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15523_ hold933/X _15559_/B vssd1 vssd1 vccd1 vccd1 _15523_/X sky130_fd_sc_hd__or2_1
XFILLER_0_214_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _12753_/A _12735_/B vssd1 vssd1 vccd1 vccd1 _17421_/D sky130_fd_sc_hd__and2_1
XFILLER_0_31_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ _18242_/CLK _18242_/D vssd1 vssd1 vccd1 vccd1 _18242_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _15482_/A _15454_/B vssd1 vssd1 vccd1 vccd1 _18421_/D sky130_fd_sc_hd__and2_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12873_/A _12666_/B vssd1 vssd1 vccd1 vccd1 _17398_/D sky130_fd_sc_hd__and2_1
XFILLER_0_182_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14405_ _15193_/A _14443_/B vssd1 vssd1 vccd1 vccd1 _14405_/X sky130_fd_sc_hd__or2_1
XFILLER_0_115_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11617_ hold5630/X _12305_/B _11616_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _17029_/D
+ sky130_fd_sc_hd__o211a_1
X_18173_ _18203_/CLK _18173_/D vssd1 vssd1 vccd1 vccd1 _18173_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_1_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_15385_ hold477/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15385_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12597_ _12597_/A _12597_/B vssd1 vssd1 vccd1 vccd1 _17375_/D sky130_fd_sc_hd__and2_1
XFILLER_0_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17124_ _17260_/CLK _17124_/D vssd1 vssd1 vccd1 vccd1 _17124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11548_ hold5315/X _11744_/B _11547_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _11548_/X
+ sky130_fd_sc_hd__o211a_1
X_14336_ _14443_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14336_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold508 input58/X vssd1 vssd1 vccd1 vccd1 hold508/X sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_334_wb_clk_i clkbuf_6_41_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17154_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14267_ hold2995/X _14268_/B _14266_/Y _14372_/A vssd1 vssd1 vccd1 vccd1 _14267_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold519 hold519/A vssd1 vssd1 vccd1 vccd1 hold519/X sky130_fd_sc_hd__dlygate4sd3_1
X_17055_ _18064_/CLK _17055_/D vssd1 vssd1 vccd1 vccd1 _17055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11479_ hold5004/X _11765_/B _11478_/X _14346_/A vssd1 vssd1 vccd1 vccd1 _11479_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16006_ _18413_/CLK _16006_/D vssd1 vssd1 vccd1 vccd1 _16006_/Q sky130_fd_sc_hd__dfxtp_1
X_13218_ _17578_/Q _17112_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13218_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_204_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14198_ _15163_/A _14198_/B vssd1 vssd1 vccd1 vccd1 _14198_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_221_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _13148_/X hold5996/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13149_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_196_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1208 _08444_/X vssd1 vssd1 vccd1 vccd1 _15852_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ _18020_/CLK _17957_/D vssd1 vssd1 vccd1 vccd1 _17957_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1219 _08326_/X vssd1 vssd1 vccd1 vccd1 _15796_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16908_ _17820_/CLK _16908_/D vssd1 vssd1 vccd1 vccd1 _16908_/Q sky130_fd_sc_hd__dfxtp_1
X_08690_ _12416_/A _08690_/B vssd1 vssd1 vccd1 vccd1 _15966_/D sky130_fd_sc_hd__and2_1
XFILLER_0_79_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17888_ _17888_/CLK _17888_/D vssd1 vssd1 vccd1 vccd1 _17888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16839_ _18042_/CLK _16839_/D vssd1 vssd1 vccd1 vccd1 _16839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_50_wb_clk_i clkbuf_6_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17853_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_180_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09311_ _15099_/A _09315_/B vssd1 vssd1 vccd1 vccd1 _09311_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09242_ _12786_/A _09242_/B vssd1 vssd1 vccd1 vccd1 _16232_/D sky130_fd_sc_hd__and2_1
XFILLER_0_185_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09173_ hold1626/X _09177_/A2 _09172_/X _12924_/A vssd1 vssd1 vccd1 vccd1 _09173_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_185_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08124_ _15529_/A hold2902/X hold108/X vssd1 vssd1 vccd1 vccd1 _08125_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_185_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08055_ hold2938/X _08097_/A2 _08054_/X _12103_/C1 vssd1 vssd1 vccd1 vccd1 _08055_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3100 _18252_/Q vssd1 vssd1 vccd1 vccd1 hold3100/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3111 _14466_/X vssd1 vssd1 vccd1 vccd1 _18030_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3122 _17400_/Q vssd1 vssd1 vccd1 vccd1 hold3122/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3133 _17397_/Q vssd1 vssd1 vccd1 vccd1 hold3133/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3144 _12656_/X vssd1 vssd1 vccd1 vccd1 _12657_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2410 _15570_/Q vssd1 vssd1 vccd1 vccd1 hold2410/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3155 _12677_/X vssd1 vssd1 vccd1 vccd1 _12678_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2421 _08269_/X vssd1 vssd1 vccd1 vccd1 _15769_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3166 _12731_/X vssd1 vssd1 vccd1 vccd1 _12732_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3177 _17423_/Q vssd1 vssd1 vccd1 vccd1 hold3177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2432 _07895_/X vssd1 vssd1 vccd1 vccd1 _15591_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08957_ hold163/X _16096_/Q _08997_/S vssd1 vssd1 vccd1 vccd1 hold164/A sky130_fd_sc_hd__mux2_1
Xhold3188 _16348_/Q vssd1 vssd1 vccd1 vccd1 _13254_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2443 _18066_/Q vssd1 vssd1 vccd1 vccd1 hold2443/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2454 _07985_/X vssd1 vssd1 vccd1 vccd1 _15635_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3199 _10039_/Y vssd1 vssd1 vccd1 vccd1 _16503_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1720 _15869_/Q vssd1 vssd1 vccd1 vccd1 hold1720/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2465 _09165_/X vssd1 vssd1 vccd1 vccd1 _16195_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1731 _14577_/X vssd1 vssd1 vccd1 vccd1 _18082_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07908_ _15531_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07908_/X sky130_fd_sc_hd__or2_1
Xhold2476 _15632_/Q vssd1 vssd1 vccd1 vccd1 hold2476/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08888_ hold673/X hold825/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold826/A sky130_fd_sc_hd__mux2_1
XFILLER_0_192_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1742 _17834_/Q vssd1 vssd1 vccd1 vccd1 hold1742/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2487 _17890_/Q vssd1 vssd1 vccd1 vccd1 hold2487/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2498 _14911_/X vssd1 vssd1 vccd1 vccd1 _18243_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1753 _07971_/X vssd1 vssd1 vccd1 vccd1 _15628_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1764 _18101_/Q vssd1 vssd1 vccd1 vccd1 hold1764/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1775 _15562_/Q vssd1 vssd1 vccd1 vccd1 hold1775/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07839_ _14457_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07839_/X sky130_fd_sc_hd__or2_1
Xhold1786 _14765_/X vssd1 vssd1 vccd1 vccd1 _18173_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1797 _18281_/Q vssd1 vssd1 vccd1 vccd1 hold1797/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10850_ hold1281/X hold4068/X _11732_/C vssd1 vssd1 vccd1 vccd1 _10851_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_196_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09509_ hold1779/X _13086_/A _10004_/C vssd1 vssd1 vccd1 vccd1 _09510_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10781_ hold2969/X hold5631/X _11654_/S vssd1 vssd1 vccd1 vccd1 _10782_/B sky130_fd_sc_hd__mux2_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12520_ hold1635/X hold4474/X _12925_/S vssd1 vssd1 vccd1 vccd1 _12520_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ hold131/X _12509_/A2 _12501_/A3 _12450_/X _12410_/A vssd1 vssd1 vccd1 vccd1
+ hold39/A sky130_fd_sc_hd__o311a_1
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11402_ hold1085/X hold4131/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11403_/B sky130_fd_sc_hd__mux2_1
X_15170_ hold1607/X _15165_/B _15169_/X _15042_/A vssd1 vssd1 vccd1 vccd1 _15170_/X
+ sky130_fd_sc_hd__o211a_1
X_12382_ _15244_/A hold727/X vssd1 vssd1 vccd1 vccd1 _17284_/D sky130_fd_sc_hd__and2_1
XFILLER_0_23_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_90 hold5959/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14121_ hold2530/X _14142_/B _14120_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14121_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11333_ hold3063/X hold4105/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11334_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14052_ _14732_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14052_/X sky130_fd_sc_hd__or2_1
X_11264_ hold957/X _16912_/Q _11741_/C vssd1 vssd1 vccd1 vccd1 _11265_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_219_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5080 _16464_/Q vssd1 vssd1 vccd1 vccd1 hold5080/X sky130_fd_sc_hd__dlygate4sd3_1
X_13003_ _14897_/A hold363/X vssd1 vssd1 vccd1 vccd1 _13003_/Y sky130_fd_sc_hd__nor2_2
X_10215_ _10563_/A _10215_/B vssd1 vssd1 vccd1 vccd1 _10215_/X sky130_fd_sc_hd__or2_1
Xhold5091 _12097_/X vssd1 vssd1 vccd1 vccd1 _17189_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_2_3_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_6530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11195_ _16889_/Q _11195_/B _11210_/C vssd1 vssd1 vccd1 vccd1 _11195_/X sky130_fd_sc_hd__and3_1
XTAP_6541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17811_ _17840_/CLK _17811_/D vssd1 vssd1 vccd1 vccd1 _17811_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4390 _16927_/Q vssd1 vssd1 vccd1 vccd1 hold4390/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_238_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10146_ _10530_/A _10146_/B vssd1 vssd1 vccd1 vccd1 _10146_/X sky130_fd_sc_hd__or2_1
XTAP_6574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17742_ _17742_/CLK _17742_/D vssd1 vssd1 vccd1 vccd1 _17742_/Q sky130_fd_sc_hd__dfxtp_1
X_14954_ hold484/A hold407/X vssd1 vssd1 vccd1 vccd1 hold240/A sky130_fd_sc_hd__or2_1
XTAP_5873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10077_ _10563_/A _10077_/B vssd1 vssd1 vccd1 vccd1 _10077_/X sky130_fd_sc_hd__or2_1
XTAP_5884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13905_ _13905_/A hold958/X vssd1 vssd1 vccd1 vccd1 _17760_/D sky130_fd_sc_hd__and2_1
X_17673_ _17705_/CLK _17673_/D vssd1 vssd1 vccd1 vccd1 _17673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14885_ hold6081/X hold332/X _14884_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 hold333/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16624_ _18214_/CLK _16624_/D vssd1 vssd1 vccd1 vccd1 _16624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13836_ hold4378/X _13773_/A _13835_/X vssd1 vssd1 vccd1 vccd1 _13836_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16555_ _18081_/CLK _16555_/D vssd1 vssd1 vccd1 vccd1 _16555_/Q sky130_fd_sc_hd__dfxtp_1
X_10979_ hold1342/X _16817_/Q _11654_/S vssd1 vssd1 vccd1 vccd1 _10980_/B sky130_fd_sc_hd__mux2_1
X_13767_ _13794_/A _13767_/B vssd1 vssd1 vccd1 vccd1 _13767_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15506_ _15506_/A _15506_/B vssd1 vssd1 vccd1 vccd1 _18432_/D sky130_fd_sc_hd__and2_1
X_12718_ _16237_/Q _17417_/Q _12766_/S vssd1 vssd1 vccd1 vccd1 _12718_/X sky130_fd_sc_hd__mux2_1
X_16486_ _18271_/CLK _16486_/D vssd1 vssd1 vccd1 vccd1 _16486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13698_ _13794_/A _13698_/B vssd1 vssd1 vccd1 vccd1 _13698_/X sky130_fd_sc_hd__or2_1
XFILLER_0_210_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18225_ _18225_/CLK _18225_/D vssd1 vssd1 vccd1 vccd1 _18225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15437_ _16096_/Q _09392_/B _09392_/C hold261/X vssd1 vssd1 vccd1 vccd1 _15437_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12649_ hold2745/X hold3146/X _12850_/S vssd1 vssd1 vccd1 vccd1 _12649_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18156_ _18156_/CLK _18156_/D vssd1 vssd1 vccd1 vccd1 _18156_/Q sky130_fd_sc_hd__dfxtp_1
X_15368_ hold102/X _15484_/A2 _09392_/D _17297_/Q vssd1 vssd1 vccd1 vccd1 _15368_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17107_ _17107_/CLK _17107_/D vssd1 vssd1 vccd1 vccd1 _17107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14319_ hold2151/X _14333_/A2 _14318_/X _14462_/C1 vssd1 vssd1 vccd1 vccd1 _14319_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold305 hold443/X vssd1 vssd1 vccd1 vccd1 hold444/A sky130_fd_sc_hd__buf_4
XFILLER_0_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18087_ _18087_/CLK _18087_/D vssd1 vssd1 vccd1 vccd1 _18087_/Q sky130_fd_sc_hd__dfxtp_1
Xhold316 hold316/A vssd1 vssd1 vccd1 vccd1 hold316/X sky130_fd_sc_hd__dlygate4sd3_1
X_15299_ hold263/X _15485_/A2 _15488_/A2 hold379/X _15298_/X vssd1 vssd1 vccd1 vccd1
+ _15302_/C sky130_fd_sc_hd__a221o_1
Xhold327 hold327/A vssd1 vssd1 vccd1 vccd1 hold327/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold338 hold338/A vssd1 vssd1 vccd1 vccd1 hold338/X sky130_fd_sc_hd__clkbuf_8
Xhold349 hold349/A vssd1 vssd1 vccd1 vccd1 hold349/X sky130_fd_sc_hd__dlygate4sd3_1
X_17038_ _17886_/CLK _17038_/D vssd1 vssd1 vccd1 vccd1 _17038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout807 _15070_/A vssd1 vssd1 vccd1 vccd1 _15050_/A sky130_fd_sc_hd__buf_4
X_09860_ hold3080/X hold4152/X _10040_/C vssd1 vssd1 vccd1 vccd1 _09861_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout818 _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14342_/A sky130_fd_sc_hd__buf_4
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout829 _14863_/C1 vssd1 vssd1 vccd1 vccd1 _14885_/C1 sky130_fd_sc_hd__clkbuf_4
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _12410_/A hold828/X vssd1 vssd1 vccd1 vccd1 _16024_/D sky130_fd_sc_hd__and2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ hold2695/X hold3601/X _10031_/C vssd1 vssd1 vccd1 vccd1 _09792_/B sky130_fd_sc_hd__mux2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 hold519/X vssd1 vssd1 vccd1 vccd1 input39/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1016 _08114_/X vssd1 vssd1 vccd1 vccd1 _08115_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ _12420_/A _08742_/B vssd1 vssd1 vccd1 vccd1 _15991_/D sky130_fd_sc_hd__and2_1
Xhold1027 _18029_/Q vssd1 vssd1 vccd1 vccd1 hold1027/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1038 _08300_/X vssd1 vssd1 vccd1 vccd1 _15783_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 _15781_/Q vssd1 vssd1 vccd1 vccd1 hold1049/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08673_ hold71/X _15958_/Q _08721_/S vssd1 vssd1 vccd1 vccd1 hold260/A sky130_fd_sc_hd__mux2_1
XFILLER_0_178_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_256_wb_clk_i clkbuf_6_58_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18056_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09225_ hold2809/X _09218_/B _09224_/X _12843_/A vssd1 vssd1 vccd1 vccd1 _09225_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09156_ _15539_/A _09156_/B vssd1 vssd1 vccd1 vccd1 _09156_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08107_ _08171_/A _08107_/B vssd1 vssd1 vccd1 vccd1 _15692_/D sky130_fd_sc_hd__and2_1
XFILLER_0_146_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_6_32_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_32_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_09087_ hold1386/X _09102_/B _09086_/X _14358_/A vssd1 vssd1 vccd1 vccd1 _09087_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08038_ hold1173/X _08033_/B _08037_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _08038_/X
+ sky130_fd_sc_hd__o211a_1
Xhold850 hold850/A vssd1 vssd1 vccd1 vccd1 hold850/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold861 hold861/A vssd1 vssd1 vccd1 vccd1 hold861/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold872 hold872/A vssd1 vssd1 vccd1 vccd1 hold872/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 hold883/A vssd1 vssd1 vccd1 vccd1 hold883/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 hold902/X vssd1 vssd1 vccd1 vccd1 hold894/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10000_ _11158_/A _10000_/B vssd1 vssd1 vccd1 vccd1 _16490_/D sky130_fd_sc_hd__nor2_1
XTAP_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09989_ _16487_/Q _10004_/B _10004_/C vssd1 vssd1 vccd1 vccd1 _09989_/X sky130_fd_sc_hd__and3_1
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2240 _14571_/X vssd1 vssd1 vccd1 vccd1 _18080_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2251 hold919/X vssd1 vssd1 vccd1 vccd1 input4/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2262 _14861_/X vssd1 vssd1 vccd1 vccd1 _18219_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2273 _12617_/X vssd1 vssd1 vccd1 vccd1 _12618_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2284 _16232_/Q vssd1 vssd1 vccd1 vccd1 hold2284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2295 _18124_/Q vssd1 vssd1 vccd1 vccd1 hold2295/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1550 _17822_/Q vssd1 vssd1 vccd1 vccd1 hold1550/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1561 _14159_/X vssd1 vssd1 vccd1 vccd1 _17883_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1572 _16215_/Q vssd1 vssd1 vccd1 vccd1 hold1572/X sky130_fd_sc_hd__dlygate4sd3_1
X_11951_ hold3047/X hold5462/X _12335_/C vssd1 vssd1 vccd1 vccd1 _11952_/B sky130_fd_sc_hd__mux2_1
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1583 _17968_/Q vssd1 vssd1 vccd1 vccd1 hold1583/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1594 _15829_/Q vssd1 vssd1 vccd1 vccd1 hold1594/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10902_ _11121_/A _10902_/B vssd1 vssd1 vccd1 vccd1 _10902_/X sky130_fd_sc_hd__or2_1
X_14670_ _15225_/A _14672_/B vssd1 vssd1 vccd1 vccd1 _14670_/X sky130_fd_sc_hd__or2_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11882_ _15710_/Q hold5717/X _12362_/C vssd1 vssd1 vccd1 vccd1 _11883_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10833_ _11121_/A _10833_/B vssd1 vssd1 vccd1 vccd1 _10833_/X sky130_fd_sc_hd__or2_1
X_13621_ hold4756/X _13811_/B _13620_/X _12822_/A vssd1 vssd1 vccd1 vccd1 _13621_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16340_ _18387_/CLK _16340_/D vssd1 vssd1 vccd1 vccd1 _16340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10764_ _11049_/A _10764_/B vssd1 vssd1 vccd1 vccd1 _10764_/X sky130_fd_sc_hd__or2_1
X_13552_ hold5432/X _13856_/B _13551_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13552_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12503_ hold8/X _12445_/A _12445_/B _12502_/X _09057_/A vssd1 vssd1 vccd1 vccd1 hold9/A
+ sky130_fd_sc_hd__o311a_1
X_13483_ hold5211/X _12356_/B _13482_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _13483_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16271_ _18013_/CLK _16271_/D vssd1 vssd1 vccd1 vccd1 _16271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10695_ _11658_/A _10695_/B vssd1 vssd1 vccd1 vccd1 _10695_/X sky130_fd_sc_hd__or2_1
X_18010_ _18010_/CLK _18010_/D vssd1 vssd1 vccd1 vccd1 _18010_/Q sky130_fd_sc_hd__dfxtp_1
X_12434_ _15274_/A _12434_/B vssd1 vssd1 vccd1 vccd1 _17310_/D sky130_fd_sc_hd__and2_1
X_15222_ hold2306/X _15221_/B _15221_/Y _15226_/C1 vssd1 vssd1 vccd1 vccd1 _15222_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15153_ _15207_/A _15157_/B vssd1 vssd1 vccd1 vccd1 _15153_/X sky130_fd_sc_hd__or2_1
XFILLER_0_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12365_ _17279_/Q _12365_/B _12371_/C vssd1 vssd1 vccd1 vccd1 _12365_/X sky130_fd_sc_hd__and3_1
XFILLER_0_129_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11316_ _12240_/A _11316_/B vssd1 vssd1 vccd1 vccd1 _11316_/X sky130_fd_sc_hd__or2_1
X_14104_ _14443_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14104_/X sky130_fd_sc_hd__or2_1
X_15084_ hold2345/X hold341/X _15083_/X _15212_/C1 vssd1 vssd1 vccd1 vccd1 _15084_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12296_ _17256_/Q _13811_/B _13811_/C vssd1 vssd1 vccd1 vccd1 _12296_/X sky130_fd_sc_hd__and3_1
XFILLER_0_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14035_ hold2779/X _14038_/B _14034_/Y _14193_/C1 vssd1 vssd1 vccd1 vccd1 _14035_/X
+ sky130_fd_sc_hd__o211a_1
X_11247_ _11631_/A _11247_/B vssd1 vssd1 vccd1 vccd1 _11247_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11178_ hold4341/X _11109_/A _11177_/X vssd1 vssd1 vccd1 vccd1 _11178_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10129_ hold3811/X _10631_/B _10128_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10129_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15986_ _16125_/CLK _15986_/D vssd1 vssd1 vccd1 vccd1 hold757/A sky130_fd_sc_hd__dfxtp_1
XTAP_5670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17725_ _17725_/CLK _17725_/D vssd1 vssd1 vccd1 vccd1 _17725_/Q sky130_fd_sc_hd__dfxtp_1
X_14937_ hold1315/X _14952_/B _14936_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _14937_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17656_ _17726_/CLK _17656_/D vssd1 vssd1 vccd1 vccd1 _17656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14868_ _15099_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14868_/X sky130_fd_sc_hd__or2_1
XFILLER_0_187_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_230_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16607_ _18197_/CLK _16607_/D vssd1 vssd1 vccd1 vccd1 _16607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13819_ _13819_/A _13819_/B vssd1 vssd1 vccd1 vccd1 _13819_/Y sky130_fd_sc_hd__nor2_1
X_17587_ _17747_/CLK _17587_/D vssd1 vssd1 vccd1 vccd1 _17587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14799_ hold2522/X _14826_/B _14798_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14799_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16538_ _18180_/CLK _16538_/D vssd1 vssd1 vccd1 vccd1 _16538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16469_ _18382_/CLK _16469_/D vssd1 vssd1 vccd1 vccd1 _16469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09010_ hold147/X hold665/X _09060_/S vssd1 vssd1 vccd1 vccd1 _09011_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_128_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18208_ _18208_/CLK _18208_/D vssd1 vssd1 vccd1 vccd1 _18208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18139_ _18262_/CLK _18139_/D vssd1 vssd1 vccd1 vccd1 _18139_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5805 _17202_/Q vssd1 vssd1 vccd1 vccd1 hold5805/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5816 _13327_/X vssd1 vssd1 vccd1 vccd1 _17562_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold102 hold102/A vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5827 _16494_/Q vssd1 vssd1 vccd1 vccd1 hold5827/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5838 _09538_/X vssd1 vssd1 vccd1 vccd1 _16336_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 hold113/A vssd1 vssd1 vccd1 vccd1 hold113/X sky130_fd_sc_hd__clkbuf_4
Xhold5849 hold6010/X vssd1 vssd1 vccd1 vccd1 _13273_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 hold124/A vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold135 hold135/A vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 hold392/X vssd1 vssd1 vccd1 vccd1 hold393/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 hold681/X vssd1 vssd1 vccd1 vccd1 hold682/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 input9/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__buf_1
Xhold179 input11/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__buf_1
X_09912_ _09912_/A _09912_/B vssd1 vssd1 vccd1 vccd1 _09912_/X sky130_fd_sc_hd__or2_1
Xfanout604 _15484_/B1 vssd1 vssd1 vccd1 vccd1 _09386_/D sky130_fd_sc_hd__buf_8
Xfanout615 _09358_/Y vssd1 vssd1 vccd1 vccd1 _09392_/B sky130_fd_sc_hd__clkbuf_8
Xfanout626 _09339_/Y vssd1 vssd1 vccd1 vccd1 _15490_/A1 sky130_fd_sc_hd__buf_8
X_09843_ _09981_/A _09843_/B vssd1 vssd1 vccd1 vccd1 _09843_/X sky130_fd_sc_hd__or2_1
Xfanout637 _12199_/C1 vssd1 vssd1 vccd1 vccd1 _12798_/A sky130_fd_sc_hd__buf_2
Xfanout648 fanout739/X vssd1 vssd1 vccd1 vccd1 _12199_/C1 sky130_fd_sc_hd__buf_4
Xfanout659 _12588_/A vssd1 vssd1 vccd1 vccd1 _12894_/A sky130_fd_sc_hd__buf_4
XFILLER_0_77_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _09954_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09774_/X sky130_fd_sc_hd__or2_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ hold320/X hold389/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08726_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_197_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _12438_/A hold103/X vssd1 vssd1 vccd1 vccd1 _15950_/D sky130_fd_sc_hd__and2_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_437_wb_clk_i clkbuf_6_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17426_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _15284_/A hold499/X vssd1 vssd1 vccd1 vccd1 _15917_/D sky130_fd_sc_hd__and2_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09208_ _15537_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09208_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10480_ hold5144/X _11204_/B _10479_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _10480_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09139_ hold2657/X _09177_/A2 _09138_/X _12888_/A vssd1 vssd1 vccd1 vccd1 _09139_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12150_ _12273_/A _12150_/B vssd1 vssd1 vccd1 vccd1 _12150_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11101_ hold4113/X _11195_/B _11100_/X _14528_/C1 vssd1 vssd1 vccd1 vccd1 _11101_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12081_ _13407_/A _12081_/B vssd1 vssd1 vccd1 vccd1 _12081_/X sky130_fd_sc_hd__or2_1
Xhold680 hold680/A vssd1 vssd1 vccd1 vccd1 hold680/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold691 hold691/A vssd1 vssd1 vccd1 vccd1 hold691/X sky130_fd_sc_hd__buf_4
XFILLER_0_198_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11032_ hold3958/X _11789_/B _11031_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _11032_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_217_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ _17731_/CLK _15840_/D vssd1 vssd1 vccd1 vccd1 _15840_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2070 _17769_/Q vssd1 vssd1 vccd1 vccd1 hold2070/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2081 _18291_/Q vssd1 vssd1 vccd1 vccd1 hold2081/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2092 _16190_/Q vssd1 vssd1 vccd1 vccd1 hold2092/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _17690_/CLK _15771_/D vssd1 vssd1 vccd1 vccd1 _15771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12983_ hold4479/X _12982_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12984_/B sky130_fd_sc_hd__mux2_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ _18400_/CLK _17510_/D vssd1 vssd1 vccd1 vccd1 _17510_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1380 _15866_/Q vssd1 vssd1 vccd1 vccd1 hold1380/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14722_ _15169_/A _14730_/B vssd1 vssd1 vccd1 vccd1 _14722_/X sky130_fd_sc_hd__or2_1
Xhold1391 _13889_/Y vssd1 vssd1 vccd1 vccd1 hold1391/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _12285_/A _11934_/B vssd1 vssd1 vccd1 vccd1 _11934_/X sky130_fd_sc_hd__or2_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_178_wb_clk_i clkbuf_6_49_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18357_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_131_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _17445_/CLK _17441_/D vssd1 vssd1 vccd1 vccd1 _17441_/Q sky130_fd_sc_hd__dfxtp_1
X_14653_ hold2918/X _14664_/B _14652_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14653_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11865_ _12273_/A _11865_/B vssd1 vssd1 vccd1 vccd1 _11865_/X sky130_fd_sc_hd__or2_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_107_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18413_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13604_ hold2857/X _17655_/Q _13817_/C vssd1 vssd1 vccd1 vccd1 _13605_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10816_ hold5549/X _11213_/B _10815_/X _14342_/A vssd1 vssd1 vccd1 vccd1 _10816_/X
+ sky130_fd_sc_hd__o211a_1
X_17372_ _17881_/CLK _17372_/D vssd1 vssd1 vccd1 vccd1 _17372_/Q sky130_fd_sc_hd__dfxtp_1
X_14584_ _15193_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14584_/X sky130_fd_sc_hd__or2_1
X_11796_ hold4411/X _12240_/A _11795_/X vssd1 vssd1 vccd1 vccd1 _11796_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16323_ _16323_/CLK _16323_/D vssd1 vssd1 vccd1 vccd1 _16323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13535_ hold1263/X _17632_/Q _13862_/C vssd1 vssd1 vccd1 vccd1 _13536_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_171_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10747_ hold5018/X _11222_/B _10746_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _10747_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16254_ _17517_/CLK _16254_/D vssd1 vssd1 vccd1 vccd1 _16254_/Q sky130_fd_sc_hd__dfxtp_1
X_10678_ hold4905/X _11162_/B _10677_/X _15176_/C1 vssd1 vssd1 vccd1 vccd1 _10678_/X
+ sky130_fd_sc_hd__o211a_1
X_13466_ hold1330/X hold5472/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13467_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15205_ _15205_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15205_/X sky130_fd_sc_hd__or2_1
X_12417_ hold245/X hold489/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12418_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_112_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16185_ _17471_/CLK _16185_/D vssd1 vssd1 vccd1 vccd1 _16185_/Q sky130_fd_sc_hd__dfxtp_1
X_13397_ hold1442/X hold3547/X _13877_/C vssd1 vssd1 vccd1 vccd1 _13398_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15136_ hold3184/X _15167_/B _15135_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _15136_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12348_ hold5705/X _12255_/A _12347_/X vssd1 vssd1 vccd1 vccd1 _12348_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15067_ _15229_/A hold2751/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15068_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12279_ _13749_/A _12279_/B vssd1 vssd1 vccd1 vccd1 _12279_/X sky130_fd_sc_hd__or2_1
XFILLER_0_208_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14018_ _15525_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14018_/X sky130_fd_sc_hd__or2_1
XTAP_6190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_235_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15969_ _17284_/CLK _15969_/D vssd1 vssd1 vccd1 vccd1 hold558/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08510_ hold2320/X _08503_/Y _08509_/X _13417_/C1 vssd1 vssd1 vccd1 vccd1 _08510_/X
+ sky130_fd_sc_hd__o211a_1
X_17708_ _17734_/CLK _17708_/D vssd1 vssd1 vccd1 vccd1 _17708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09490_ hold935/X _09490_/B hold937/X vssd1 vssd1 vccd1 vccd1 _13055_/C sky130_fd_sc_hd__and3_4
XFILLER_0_72_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08441_ _14960_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08441_/X sky130_fd_sc_hd__or2_1
X_17639_ _17639_/CLK _17639_/D vssd1 vssd1 vccd1 vccd1 _17639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08372_ hold384/A _15818_/Q hold115/X vssd1 vssd1 vccd1 vccd1 hold230/A sky130_fd_sc_hd__mux2_1
XFILLER_0_59_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5602 _11998_/X vssd1 vssd1 vccd1 vccd1 _17156_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5613 _11923_/X vssd1 vssd1 vccd1 vccd1 _17131_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5624 _16934_/Q vssd1 vssd1 vccd1 vccd1 hold5624/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5635 _16964_/Q vssd1 vssd1 vccd1 vccd1 hold5635/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5646 _11275_/X vssd1 vssd1 vccd1 vccd1 _16915_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4901 _16939_/Q vssd1 vssd1 vccd1 vccd1 hold4901/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4912 _10900_/X vssd1 vssd1 vccd1 vccd1 _16790_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5657 _17073_/Q vssd1 vssd1 vccd1 vccd1 hold5657/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4923 _17093_/Q vssd1 vssd1 vccd1 vccd1 hold4923/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5668 _11659_/X vssd1 vssd1 vccd1 vccd1 _17043_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4934 _11311_/X vssd1 vssd1 vccd1 vccd1 _16927_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5679 _17049_/Q vssd1 vssd1 vccd1 vccd1 hold5679/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4945 _16787_/Q vssd1 vssd1 vccd1 vccd1 hold4945/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4956 _10918_/X vssd1 vssd1 vccd1 vccd1 _16796_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4967 _11899_/X vssd1 vssd1 vccd1 vccd1 _17123_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4978 _17731_/Q vssd1 vssd1 vccd1 vccd1 hold4978/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout401 _14443_/B vssd1 vssd1 vccd1 vccd1 _14445_/B sky130_fd_sc_hd__buf_6
Xfanout412 _14204_/B vssd1 vssd1 vccd1 vccd1 _14214_/B sky130_fd_sc_hd__buf_6
Xhold4989 _17013_/Q vssd1 vssd1 vccd1 vccd1 hold4989/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout423 _14000_/Y vssd1 vssd1 vccd1 vccd1 _14040_/B sky130_fd_sc_hd__buf_8
Xfanout434 _13052_/X vssd1 vssd1 vccd1 vccd1 _13311_/A1 sky130_fd_sc_hd__buf_12
Xfanout445 _12227_/S vssd1 vssd1 vccd1 vccd1 _13481_/S sky130_fd_sc_hd__buf_6
Xfanout456 _11168_/C vssd1 vssd1 vccd1 vccd1 _11738_/C sky130_fd_sc_hd__clkbuf_8
X_09826_ hold5080/X _11171_/B _09825_/X _15176_/C1 vssd1 vssd1 vccd1 vccd1 _09826_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout467 _13877_/C vssd1 vssd1 vccd1 vccd1 _13874_/C sky130_fd_sc_hd__clkbuf_4
Xfanout478 fanout485/X vssd1 vssd1 vccd1 vccd1 _11210_/C sky130_fd_sc_hd__buf_4
Xfanout489 _11201_/C vssd1 vssd1 vccd1 vccd1 _11171_/C sky130_fd_sc_hd__buf_6
XFILLER_0_225_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09757_ hold4741/X _10031_/B _09756_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09757_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_216_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_wb_clk_i clkbuf_6_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18453_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_240_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _15344_/A _08708_/B vssd1 vssd1 vccd1 vccd1 _15975_/D sky130_fd_sc_hd__and2_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ hold3982/X _11204_/B _09687_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _09688_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_271_wb_clk_i clkbuf_6_57_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18228_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ hold5/X hold165/X _08657_/S vssd1 vssd1 vccd1 vccd1 _08640_/B sky130_fd_sc_hd__mux2_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_200_wb_clk_i clkbuf_6_53_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18352_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_83_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11650_ hold5622/X _11744_/B _11649_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _11650_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10601_ _10601_/A _10601_/B _10601_/C vssd1 vssd1 vccd1 vccd1 _10601_/X sky130_fd_sc_hd__and3_1
XFILLER_0_166_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11581_ hold5679/X _11771_/B _11580_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _11581_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10532_ hold2207/X _16668_/Q _11213_/C vssd1 vssd1 vccd1 vccd1 _10533_/B sky130_fd_sc_hd__mux2_1
X_13320_ _13800_/A _13320_/B vssd1 vssd1 vccd1 vccd1 _13320_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10463_ hold2528/X _16645_/Q _10475_/S vssd1 vssd1 vccd1 vccd1 _10464_/B sky130_fd_sc_hd__mux2_1
X_13251_ _13250_/X _16924_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13251_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_161_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12202_ hold4859/X _13811_/B _12201_/X _12822_/A vssd1 vssd1 vccd1 vccd1 _12202_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13182_ _13182_/A _13294_/B vssd1 vssd1 vccd1 vccd1 _13182_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10394_ hold2161/X hold3556/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10395_/B sky130_fd_sc_hd__mux2_1
X_12133_ hold5795/X _12362_/B _12132_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _12133_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17990_ _18347_/CLK _17990_/D vssd1 vssd1 vccd1 vccd1 _17990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12064_ hold5775/X _12350_/B _12063_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _12064_/X
+ sky130_fd_sc_hd__o211a_1
X_16941_ _17853_/CLK _16941_/D vssd1 vssd1 vccd1 vccd1 _16941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_236_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11015_ hold1487/X hold5154/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11016_/B sky130_fd_sc_hd__mux2_1
X_16872_ _18046_/CLK _16872_/D vssd1 vssd1 vccd1 vccd1 _16872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15823_ _17702_/CLK _15823_/D vssd1 vssd1 vccd1 vccd1 _15823_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_359_wb_clk_i clkbuf_6_41_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17242_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_205_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _17737_/CLK _15754_/D vssd1 vssd1 vccd1 vccd1 _15754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12966_ _14362_/A _12966_/B vssd1 vssd1 vccd1 vccd1 _17498_/D sky130_fd_sc_hd__and2_1
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ hold2035/X _14720_/B _14704_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _14705_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11917_ hold5673/X _12299_/B _11916_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _11917_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15685_ _17268_/CLK _15685_/D vssd1 vssd1 vccd1 vccd1 _15685_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _12906_/A _12897_/B vssd1 vssd1 vccd1 vccd1 _17475_/D sky130_fd_sc_hd__and2_1
XFILLER_0_142_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17424_ _17426_/CLK _17424_/D vssd1 vssd1 vccd1 vccd1 _17424_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _15191_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14636_/X sky130_fd_sc_hd__or2_1
XFILLER_0_158_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11848_ hold4491/X _12332_/B _11847_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _11848_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _17517_/CLK _17355_/D vssd1 vssd1 vccd1 vccd1 _17355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14567_ _15191_/A _14557_/Y hold2232/X _15218_/C1 vssd1 vssd1 vccd1 vccd1 _14567_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11779_ _13864_/A _11779_/B vssd1 vssd1 vccd1 vccd1 _11779_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_83_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16306_ _16315_/CLK _16306_/D vssd1 vssd1 vccd1 vccd1 _16306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13518_ _13719_/A _13518_/B vssd1 vssd1 vccd1 vccd1 _13518_/X sky130_fd_sc_hd__or2_1
X_17286_ _18409_/CLK _17286_/D vssd1 vssd1 vccd1 vccd1 hold390/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14498_ hold2127/X _14487_/B _14497_/X _14354_/A vssd1 vssd1 vccd1 vccd1 _14498_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16237_ _17429_/CLK hold953/X vssd1 vssd1 vccd1 vccd1 _16237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13449_ _13737_/A _13449_/B vssd1 vssd1 vccd1 vccd1 _13449_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_75_wb_clk_i clkbuf_6_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17978_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_152_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4208 _15472_/X vssd1 vssd1 vccd1 vccd1 _15473_/B sky130_fd_sc_hd__dlygate4sd3_1
X_16168_ _17493_/CLK _16168_/D vssd1 vssd1 vccd1 vccd1 _16168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4219 _16012_/Q vssd1 vssd1 vccd1 vccd1 _15425_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15119_ _15227_/A _15119_/B vssd1 vssd1 vccd1 vccd1 _15119_/X sky130_fd_sc_hd__or2_1
Xhold3507 _12373_/Y vssd1 vssd1 vccd1 vccd1 _17281_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_227_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08990_ _15374_/A hold83/X vssd1 vssd1 vccd1 vccd1 _16112_/D sky130_fd_sc_hd__and2_1
X_16099_ _17303_/CLK _16099_/D vssd1 vssd1 vccd1 vccd1 hold688/A sky130_fd_sc_hd__dfxtp_1
Xhold3518 _11199_/Y vssd1 vssd1 vccd1 vccd1 _11200_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3529 _13849_/Y vssd1 vssd1 vccd1 vccd1 _17736_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2806 _14416_/X vssd1 vssd1 vccd1 vccd1 _18006_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07941_ hold1336/X _07991_/A2 _07940_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _07941_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_220_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2817 _17868_/Q vssd1 vssd1 vccd1 vccd1 hold2817/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2828 _15625_/Q vssd1 vssd1 vccd1 vccd1 hold2828/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2839 _14959_/X vssd1 vssd1 vccd1 vccd1 _18266_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07872_ hold1554/X _07869_/B _07871_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _07872_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09611_ _18274_/Q _16361_/Q _10004_/C vssd1 vssd1 vccd1 vccd1 _09612_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09542_ hold1960/X _13174_/A _10022_/C vssd1 vssd1 vccd1 vccd1 _09543_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_218_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_1310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09473_ _09477_/C _09478_/B _09473_/C vssd1 vssd1 vccd1 vccd1 _16318_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_231_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08424_ hold1704/X _08433_/B _08423_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08424_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08355_ _12750_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _15809_/D sky130_fd_sc_hd__and2_1
XFILLER_0_18_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08286_ hold1770/X _08336_/A2 _08285_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08286_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6100 la_data_in[20] vssd1 vssd1 vccd1 vccd1 hold481/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold6111 _17522_/Q vssd1 vssd1 vccd1 vccd1 hold6111/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6122 _16319_/Q vssd1 vssd1 vccd1 vccd1 hold6122/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6133 _16306_/Q vssd1 vssd1 vccd1 vccd1 hold6133/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5410 _17022_/Q vssd1 vssd1 vccd1 vccd1 hold5410/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5421 _10426_/X vssd1 vssd1 vccd1 vccd1 _16632_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5432 _17669_/Q vssd1 vssd1 vccd1 vccd1 hold5432/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5443 _12211_/X vssd1 vssd1 vccd1 vccd1 _17227_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5454 _17089_/Q vssd1 vssd1 vccd1 vccd1 hold5454/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4720 _16457_/Q vssd1 vssd1 vccd1 vccd1 hold4720/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5465 _13786_/X vssd1 vssd1 vccd1 vccd1 _17715_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4731 _17665_/Q vssd1 vssd1 vccd1 vccd1 hold4731/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5476 _17675_/Q vssd1 vssd1 vccd1 vccd1 hold5476/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4742 _09757_/X vssd1 vssd1 vccd1 vccd1 _16409_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5487 _13753_/X vssd1 vssd1 vccd1 vccd1 _17704_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4753 _11755_/Y vssd1 vssd1 vccd1 vccd1 _17075_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5498 _17706_/Q vssd1 vssd1 vccd1 vccd1 hold5498/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4764 _17699_/Q vssd1 vssd1 vccd1 vccd1 hold4764/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4775 _16424_/Q vssd1 vssd1 vccd1 vccd1 hold4775/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4786 _13414_/X vssd1 vssd1 vccd1 vccd1 _17591_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout220 _10025_/B vssd1 vssd1 vccd1 vccd1 _10031_/B sky130_fd_sc_hd__clkbuf_8
Xhold4797 _17224_/Q vssd1 vssd1 vccd1 vccd1 hold4797/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout231 _10604_/B vssd1 vssd1 vccd1 vccd1 _10628_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout242 _10589_/B vssd1 vssd1 vccd1 vccd1 _10649_/B sky130_fd_sc_hd__buf_4
Xfanout253 fanout299/X vssd1 vssd1 vccd1 vccd1 _13800_/A sky130_fd_sc_hd__buf_4
XFILLER_0_227_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout264 _11043_/A vssd1 vssd1 vccd1 vccd1 _11637_/A sky130_fd_sc_hd__buf_4
XFILLER_0_227_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout275 _12159_/A vssd1 vssd1 vccd1 vccd1 _13581_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_236_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout286 _11667_/A vssd1 vssd1 vccd1 vccd1 _12234_/A sky130_fd_sc_hd__buf_4
X_09809_ hold2534/X _16427_/Q _10025_/C vssd1 vssd1 vccd1 vccd1 _09810_/B sky130_fd_sc_hd__mux2_1
Xfanout297 _11127_/A vssd1 vssd1 vccd1 vccd1 _11124_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_452_wb_clk_i clkbuf_6_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17722_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_226_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12820_ hold2754/X hold3127/X _12871_/S vssd1 vssd1 vccd1 vccd1 _12820_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ hold1264/X hold3394/X _12766_/S vssd1 vssd1 vccd1 vccd1 _12751_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ hold1285/X hold3866/X _12173_/S vssd1 vssd1 vccd1 vccd1 _11703_/B sky130_fd_sc_hd__mux2_1
X_15470_ hold401/X _09392_/C _15467_/X vssd1 vssd1 vccd1 vccd1 _15471_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_167_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ hold1937/X hold3372/X _12844_/S vssd1 vssd1 vccd1 vccd1 _12682_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_166_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14421_ _15535_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14421_/X sky130_fd_sc_hd__or2_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ hold1560/X hold5002/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11634_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17140_ _17270_/CLK _17140_/D vssd1 vssd1 vccd1 vccd1 _17140_/Q sky130_fd_sc_hd__dfxtp_1
X_14352_ _14352_/A hold418/X vssd1 vssd1 vccd1 vccd1 hold419/A sky130_fd_sc_hd__and2_1
XFILLER_0_37_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11564_ hold2117/X _17012_/Q _11660_/S vssd1 vssd1 vccd1 vccd1 _11565_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13303_ _13052_/X _13301_/X _13302_/X _13049_/Y vssd1 vssd1 vccd1 vccd1 _13303_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_208_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10515_ _10515_/A _10515_/B vssd1 vssd1 vccd1 vccd1 _10515_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17071_ _17887_/CLK _17071_/D vssd1 vssd1 vccd1 vccd1 _17071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14283_ hold1420/X _14272_/B _14282_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _14283_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11495_ hold2577/X _16989_/Q _12329_/C vssd1 vssd1 vccd1 vccd1 _11496_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16022_ _16090_/CLK _16022_/D vssd1 vssd1 vccd1 vccd1 hold794/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10446_ _10536_/A _10446_/B vssd1 vssd1 vccd1 vccd1 _10446_/X sky130_fd_sc_hd__or2_1
X_13234_ _17580_/Q _17114_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13234_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13165_ _13164_/X hold3499/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13165_/X sky130_fd_sc_hd__mux2_1
X_10377_ _10476_/A _10377_/B vssd1 vssd1 vccd1 vccd1 _10377_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12116_ hold2476/X _17196_/Q _13721_/S vssd1 vssd1 vccd1 vccd1 _12117_/B sky130_fd_sc_hd__mux2_1
X_13096_ _13089_/X _13095_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17530_/D sky130_fd_sc_hd__o21a_1
X_17973_ _17973_/CLK _17973_/D vssd1 vssd1 vccd1 vccd1 _17973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12047_ hold2775/X hold5575/X _12335_/C vssd1 vssd1 vccd1 vccd1 _12048_/B sky130_fd_sc_hd__mux2_1
X_16924_ _17838_/CLK _16924_/D vssd1 vssd1 vccd1 vccd1 _16924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_193_wb_clk_i clkbuf_6_52_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18250_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_40_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16855_ _18056_/CLK _16855_/D vssd1 vssd1 vccd1 vccd1 _16855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_122_wb_clk_i clkbuf_6_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17324_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15806_ _17703_/CLK _15806_/D vssd1 vssd1 vccd1 vccd1 _15806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16786_ _18021_/CLK _16786_/D vssd1 vssd1 vccd1 vccd1 _16786_/Q sky130_fd_sc_hd__dfxtp_1
X_13998_ _14732_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13998_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15737_ _17748_/CLK _15737_/D vssd1 vssd1 vccd1 vccd1 _15737_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12949_ hold3070/X hold3759/X _12985_/S vssd1 vssd1 vccd1 vccd1 _12949_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18456_ _18457_/CLK _18456_/D vssd1 vssd1 vccd1 vccd1 _18456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15668_ _17628_/CLK _15668_/D vssd1 vssd1 vccd1 vccd1 _15668_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17407_ _18458_/CLK _17407_/D vssd1 vssd1 vccd1 vccd1 _17407_/Q sky130_fd_sc_hd__dfxtp_1
X_14619_ hold2585/X _14612_/B _14618_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14619_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18387_ _18387_/CLK _18387_/D vssd1 vssd1 vccd1 vccd1 _18387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15599_ _17247_/CLK _15599_/D vssd1 vssd1 vccd1 vccd1 _15599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08140_ hold220/X _15709_/Q hold108/X vssd1 vssd1 vccd1 vccd1 hold356/A sky130_fd_sc_hd__mux2_1
X_17338_ _17338_/CLK hold54/X vssd1 vssd1 vccd1 vccd1 _17338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08071_ hold2655/X _08097_/A2 _08070_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _08071_/X
+ sky130_fd_sc_hd__o211a_1
X_17269_ _17269_/CLK _17269_/D vssd1 vssd1 vccd1 vccd1 _17269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4005 _17279_/Q vssd1 vssd1 vccd1 vccd1 hold4005/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4016 _16754_/Q vssd1 vssd1 vccd1 vccd1 hold4016/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4027 _11929_/X vssd1 vssd1 vccd1 vccd1 _17133_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4038 _12151_/X vssd1 vssd1 vccd1 vccd1 _17207_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3304 _10477_/X vssd1 vssd1 vccd1 vccd1 _16649_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4049 _13675_/X vssd1 vssd1 vccd1 vccd1 _17678_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3315 _12923_/X vssd1 vssd1 vccd1 vccd1 _12924_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3326 _16611_/Q vssd1 vssd1 vccd1 vccd1 hold3326/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3337 _16655_/Q vssd1 vssd1 vccd1 vccd1 hold3337/X sky130_fd_sc_hd__dlygate4sd3_1
X_08973_ hold215/X _16104_/Q _08991_/S vssd1 vssd1 vccd1 vccd1 hold216/A sky130_fd_sc_hd__mux2_1
Xhold2603 _17904_/Q vssd1 vssd1 vccd1 vccd1 hold2603/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3348 _10555_/X vssd1 vssd1 vccd1 vccd1 _16675_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2614 _14434_/X vssd1 vssd1 vccd1 vccd1 _18015_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3359 _17391_/Q vssd1 vssd1 vccd1 vccd1 hold3359/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__buf_4
Xhold2625 _16204_/Q vssd1 vssd1 vccd1 vccd1 hold2625/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ _15547_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _07924_/Y sky130_fd_sc_hd__nand2_1
Xhold2636 _14243_/X vssd1 vssd1 vccd1 vccd1 _17922_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1902 _14476_/X vssd1 vssd1 vccd1 vccd1 _18035_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2647 _14440_/X vssd1 vssd1 vccd1 vccd1 _18018_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1913 _18239_/Q vssd1 vssd1 vccd1 vccd1 hold1913/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2658 _09139_/X vssd1 vssd1 vccd1 vccd1 _16182_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1924 _09221_/X vssd1 vssd1 vccd1 vccd1 _16222_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2669 _15792_/Q vssd1 vssd1 vccd1 vccd1 hold2669/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1935 _15752_/Q vssd1 vssd1 vccd1 vccd1 hold1935/X sky130_fd_sc_hd__dlygate4sd3_1
X_07855_ _15533_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07855_/X sky130_fd_sc_hd__or2_1
Xhold1946 _07927_/X vssd1 vssd1 vccd1 vccd1 _15607_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1957 _14492_/X vssd1 vssd1 vccd1 vccd1 _18043_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1968 _18374_/Q vssd1 vssd1 vccd1 vccd1 hold1968/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1979 _14803_/X vssd1 vssd1 vccd1 vccd1 _18191_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07786_ _07786_/A vssd1 vssd1 vccd1 vccd1 _07786_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_223_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09525_ _09933_/A _09525_/B vssd1 vssd1 vccd1 vccd1 _09525_/X sky130_fd_sc_hd__or2_1
XFILLER_0_56_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09456_ _09456_/A _09456_/B _09456_/C _09456_/D vssd1 vssd1 vccd1 vccd1 _09463_/D
+ sky130_fd_sc_hd__and4_2
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08407_ _15521_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08407_/X sky130_fd_sc_hd__or2_1
X_09387_ _15480_/A _09386_/X _07809_/B vssd1 vssd1 vccd1 vccd1 _09387_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_46_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08338_ hold337/A hold509/A _09399_/C vssd1 vssd1 vccd1 vccd1 hold113/A sky130_fd_sc_hd__or3_1
XFILLER_0_34_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08269_ hold2420/X _08268_/B _08268_/Y _09272_/A vssd1 vssd1 vccd1 vccd1 _08269_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10300_ hold3556/X _10604_/B _10299_/X _14863_/C1 vssd1 vssd1 vccd1 vccd1 _10300_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11280_ _11670_/A _11280_/B vssd1 vssd1 vccd1 vccd1 _11280_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5240 _11569_/X vssd1 vssd1 vccd1 vccd1 _17013_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10231_ hold3330/X _10637_/B _10230_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10231_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5251 _17152_/Q vssd1 vssd1 vccd1 vccd1 hold5251/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5262 _11371_/X vssd1 vssd1 vccd1 vccd1 _16947_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5273 _16870_/Q vssd1 vssd1 vccd1 vccd1 hold5273/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5284 _13567_/X vssd1 vssd1 vccd1 vccd1 _17642_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5295 _17199_/Q vssd1 vssd1 vccd1 vccd1 hold5295/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4550 _11757_/Y vssd1 vssd1 vccd1 vccd1 _11758_/B sky130_fd_sc_hd__dlygate4sd3_1
X_10162_ hold3987/X _10646_/B _10161_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10162_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4561 _17260_/Q vssd1 vssd1 vccd1 vccd1 hold4561/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4572 _10549_/X vssd1 vssd1 vccd1 vccd1 _16673_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4583 _17268_/Q vssd1 vssd1 vccd1 vccd1 hold4583/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4594 _16608_/Q vssd1 vssd1 vccd1 vccd1 hold4594/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3860 _16407_/Q vssd1 vssd1 vccd1 vccd1 hold3860/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10093_ hold3274/X _10571_/B _10092_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _10093_/X
+ sky130_fd_sc_hd__o211a_1
X_14970_ _14970_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14970_/X sky130_fd_sc_hd__or2_1
Xhold3871 _12118_/X vssd1 vssd1 vccd1 vccd1 _17196_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3882 _16644_/Q vssd1 vssd1 vccd1 vccd1 hold3882/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3893 hold6124/X vssd1 vssd1 vccd1 vccd1 hold3893/X sky130_fd_sc_hd__buf_2
XFILLER_0_156_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13921_ _13941_/A _13921_/B vssd1 vssd1 vccd1 vccd1 _17768_/D sky130_fd_sc_hd__and2_1
XFILLER_0_215_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16640_ _18231_/CLK _16640_/D vssd1 vssd1 vccd1 vccd1 _16640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13852_ _13888_/A _13852_/B vssd1 vssd1 vccd1 vccd1 _13852_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12803_ hold3752/X _12802_/X _12839_/S vssd1 vssd1 vccd1 vccd1 _12804_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_230_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16571_ _18129_/CLK _16571_/D vssd1 vssd1 vccd1 vccd1 _16571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13783_ hold5573/X _13877_/B _13782_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _13783_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_230_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10995_ _11091_/A _10995_/B vssd1 vssd1 vccd1 vccd1 _10995_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18310_ _18342_/CLK _18310_/D vssd1 vssd1 vccd1 vccd1 _18310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15522_ hold2683/X _15560_/A2 _15521_/X _12873_/A vssd1 vssd1 vccd1 vccd1 _15522_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12734_ hold3156/X _12733_/X _12749_/S vssd1 vssd1 vccd1 vccd1 _12734_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18241_ _18373_/CLK _18241_/D vssd1 vssd1 vccd1 vccd1 _18241_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _15481_/A1 _15445_/X _15452_/X _15481_/B1 hold5955/A vssd1 vssd1 vccd1 vccd1
+ _15453_/X sky130_fd_sc_hd__a32o_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ hold3151/X _12664_/X _12851_/S vssd1 vssd1 vccd1 vccd1 _12666_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14404_ hold2392/X _14446_/A2 _14403_/X _14526_/C1 vssd1 vssd1 vccd1 vccd1 _14404_/X
+ sky130_fd_sc_hd__o211a_1
X_18172_ _18172_/CLK _18172_/D vssd1 vssd1 vccd1 vccd1 _18172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11616_ _12093_/A _11616_/B vssd1 vssd1 vccd1 vccd1 _11616_/X sky130_fd_sc_hd__or2_1
X_15384_ _15482_/A _15384_/B vssd1 vssd1 vccd1 vccd1 _18414_/D sky130_fd_sc_hd__and2_1
X_12596_ hold3290/X _12595_/X _12923_/S vssd1 vssd1 vccd1 vccd1 _12596_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17123_ _17735_/CLK _17123_/D vssd1 vssd1 vccd1 vccd1 _17123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14335_ hold2813/X _14326_/B _14334_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _14335_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11547_ _11649_/A _11547_/B vssd1 vssd1 vccd1 vccd1 _11547_/X sky130_fd_sc_hd__or2_1
XFILLER_0_167_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_1410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold509 hold509/A vssd1 vssd1 vccd1 vccd1 hold509/X sky130_fd_sc_hd__buf_2
X_17054_ _17902_/CLK _17054_/D vssd1 vssd1 vccd1 vccd1 _17054_/Q sky130_fd_sc_hd__dfxtp_1
X_14266_ _15541_/A _14268_/B vssd1 vssd1 vccd1 vccd1 _14266_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_204_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11478_ _11670_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11478_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_1416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16005_ _18425_/CLK _16005_/D vssd1 vssd1 vccd1 vccd1 hold660/A sky130_fd_sc_hd__dfxtp_1
X_13217_ _13217_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13217_/X sky130_fd_sc_hd__and2_1
XFILLER_0_21_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10429_ hold3296/X _10619_/B _10428_/X _14853_/C1 vssd1 vssd1 vccd1 vccd1 _10429_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14197_ hold3014/X _14198_/B _14196_/Y _13931_/A vssd1 vssd1 vccd1 vccd1 _14197_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_221_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_374_wb_clk_i clkbuf_6_32_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17697_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ hold4309/X _13147_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13148_/X sky130_fd_sc_hd__mux2_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_303_wb_clk_i clkbuf_6_44_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17834_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13079_ _13199_/A1 _13077_/X _13078_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13079_/X
+ sky130_fd_sc_hd__o211a_1
X_17956_ _18052_/CLK _17956_/D vssd1 vssd1 vccd1 vccd1 _17956_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1209 _18140_/Q vssd1 vssd1 vccd1 vccd1 hold1209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16907_ _17883_/CLK _16907_/D vssd1 vssd1 vccd1 vccd1 _16907_/Q sky130_fd_sc_hd__dfxtp_1
X_17887_ _17887_/CLK _17887_/D vssd1 vssd1 vccd1 vccd1 _17887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16838_ _18041_/CLK _16838_/D vssd1 vssd1 vccd1 vccd1 _16838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16769_ _18036_/CLK _16769_/D vssd1 vssd1 vccd1 vccd1 _16769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09310_ hold1400/X _09323_/B _09309_/X _14358_/A vssd1 vssd1 vccd1 vccd1 _09310_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09241_ _15517_/A hold2284/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09242_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_118_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18439_ _18452_/CLK _18439_/D vssd1 vssd1 vccd1 vccd1 _18439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_90_wb_clk_i clkbuf_6_17_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16093_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_134_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09172_ _15555_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09172_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08123_ _08133_/A _08123_/B vssd1 vssd1 vccd1 vccd1 _15700_/D sky130_fd_sc_hd__and2_1
XFILLER_0_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_6_22_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_22_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08054_ _15513_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08054_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_228_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3101 _14931_/X vssd1 vssd1 vccd1 vccd1 _18252_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3112 _17952_/Q vssd1 vssd1 vccd1 vccd1 hold3112/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3123 _12671_/X vssd1 vssd1 vccd1 vccd1 _12672_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3134 _12662_/X vssd1 vssd1 vccd1 vccd1 _12663_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2400 _15754_/Q vssd1 vssd1 vccd1 vccd1 hold2400/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3145 _17399_/Q vssd1 vssd1 vccd1 vccd1 hold3145/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3156 _17421_/Q vssd1 vssd1 vccd1 vccd1 hold3156/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2411 _07850_/X vssd1 vssd1 vccd1 vccd1 _15570_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2422 _18365_/Q vssd1 vssd1 vccd1 vccd1 hold2422/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3167 _18025_/Q vssd1 vssd1 vccd1 vccd1 hold3167/X sky130_fd_sc_hd__dlygate4sd3_1
X_08956_ _15473_/A hold211/X vssd1 vssd1 vccd1 vccd1 _16095_/D sky130_fd_sc_hd__and2_1
Xhold3178 _17425_/Q vssd1 vssd1 vccd1 vccd1 hold3178/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2433 _15658_/Q vssd1 vssd1 vccd1 vccd1 hold2433/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3189 _10053_/Y vssd1 vssd1 vccd1 vccd1 _10054_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2444 _14540_/X vssd1 vssd1 vccd1 vccd1 _18066_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1710 _18428_/Q vssd1 vssd1 vccd1 vccd1 hold1710/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2455 _17799_/Q vssd1 vssd1 vccd1 vccd1 hold2455/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1721 _08481_/X vssd1 vssd1 vccd1 vccd1 _15869_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2466 _15767_/Q vssd1 vssd1 vccd1 vccd1 hold2466/X sky130_fd_sc_hd__dlygate4sd3_1
X_07907_ hold2567/X _07918_/B _07906_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _07907_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1732 _18127_/Q vssd1 vssd1 vccd1 vccd1 hold1732/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2477 _07979_/X vssd1 vssd1 vccd1 vccd1 _15632_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08887_ _15414_/A _08887_/B vssd1 vssd1 vccd1 vccd1 _16061_/D sky130_fd_sc_hd__and2_1
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1743 _14059_/X vssd1 vssd1 vccd1 vccd1 _17834_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2488 _14175_/X vssd1 vssd1 vccd1 vccd1 _17890_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1754 _18201_/Q vssd1 vssd1 vccd1 vccd1 hold1754/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2499 _15798_/Q vssd1 vssd1 vccd1 vccd1 hold2499/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1765 _14615_/X vssd1 vssd1 vccd1 vccd1 _18101_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07838_ hold2993/X _07865_/B _07837_/X _12289_/C1 vssd1 vssd1 vccd1 vccd1 _07838_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1776 _07834_/X vssd1 vssd1 vccd1 vccd1 _15562_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1787 _17790_/Q vssd1 vssd1 vccd1 vccd1 hold1787/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1798 _14991_/X vssd1 vssd1 vccd1 vccd1 _18281_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09508_ hold4847/X _09992_/B _09507_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _09508_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10780_ hold5215/X _11162_/B _10779_/X _14372_/A vssd1 vssd1 vccd1 vccd1 _10780_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_6_61_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_61_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ hold1418/X _07804_/A _15284_/A _09438_/X vssd1 vssd1 vccd1 vccd1 _09439_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _17318_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12450_/X sky130_fd_sc_hd__or2_1
XFILLER_0_227_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11401_ hold5665/X _12329_/B _11400_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _11401_/X
+ sky130_fd_sc_hd__o211a_1
X_12381_ hold226/X hold726/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold727/A sky130_fd_sc_hd__mux2_1
XFILLER_0_35_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_80 hold1253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_91 hold5974/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14120_ _15193_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14120_/X sky130_fd_sc_hd__or2_1
X_11332_ hold5614/X _11717_/B _11331_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11332_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14051_ hold1201/X _14040_/B _14050_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _14051_/X
+ sky130_fd_sc_hd__o211a_1
X_11263_ hold4877/X _11165_/B _11262_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _11263_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5070 _16855_/Q vssd1 vssd1 vccd1 vccd1 hold5070/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13002_ _15244_/A _13002_/B vssd1 vssd1 vccd1 vccd1 _17510_/D sky130_fd_sc_hd__and2_1
Xhold5081 _09826_/X vssd1 vssd1 vccd1 vccd1 _16432_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10214_ hold2047/X _16562_/Q _10634_/C vssd1 vssd1 vccd1 vccd1 _10215_/B sky130_fd_sc_hd__mux2_1
Xhold5092 _16600_/Q vssd1 vssd1 vccd1 vccd1 hold5092/X sky130_fd_sc_hd__dlygate4sd3_1
X_11194_ _11218_/A _11194_/B vssd1 vssd1 vccd1 vccd1 _11194_/Y sky130_fd_sc_hd__nor2_1
XTAP_6520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4380 _13837_/Y vssd1 vssd1 vccd1 vccd1 _17732_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10145_ hold2824/X hold3420/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10146_/B sky130_fd_sc_hd__mux2_1
X_17810_ _17873_/CLK _17810_/D vssd1 vssd1 vccd1 vccd1 _17810_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4391 _11790_/Y vssd1 vssd1 vccd1 vccd1 _11791_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3690 _16645_/Q vssd1 vssd1 vccd1 vccd1 hold3690/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17741_ _17741_/CLK _17741_/D vssd1 vssd1 vccd1 vccd1 _17741_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14953_ hold1000/X _14952_/B _14952_/Y _15226_/C1 vssd1 vssd1 vccd1 vccd1 _14953_/X
+ sky130_fd_sc_hd__o211a_1
X_10076_ _18074_/Q _16516_/Q _10634_/C vssd1 vssd1 vccd1 vccd1 _10077_/B sky130_fd_sc_hd__mux2_1
XTAP_5874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13904_ _15085_/A hold957/X hold297/X vssd1 vssd1 vccd1 vccd1 hold958/A sky130_fd_sc_hd__mux2_1
X_17672_ _17672_/CLK _17672_/D vssd1 vssd1 vccd1 vccd1 _17672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14884_ hold484/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14884_/X sky130_fd_sc_hd__or2_1
XFILLER_0_72_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16623_ _18149_/CLK _16623_/D vssd1 vssd1 vccd1 vccd1 _16623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13835_ _17732_/Q _13856_/B _13871_/C vssd1 vssd1 vccd1 vccd1 _13835_/X sky130_fd_sc_hd__and3_1
XFILLER_0_159_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16554_ _18176_/CLK _16554_/D vssd1 vssd1 vccd1 vccd1 _16554_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13766_ hold1397/X hold3696/X _13766_/S vssd1 vssd1 vccd1 vccd1 _13767_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10978_ hold5523/X _11071_/A2 _10977_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _10978_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15505_ _15521_/A hold2222/X _15505_/S vssd1 vssd1 vccd1 vccd1 _15506_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_128_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12717_ _12810_/A _12717_/B vssd1 vssd1 vccd1 vccd1 _17415_/D sky130_fd_sc_hd__and2_1
X_16485_ _18398_/CLK _16485_/D vssd1 vssd1 vccd1 vccd1 _16485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13697_ hold2466/X hold3728/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13698_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_72_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18224_ _18224_/CLK _18224_/D vssd1 vssd1 vccd1 vccd1 _18224_/Q sky130_fd_sc_hd__dfxtp_1
X_15436_ _17319_/Q _15487_/A2 _09392_/A hold283/X vssd1 vssd1 vccd1 vccd1 _15436_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12648_ _12822_/A _12648_/B vssd1 vssd1 vccd1 vccd1 _17392_/D sky130_fd_sc_hd__and2_1
XFILLER_0_25_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18155_ _18181_/CLK _18155_/D vssd1 vssd1 vccd1 vccd1 _18155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15367_ hold124/X _15487_/A2 _15484_/B1 hold324/X _15366_/X vssd1 vssd1 vccd1 vccd1
+ _15372_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_136_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12579_ _12894_/A _12579_/B vssd1 vssd1 vccd1 vccd1 _17369_/D sky130_fd_sc_hd__and2_1
XFILLER_0_68_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17106_ _17209_/CLK _17106_/D vssd1 vssd1 vccd1 vccd1 _17106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14318_ _14604_/A _14334_/B vssd1 vssd1 vccd1 vccd1 _14318_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_230_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18086_ _18106_/CLK _18086_/D vssd1 vssd1 vccd1 vccd1 _18086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15298_ hold497/X _15484_/A2 _09392_/D hold274/X vssd1 vssd1 vccd1 vccd1 _15298_/X
+ sky130_fd_sc_hd__a22o_1
Xhold306 hold306/A vssd1 vssd1 vccd1 vccd1 hold306/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 hold317/A vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold328 hold402/X vssd1 vssd1 vccd1 vccd1 hold403/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold339 hold339/A vssd1 vssd1 vccd1 vccd1 hold339/X sky130_fd_sc_hd__dlygate4sd3_1
X_17037_ _17885_/CLK _17037_/D vssd1 vssd1 vccd1 vccd1 _17037_/Q sky130_fd_sc_hd__dfxtp_1
X_14249_ hold1047/X _14268_/B _14248_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _14249_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout808 _15070_/A vssd1 vssd1 vccd1 vccd1 _15146_/C1 sky130_fd_sc_hd__buf_4
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout819 _10564_/C1 vssd1 vssd1 vccd1 vccd1 _14875_/C1 sky130_fd_sc_hd__buf_4
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_237_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08810_ hold684/X hold827/X _08866_/S vssd1 vssd1 vccd1 vccd1 hold828/A sky130_fd_sc_hd__mux2_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09790_ hold5829/X _10022_/B _09789_/X _15202_/C1 vssd1 vssd1 vccd1 vccd1 _09790_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1006 input39/X vssd1 vssd1 vccd1 vccd1 hold520/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1017 _18241_/Q vssd1 vssd1 vccd1 vccd1 hold1017/X sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ hold147/X hold593/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08742_/B sky130_fd_sc_hd__mux2_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1028 _14464_/X vssd1 vssd1 vccd1 vccd1 _18029_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17939_ _17971_/CLK _17939_/D vssd1 vssd1 vccd1 vccd1 _17939_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1039 _15568_/Q vssd1 vssd1 vccd1 vccd1 hold1039/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08672_ _15434_/A hold719/X vssd1 vssd1 vccd1 vccd1 _15957_/D sky130_fd_sc_hd__and2_1
XFILLER_0_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09224_ _15553_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09224_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09155_ hold2092/X _09164_/B _09154_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _09155_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08106_ _14166_/A hold1305/X hold108/X vssd1 vssd1 vccd1 vccd1 _08106_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_296_wb_clk_i clkbuf_6_39_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18060_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09086_ hold951/X _09098_/B vssd1 vssd1 vccd1 vccd1 _09086_/X sky130_fd_sc_hd__or2_1
XFILLER_0_13_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_225_wb_clk_i clkbuf_6_63_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18229_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08037_ _14330_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08037_/X sky130_fd_sc_hd__or2_1
Xhold840 hold988/X vssd1 vssd1 vccd1 vccd1 hold989/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 hold851/A vssd1 vssd1 vccd1 vccd1 hold851/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 hold862/A vssd1 vssd1 vccd1 vccd1 hold862/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold873 hold873/A vssd1 vssd1 vccd1 vccd1 hold873/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold884 hold884/A vssd1 vssd1 vccd1 vccd1 hold884/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold895 hold903/X vssd1 vssd1 vccd1 vccd1 hold904/A sky130_fd_sc_hd__clkbuf_2
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09988_ _13078_/A _09992_/B _09987_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _16486_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2230 _08302_/X vssd1 vssd1 vccd1 vccd1 _15784_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2241 _18079_/Q vssd1 vssd1 vccd1 vccd1 hold2241/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2252 input4/X vssd1 vssd1 vccd1 vccd1 hold920/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08939_ hold131/X hold663/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold664/A sky130_fd_sc_hd__mux2_1
Xhold2263 hold2268/X vssd1 vssd1 vccd1 vccd1 hold2269/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2274 _18462_/Q vssd1 vssd1 vccd1 vccd1 _07789_/A sky130_fd_sc_hd__buf_1
XFILLER_0_235_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1540 la_data_in[6] vssd1 vssd1 vccd1 vccd1 hold1540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2285 _15845_/Q vssd1 vssd1 vccd1 vccd1 hold2285/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2296 _14663_/X vssd1 vssd1 vccd1 vccd1 _18124_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1551 _14033_/X vssd1 vssd1 vccd1 vccd1 _17822_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ hold5749/X _12350_/B _11949_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _11950_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1562 _15587_/Q vssd1 vssd1 vccd1 vccd1 hold1562/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1573 _09207_/X vssd1 vssd1 vccd1 vccd1 _16215_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1584 _14337_/X vssd1 vssd1 vccd1 vccd1 _17968_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10901_ hold1169/X _16791_/Q _11216_/C vssd1 vssd1 vccd1 vccd1 _10902_/B sky130_fd_sc_hd__mux2_1
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1595 _08398_/X vssd1 vssd1 vccd1 vccd1 _15829_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11881_ hold5735/X _12332_/B _11880_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _11881_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13620_ _13716_/A _13620_/B vssd1 vssd1 vccd1 vccd1 _13620_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10832_ hold1620/X hold5227/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10833_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13551_ _13773_/A _13551_/B vssd1 vssd1 vccd1 vccd1 _13551_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10763_ hold1101/X _16745_/Q _11144_/C vssd1 vssd1 vccd1 vccd1 _10764_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_94_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12502_ _17344_/Q _12506_/B vssd1 vssd1 vccd1 vccd1 _12502_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16270_ _17881_/CLK _16270_/D vssd1 vssd1 vccd1 vccd1 _16270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13482_ _13482_/A _13482_/B vssd1 vssd1 vccd1 vccd1 _13482_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10694_ hold1047/X hold3483/X _11210_/C vssd1 vssd1 vccd1 vccd1 _10695_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15221_ _15221_/A _15221_/B vssd1 vssd1 vccd1 vccd1 _15221_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12433_ hold315/X hold514/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12434_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15152_ hold1374/X _15167_/B _15151_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _15152_/X
+ sky130_fd_sc_hd__o211a_1
X_12364_ _13873_/A _12364_/B vssd1 vssd1 vccd1 vccd1 _12364_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_65_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14103_ hold6057/X _14107_/A2 hold709/X _13905_/A vssd1 vssd1 vccd1 vccd1 hold710/A
+ sky130_fd_sc_hd__o211a_1
X_11315_ hold2821/X hold4411/X _12335_/C vssd1 vssd1 vccd1 vccd1 _11316_/B sky130_fd_sc_hd__mux2_1
X_15083_ _15191_/A _15119_/B vssd1 vssd1 vccd1 vccd1 _15083_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12295_ _13819_/A _12295_/B vssd1 vssd1 vccd1 vccd1 _12295_/Y sky130_fd_sc_hd__nor2_1
X_14034_ _15541_/A _14038_/B vssd1 vssd1 vccd1 vccd1 _14034_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_238_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11246_ hold2222/X hold4454/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11247_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11177_ _16883_/Q _11204_/B _11204_/C vssd1 vssd1 vccd1 vccd1 _11177_/X sky130_fd_sc_hd__and3_1
XTAP_6361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10128_ _10536_/A _10128_/B vssd1 vssd1 vccd1 vccd1 _10128_/X sky130_fd_sc_hd__or2_1
XFILLER_0_101_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15985_ _16147_/CLK _15985_/D vssd1 vssd1 vccd1 vccd1 hold523/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10059_ _13270_/A _10539_/A _10058_/X vssd1 vssd1 vccd1 vccd1 _10059_/Y sky130_fd_sc_hd__a21oi_1
X_14936_ _15205_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14936_/X sky130_fd_sc_hd__or2_1
X_17724_ _17724_/CLK _17724_/D vssd1 vssd1 vccd1 vccd1 _17724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_wb_clk_i clkbuf_6_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17881_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14867_ hold1980/X hold332/X _14866_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14867_/X
+ sky130_fd_sc_hd__o211a_1
X_17655_ _17720_/CLK _17655_/D vssd1 vssd1 vccd1 vccd1 _17655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16606_ _18164_/CLK _16606_/D vssd1 vssd1 vccd1 vccd1 _16606_/Q sky130_fd_sc_hd__dfxtp_1
X_13818_ hold4335/X _13722_/A _13817_/X vssd1 vssd1 vccd1 vccd1 _13819_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_230_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17586_ _17653_/CLK _17586_/D vssd1 vssd1 vccd1 vccd1 _17586_/Q sky130_fd_sc_hd__dfxtp_1
X_14798_ _15191_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14798_/X sky130_fd_sc_hd__or2_1
XFILLER_0_159_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16537_ _18223_/CLK _16537_/D vssd1 vssd1 vccd1 vccd1 _16537_/Q sky130_fd_sc_hd__dfxtp_1
X_13749_ _13749_/A _13749_/B vssd1 vssd1 vccd1 vccd1 _13749_/X sky130_fd_sc_hd__or2_1
XFILLER_0_73_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16468_ _18381_/CLK _16468_/D vssd1 vssd1 vccd1 vccd1 _16468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15419_ hold791/X _09386_/A _15417_/X vssd1 vssd1 vccd1 vccd1 _15422_/B sky130_fd_sc_hd__a21o_1
X_18207_ _18235_/CLK _18207_/D vssd1 vssd1 vccd1 vccd1 _18207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16399_ _18349_/CLK _16399_/D vssd1 vssd1 vccd1 vccd1 _16399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18138_ _18234_/CLK _18138_/D vssd1 vssd1 vccd1 vccd1 _18138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5806 _12040_/X vssd1 vssd1 vccd1 vccd1 _17170_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5817 _16496_/Q vssd1 vssd1 vccd1 vccd1 hold5817/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold103 hold103/A vssd1 vssd1 vccd1 vccd1 hold103/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5828 _09916_/X vssd1 vssd1 vccd1 vccd1 _16462_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5839 _16484_/Q vssd1 vssd1 vccd1 vccd1 hold5839/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 hold114/A vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__clkbuf_2
Xhold125 hold125/A vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18069_ _18069_/CLK _18069_/D vssd1 vssd1 vccd1 vccd1 _18069_/Q sky130_fd_sc_hd__dfxtp_1
Xhold136 hold136/A vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 hold394/X vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__buf_4
Xhold158 hold683/X vssd1 vssd1 vccd1 vccd1 hold684/A sky130_fd_sc_hd__buf_1
X_09911_ hold1968/X hold3574/X _10025_/C vssd1 vssd1 vccd1 vccd1 _09912_/B sky130_fd_sc_hd__mux2_1
Xhold169 hold59/X vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__buf_4
XFILLER_0_223_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout605 _09366_/Y vssd1 vssd1 vccd1 vccd1 _15484_/B1 sky130_fd_sc_hd__buf_8
Xfanout616 _09356_/Y vssd1 vssd1 vccd1 vccd1 _15446_/B1 sky130_fd_sc_hd__buf_6
Xfanout627 _09339_/Y vssd1 vssd1 vccd1 vccd1 _15481_/A1 sky130_fd_sc_hd__clkbuf_8
X_09842_ hold3184/X hold4169/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09843_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_0_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout638 _12849_/A vssd1 vssd1 vccd1 vccd1 _12843_/A sky130_fd_sc_hd__buf_4
XFILLER_0_42_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout649 _12855_/A vssd1 vssd1 vccd1 vccd1 _12864_/A sky130_fd_sc_hd__buf_4
XFILLER_0_158_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09773_ _18328_/Q hold3216/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09774_/B sky130_fd_sc_hd__mux2_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _12420_/A hold496/X vssd1 vssd1 vccd1 vccd1 _15983_/D sky130_fd_sc_hd__and2_1
XFILLER_0_213_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ hold87/X hold102/X _08657_/S vssd1 vssd1 vccd1 vccd1 hold103/A sky130_fd_sc_hd__mux2_1
XFILLER_0_178_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08586_ hold82/X hold498/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold499/A sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_228_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09207_ hold1572/X _09214_/B _09206_/X _12822_/A vssd1 vssd1 vccd1 vccd1 _09207_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_406_wb_clk_i clkbuf_6_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17888_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_173_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09138_ _15521_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09138_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09069_ hold1618/X _09106_/B _09068_/X _12948_/A vssd1 vssd1 vccd1 vccd1 _09069_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11100_ _11100_/A _11100_/B vssd1 vssd1 vccd1 vccd1 _11100_/X sky130_fd_sc_hd__or2_1
X_12080_ hold1170/X hold4046/X _13886_/C vssd1 vssd1 vccd1 vccd1 _12081_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold670 data_in[9] vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 data_in[3] vssd1 vssd1 vccd1 vccd1 hold681/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold692 hold692/A vssd1 vssd1 vccd1 vccd1 hold692/X sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ _11694_/A _11031_/B vssd1 vssd1 vccd1 vccd1 _11031_/X sky130_fd_sc_hd__or2_1
XFILLER_0_217_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2060 _16173_/Q vssd1 vssd1 vccd1 vccd1 hold2060/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2071 _17853_/Q vssd1 vssd1 vccd1 vccd1 hold2071/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2082 _15011_/X vssd1 vssd1 vccd1 vccd1 _18291_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15770_ _17689_/CLK _15770_/D vssd1 vssd1 vccd1 vccd1 _15770_/Q sky130_fd_sc_hd__dfxtp_1
X_12982_ hold2468/X hold3748/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12982_/X sky130_fd_sc_hd__mux2_1
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2093 _09155_/X vssd1 vssd1 vccd1 vccd1 _16190_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1370 _15770_/Q vssd1 vssd1 vccd1 vccd1 hold1370/X sky130_fd_sc_hd__dlygate4sd3_1
X_14721_ hold1058/X _14720_/B _14720_/Y _14895_/C1 vssd1 vssd1 vccd1 vccd1 _14721_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1381 _08475_/X vssd1 vssd1 vccd1 vccd1 _15866_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ hold2655/X _17135_/Q _12317_/C vssd1 vssd1 vccd1 vccd1 _11934_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_99_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1392 _13890_/X vssd1 vssd1 vccd1 vccd1 _17750_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _17440_/CLK _17440_/D vssd1 vssd1 vccd1 vccd1 _17440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _15099_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14652_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ hold1411/X hold3453/X _12371_/C vssd1 vssd1 vccd1 vccd1 _11865_/B sky130_fd_sc_hd__mux2_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13603_ hold3728/X _13795_/A2 _13602_/X _13795_/C1 vssd1 vssd1 vccd1 vccd1 _13603_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10815_ _11103_/A _10815_/B vssd1 vssd1 vccd1 vccd1 _10815_/X sky130_fd_sc_hd__or2_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17371_ _17881_/CLK _17371_/D vssd1 vssd1 vccd1 vccd1 _17371_/Q sky130_fd_sc_hd__dfxtp_1
X_14583_ hold2491/X _14610_/B _14582_/X _14691_/C1 vssd1 vssd1 vccd1 vccd1 _14583_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11795_ _17089_/Q _12335_/B _12335_/C vssd1 vssd1 vccd1 vccd1 _11795_/X sky130_fd_sc_hd__and3_1
X_16322_ _16323_/CLK _16322_/D vssd1 vssd1 vccd1 vccd1 _16322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13534_ hold4685/X _13829_/B _13533_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13534_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10746_ _11124_/A _10746_/B vssd1 vssd1 vccd1 vccd1 _10746_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_147_wb_clk_i clkbuf_6_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18421_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16253_ _17434_/CLK _16253_/D vssd1 vssd1 vccd1 vccd1 hold954/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13465_ hold5733/X _13868_/B _13464_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13465_/X
+ sky130_fd_sc_hd__o211a_1
X_10677_ _11067_/A _10677_/B vssd1 vssd1 vccd1 vccd1 _10677_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15204_ hold1199/X _15221_/B _15203_/X _15204_/C1 vssd1 vssd1 vccd1 vccd1 _15204_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12416_ _12416_/A _12416_/B vssd1 vssd1 vccd1 vccd1 _17301_/D sky130_fd_sc_hd__and2_1
XFILLER_0_207_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16184_ _17477_/CLK _16184_/D vssd1 vssd1 vccd1 vccd1 _16184_/Q sky130_fd_sc_hd__dfxtp_1
X_13396_ hold5325/X _13874_/B _13395_/X _08347_/A vssd1 vssd1 vccd1 vccd1 _13396_/X
+ sky130_fd_sc_hd__o211a_1
X_15135_ _15189_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15135_/X sky130_fd_sc_hd__or2_1
X_12347_ _17273_/Q _12350_/B _13463_/S vssd1 vssd1 vccd1 vccd1 _12347_/X sky130_fd_sc_hd__and3_1
XFILLER_0_51_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15066_ _15066_/A _15066_/B vssd1 vssd1 vccd1 vccd1 _18318_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12278_ hold1325/X _17250_/Q _13748_/S vssd1 vssd1 vccd1 vccd1 _12279_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14017_ hold1481/X _14038_/B _14016_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _14017_/X
+ sky130_fd_sc_hd__o211a_1
X_11229_ _11622_/A _11229_/B vssd1 vssd1 vccd1 vccd1 _11229_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15968_ _18410_/CLK _15968_/D vssd1 vssd1 vccd1 vccd1 hold832/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_218_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17707_ _17707_/CLK _17707_/D vssd1 vssd1 vccd1 vccd1 _17707_/Q sky130_fd_sc_hd__dfxtp_1
X_14919_ hold1853/X _14946_/B _14918_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _14919_/X
+ sky130_fd_sc_hd__o211a_1
X_15899_ _17319_/CLK _15899_/D vssd1 vssd1 vccd1 vccd1 hold849/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08440_ hold2542/X _08442_/A2 _08439_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _08440_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17638_ _17702_/CLK _17638_/D vssd1 vssd1 vccd1 vccd1 _17638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08371_ _08377_/A _08371_/B vssd1 vssd1 vccd1 vccd1 _15817_/D sky130_fd_sc_hd__and2_1
XFILLER_0_4_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17569_ _17599_/CLK _17569_/D vssd1 vssd1 vccd1 vccd1 _17569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5603 _17749_/Q vssd1 vssd1 vccd1 vccd1 hold5603/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5614 _16966_/Q vssd1 vssd1 vccd1 vccd1 hold5614/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5625 _11236_/X vssd1 vssd1 vccd1 vccd1 _16902_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5636 _11326_/X vssd1 vssd1 vccd1 vccd1 _16932_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4902 _11251_/X vssd1 vssd1 vccd1 vccd1 _16907_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5647 _16783_/Q vssd1 vssd1 vccd1 vccd1 hold5647/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4913 _17240_/Q vssd1 vssd1 vccd1 vccd1 hold4913/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5658 _11653_/X vssd1 vssd1 vccd1 vccd1 _17041_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4924 _12289_/X vssd1 vssd1 vccd1 vccd1 _17253_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5669 _16999_/Q vssd1 vssd1 vccd1 vccd1 hold5669/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4935 _16813_/Q vssd1 vssd1 vccd1 vccd1 hold4935/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4946 _10795_/X vssd1 vssd1 vccd1 vccd1 _16755_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4957 _16882_/Q vssd1 vssd1 vccd1 vccd1 hold4957/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout402 _14446_/A2 vssd1 vssd1 vccd1 vccd1 _14433_/B sky130_fd_sc_hd__buf_6
Xhold4968 _17231_/Q vssd1 vssd1 vccd1 vccd1 hold4968/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4979 _16820_/Q vssd1 vssd1 vccd1 vccd1 hold4979/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout413 _14162_/Y vssd1 vssd1 vccd1 vccd1 _14198_/B sky130_fd_sc_hd__buf_8
XFILLER_0_10_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout424 _13994_/B vssd1 vssd1 vccd1 vccd1 _13998_/B sky130_fd_sc_hd__buf_6
XFILLER_0_226_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout435 _13817_/C vssd1 vssd1 vccd1 vccd1 _13814_/C sky130_fd_sc_hd__clkbuf_8
Xfanout446 fanout485/X vssd1 vssd1 vccd1 vccd1 _12227_/S sky130_fd_sc_hd__buf_4
X_09825_ _11010_/A _09825_/B vssd1 vssd1 vccd1 vccd1 _09825_/X sky130_fd_sc_hd__or2_1
Xfanout457 _11168_/C vssd1 vssd1 vccd1 vccd1 _11654_/S sky130_fd_sc_hd__buf_6
XFILLER_0_201_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout468 _13877_/C vssd1 vssd1 vccd1 vccd1 _13880_/C sky130_fd_sc_hd__clkbuf_8
Xfanout479 _11774_/C vssd1 vssd1 vccd1 vccd1 _12173_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09756_ _09948_/A _09756_/B vssd1 vssd1 vccd1 vccd1 _09756_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08707_ hold373/X hold465/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08708_/B sky130_fd_sc_hd__mux2_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _10986_/A _09687_/B vssd1 vssd1 vccd1 vccd1 _09687_/X sky130_fd_sc_hd__or2_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08638_ _12390_/A _08638_/B vssd1 vssd1 vccd1 vccd1 _15941_/D sky130_fd_sc_hd__and2_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _15364_/A _08569_/B vssd1 vssd1 vccd1 vccd1 _15908_/D sky130_fd_sc_hd__and2_1
XFILLER_0_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10600_ _11206_/A _10600_/B vssd1 vssd1 vccd1 vccd1 _16690_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11580_ _12243_/A _11580_/B vssd1 vssd1 vccd1 vccd1 _11580_/X sky130_fd_sc_hd__or2_1
XFILLER_0_119_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10531_ hold3674/X _10625_/B _10530_/X _14893_/C1 vssd1 vssd1 vccd1 vccd1 _10531_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_240_wb_clk_i clkbuf_6_60_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18146_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13250_ _17582_/Q _17116_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13250_/X sky130_fd_sc_hd__mux2_1
X_10462_ hold5229/X _10070_/B _10461_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _10462_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12201_ _13716_/A _12201_/B vssd1 vssd1 vccd1 vccd1 _12201_/X sky130_fd_sc_hd__or2_1
X_13181_ _13180_/X hold6000/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13181_/X sky130_fd_sc_hd__mux2_1
X_10393_ hold3970/X _10619_/B _10392_/X _14853_/C1 vssd1 vssd1 vccd1 vccd1 _10393_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12132_ _12267_/A _12132_/B vssd1 vssd1 vccd1 vccd1 _12132_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12063_ _12255_/A _12063_/B vssd1 vssd1 vccd1 vccd1 _12063_/X sky130_fd_sc_hd__or2_1
X_16940_ _17820_/CLK _16940_/D vssd1 vssd1 vccd1 vccd1 _16940_/Q sky130_fd_sc_hd__dfxtp_1
X_11014_ hold5044/X _11204_/B _11013_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _11014_/X
+ sky130_fd_sc_hd__o211a_1
X_16871_ _18042_/CLK _16871_/D vssd1 vssd1 vccd1 vccd1 _16871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15822_ _17733_/CLK _15822_/D vssd1 vssd1 vccd1 vccd1 _15822_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15753_ _17672_/CLK _15753_/D vssd1 vssd1 vccd1 vccd1 _15753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12965_ hold3212/X _12964_/X _12971_/S vssd1 vssd1 vccd1 vccd1 _12965_/X sky130_fd_sc_hd__mux2_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14704_ _15205_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14704_/X sky130_fd_sc_hd__or2_1
X_11916_ _12210_/A _11916_/B vssd1 vssd1 vccd1 vccd1 _11916_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_399_wb_clk_i clkbuf_6_37_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17858_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_158_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15684_ _17144_/CLK _15684_/D vssd1 vssd1 vccd1 vccd1 _15684_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ hold3316/X _12895_/X _12923_/S vssd1 vssd1 vccd1 vccd1 _12896_/X sky130_fd_sc_hd__mux2_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ hold2765/X _14666_/B _14634_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _14635_/X
+ sky130_fd_sc_hd__o211a_1
X_17423_ _17426_/CLK _17423_/D vssd1 vssd1 vccd1 vccd1 _17423_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_328_wb_clk_i clkbuf_6_44_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17905_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11847_ _12159_/A _11847_/B vssd1 vssd1 vccd1 vccd1 _11847_/X sky130_fd_sc_hd__or2_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _15492_/A _14573_/B hold2231/X vssd1 vssd1 vccd1 vccd1 _14566_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_172_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17354_ _17517_/CLK _17354_/D vssd1 vssd1 vccd1 vccd1 _17354_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11778_ hold4364/X _12285_/A _11777_/X vssd1 vssd1 vccd1 vccd1 _11778_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16305_ _16315_/CLK _16305_/D vssd1 vssd1 vccd1 vccd1 _16305_/Q sky130_fd_sc_hd__dfxtp_1
X_13517_ hold1051/X _17626_/Q _13721_/S vssd1 vssd1 vccd1 vccd1 _13518_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_83_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17285_ _17328_/CLK _17285_/D vssd1 vssd1 vccd1 vccd1 hold808/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10729_ hold5317/X _11210_/B _10728_/X _14526_/C1 vssd1 vssd1 vccd1 vccd1 _10729_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14497_ _15231_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14497_/X sky130_fd_sc_hd__or2_1
XFILLER_0_71_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16236_ _17430_/CLK _16236_/D vssd1 vssd1 vccd1 vccd1 _16236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13448_ hold1372/X hold3838/X _13862_/C vssd1 vssd1 vccd1 vccd1 _13449_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16167_ _17512_/CLK _16167_/D vssd1 vssd1 vccd1 vccd1 _16167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13379_ hold1720/X hold4458/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13380_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4209 hold5915/X vssd1 vssd1 vccd1 vccd1 hold5916/A sky130_fd_sc_hd__buf_4
X_15118_ hold2220/X hold340/X _15117_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _15118_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_239_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_224_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16098_ _16098_/CLK _16098_/D vssd1 vssd1 vccd1 vccd1 hold588/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3508 _16712_/Q vssd1 vssd1 vccd1 vccd1 hold3508/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3519 _11200_/Y vssd1 vssd1 vccd1 vccd1 _16890_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15049_ _15103_/A hold1621/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15050_/B sky130_fd_sc_hd__mux2_1
X_07940_ _14395_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07940_/X sky130_fd_sc_hd__or2_1
Xhold2807 _15779_/Q vssd1 vssd1 vccd1 vccd1 hold2807/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2818 _14129_/X vssd1 vssd1 vccd1 vccd1 _17868_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2829 _07965_/X vssd1 vssd1 vccd1 vccd1 _15625_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_44_wb_clk_i clkbuf_6_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17883_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07871_ _15549_/A _07871_/B vssd1 vssd1 vccd1 vccd1 _07871_/X sky130_fd_sc_hd__or2_1
XFILLER_0_236_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_235_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09610_ hold4679/X _09992_/B _09609_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _09610_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09541_ hold3620/X _10028_/B _09540_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _09541_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_1309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09472_ hold733/X hold739/X _09472_/C _09472_/D vssd1 vssd1 vccd1 vccd1 _09477_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_0_231_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08423_ _14477_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08423_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08354_ hold933/X hold1098/X hold115/X vssd1 vssd1 vccd1 vccd1 _08355_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_149_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08285_ _14395_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08285_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6101 la_data_in[31] vssd1 vssd1 vccd1 vccd1 hold358/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold6112 data_in[10] vssd1 vssd1 vccd1 vccd1 hold208/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6123 _16310_/Q vssd1 vssd1 vccd1 vccd1 hold6123/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6134 _17348_/Q vssd1 vssd1 vccd1 vccd1 hold6134/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5400 _17056_/Q vssd1 vssd1 vccd1 vccd1 hold5400/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5411 _11500_/X vssd1 vssd1 vccd1 vccd1 _16990_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5422 _16700_/Q vssd1 vssd1 vccd1 vccd1 hold5422/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5433 _13552_/X vssd1 vssd1 vccd1 vccd1 _17637_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5444 _17036_/Q vssd1 vssd1 vccd1 vccd1 hold5444/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4710 _13525_/X vssd1 vssd1 vccd1 vccd1 _17628_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5455 _11701_/X vssd1 vssd1 vccd1 vccd1 _17057_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4721 _09805_/X vssd1 vssd1 vccd1 vccd1 _16425_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5466 _17616_/Q vssd1 vssd1 vccd1 vccd1 hold5466/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5477 _13570_/X vssd1 vssd1 vccd1 vccd1 _17643_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4732 _13540_/X vssd1 vssd1 vccd1 vccd1 _17633_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4743 _17559_/Q vssd1 vssd1 vccd1 vccd1 hold4743/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5488 _16880_/Q vssd1 vssd1 vccd1 vccd1 hold5488/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4754 _16501_/Q vssd1 vssd1 vccd1 vccd1 hold4754/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5499 _13663_/X vssd1 vssd1 vccd1 vccd1 _17674_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4765 _13642_/X vssd1 vssd1 vccd1 vccd1 _17667_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4776 _09706_/X vssd1 vssd1 vccd1 vccd1 _16392_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout210 _09494_/X vssd1 vssd1 vccd1 vccd1 fanout210/X sky130_fd_sc_hd__buf_12
Xfanout221 _10013_/B vssd1 vssd1 vccd1 vccd1 _10025_/B sky130_fd_sc_hd__buf_4
Xhold4787 _17162_/Q vssd1 vssd1 vccd1 vccd1 hold4787/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout232 _10604_/B vssd1 vssd1 vccd1 vccd1 _10646_/B sky130_fd_sc_hd__clkbuf_8
Xhold4798 _12106_/X vssd1 vssd1 vccd1 vccd1 _17192_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout243 _10634_/B vssd1 vssd1 vccd1 vccd1 _10589_/B sky130_fd_sc_hd__buf_4
XFILLER_0_22_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout254 _13794_/A vssd1 vssd1 vccd1 vccd1 _13734_/A sky130_fd_sc_hd__buf_4
Xfanout265 fanout299/X vssd1 vssd1 vccd1 vccd1 _11043_/A sky130_fd_sc_hd__buf_2
Xfanout276 _12159_/A vssd1 vssd1 vccd1 vccd1 _12267_/A sky130_fd_sc_hd__buf_4
X_09808_ hold4650/X _11162_/B _09807_/X _14372_/A vssd1 vssd1 vccd1 vccd1 _09808_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout287 _11667_/A vssd1 vssd1 vccd1 vccd1 _12243_/A sky130_fd_sc_hd__buf_4
Xfanout298 fanout299/X vssd1 vssd1 vccd1 vccd1 _11127_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_213_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09739_ hold4618/X _10025_/B _09738_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09739_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12750_ _12750_/A _12750_/B vssd1 vssd1 vccd1 vccd1 _17426_/D sky130_fd_sc_hd__and2_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ hold5454/X _11798_/B _11700_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11701_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_421_wb_clk_i clkbuf_6_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17221_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12681_ _12843_/A _12681_/B vssd1 vssd1 vccd1 vccd1 _17403_/D sky130_fd_sc_hd__and2_1
XFILLER_0_166_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ hold2796/X _14433_/B _14419_/X _14552_/C1 vssd1 vssd1 vccd1 vccd1 _14420_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11632_ hold5663/X _11726_/B _11631_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _11632_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_182_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14351_ hold423/A _17975_/Q _14381_/S vssd1 vssd1 vccd1 vccd1 hold418/A sky130_fd_sc_hd__mux2_1
XFILLER_0_163_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11563_ hold5113/X _11753_/B _11562_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11563_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13302_ _13302_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13302_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10514_ hold2735/X _16662_/Q _10604_/C vssd1 vssd1 vccd1 vccd1 _10515_/B sky130_fd_sc_hd__mux2_1
X_17070_ _17886_/CLK _17070_/D vssd1 vssd1 vccd1 vccd1 _17070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14282_ _15231_/A _14282_/B vssd1 vssd1 vccd1 vccd1 _14282_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11494_ hold5529/X _12323_/B _11493_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _11494_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16021_ _17520_/CLK _16021_/D vssd1 vssd1 vccd1 vccd1 hold310/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13233_ _13233_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13233_/X sky130_fd_sc_hd__and2_1
XFILLER_0_165_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10445_ hold2879/X hold3785/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10446_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13164_ hold4251/X _13163_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13164_/X sky130_fd_sc_hd__mux2_2
X_10376_ hold2100/X _16616_/Q _10571_/C vssd1 vssd1 vccd1 vccd1 _10377_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_236_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12115_ hold5641/X _12299_/B _12114_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _12115_/X
+ sky130_fd_sc_hd__o211a_1
X_13095_ _13199_/A1 _13093_/X _13094_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13095_/X
+ sky130_fd_sc_hd__o211a_1
X_17972_ _18036_/CLK _17972_/D vssd1 vssd1 vccd1 vccd1 _17972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12046_ hold5743/X _12350_/B _12045_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _12046_/X
+ sky130_fd_sc_hd__o211a_1
X_16923_ _17771_/CLK _16923_/D vssd1 vssd1 vccd1 vccd1 _16923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_218_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16854_ _17929_/CLK _16854_/D vssd1 vssd1 vccd1 vccd1 _16854_/Q sky130_fd_sc_hd__dfxtp_1
X_15805_ _17716_/CLK _15805_/D vssd1 vssd1 vccd1 vccd1 _15805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13997_ hold2023/X _13986_/B _13996_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _13997_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16785_ _18020_/CLK _16785_/D vssd1 vssd1 vccd1 vccd1 _16785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12948_ _12948_/A _12948_/B vssd1 vssd1 vccd1 vccd1 _17492_/D sky130_fd_sc_hd__and2_1
X_15736_ _17733_/CLK _15736_/D vssd1 vssd1 vccd1 vccd1 _15736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_162_wb_clk_i clkbuf_6_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18416_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_158_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18455_ _18455_/CLK _18455_/D vssd1 vssd1 vccd1 vccd1 _18455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15667_ _17127_/CLK _15667_/D vssd1 vssd1 vccd1 vccd1 _15667_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ _12888_/A _12879_/B vssd1 vssd1 vccd1 vccd1 _17469_/D sky130_fd_sc_hd__and2_1
XFILLER_0_150_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_233_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17406_ _18457_/CLK _17406_/D vssd1 vssd1 vccd1 vccd1 _17406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14618_ _14726_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14618_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18386_ _18386_/CLK _18386_/D vssd1 vssd1 vccd1 vccd1 _18386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15598_ _17278_/CLK _15598_/D vssd1 vssd1 vccd1 vccd1 _15598_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17337_ _17337_/CLK hold48/X vssd1 vssd1 vccd1 vccd1 _17337_/Q sky130_fd_sc_hd__dfxtp_1
X_14549_ hold820/X _14553_/B vssd1 vssd1 vccd1 vccd1 hold821/A sky130_fd_sc_hd__or2_1
XFILLER_0_3_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_12_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_12_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_226_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08070_ _15529_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08070_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17268_ _17268_/CLK _17268_/D vssd1 vssd1 vccd1 vccd1 _17268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16219_ _17450_/CLK _16219_/D vssd1 vssd1 vccd1 vccd1 _16219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17199_ _17899_/CLK _17199_/D vssd1 vssd1 vccd1 vccd1 _17199_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4006 _12271_/X vssd1 vssd1 vccd1 vccd1 _17247_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4017 _10696_/X vssd1 vssd1 vccd1 vccd1 _16722_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4028 _17455_/Q vssd1 vssd1 vccd1 vccd1 hold4028/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4039 _17427_/Q vssd1 vssd1 vccd1 vccd1 hold4039/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3305 _17477_/Q vssd1 vssd1 vccd1 vccd1 hold3305/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3316 _17475_/Q vssd1 vssd1 vccd1 vccd1 hold3316/X sky130_fd_sc_hd__dlygate4sd3_1
X_08972_ _12420_/A hold246/X vssd1 vssd1 vccd1 vccd1 _16103_/D sky130_fd_sc_hd__and2_1
Xhold3327 _10267_/X vssd1 vssd1 vccd1 vccd1 _16579_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3338 _10399_/X vssd1 vssd1 vccd1 vccd1 _16623_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2604 _14203_/X vssd1 vssd1 vccd1 vccd1 _17904_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3349 _17461_/Q vssd1 vssd1 vccd1 vccd1 hold3349/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2615 _15808_/Q vssd1 vssd1 vccd1 vccd1 hold2615/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2626 _09185_/X vssd1 vssd1 vccd1 vccd1 _16204_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07923_ hold2474/X _07924_/B _07922_/Y _08115_/A vssd1 vssd1 vccd1 vccd1 _07923_/X
+ sky130_fd_sc_hd__o211a_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__buf_4
XFILLER_0_208_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2637 _18129_/Q vssd1 vssd1 vccd1 vccd1 hold2637/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1903 _18354_/Q vssd1 vssd1 vccd1 vccd1 hold1903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2648 _15630_/Q vssd1 vssd1 vccd1 vccd1 hold2648/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2659 _18143_/Q vssd1 vssd1 vccd1 vccd1 hold2659/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1914 _14903_/X vssd1 vssd1 vccd1 vccd1 _18239_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1925 _18217_/Q vssd1 vssd1 vccd1 vccd1 hold1925/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1936 _08235_/X vssd1 vssd1 vccd1 vccd1 _15752_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07854_ hold1205/X _07869_/B _07853_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _07854_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1947 _18081_/Q vssd1 vssd1 vccd1 vccd1 hold1947/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1958 _18270_/Q vssd1 vssd1 vccd1 vccd1 hold1958/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1969 _15184_/X vssd1 vssd1 vccd1 vccd1 _18374_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07785_ _09438_/B vssd1 vssd1 vccd1 vccd1 _07785_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_79_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09524_ hold1881/X _13126_/A _10028_/C vssd1 vssd1 vccd1 vccd1 _09525_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_51_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_51_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09455_ _09456_/A _09455_/B vssd1 vssd1 vccd1 vccd1 _09457_/C sky130_fd_sc_hd__or2_1
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08406_ hold1125/X _08442_/A2 _08405_/X _08363_/A vssd1 vssd1 vccd1 vccd1 _08406_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09386_ _09386_/A _09386_/B _09392_/C _09386_/D vssd1 vssd1 vccd1 vccd1 _09386_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_108_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08337_ hold444/X hold405/X vssd1 vssd1 vccd1 vccd1 _09399_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_163_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08268_ _15547_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08268_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_61_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08199_ _15533_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08199_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5230 _10462_/X vssd1 vssd1 vccd1 vccd1 _16644_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10230_ _10542_/A _10230_/B vssd1 vssd1 vccd1 vccd1 _10230_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5241 _16838_/Q vssd1 vssd1 vccd1 vccd1 hold5241/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5252 _11890_/X vssd1 vssd1 vccd1 vccd1 _17120_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5263 _17624_/Q vssd1 vssd1 vccd1 vccd1 hold5263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5274 _11044_/X vssd1 vssd1 vccd1 vccd1 _16838_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4540 _10264_/X vssd1 vssd1 vccd1 vccd1 _16578_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5285 _17680_/Q vssd1 vssd1 vccd1 vccd1 hold5285/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10161_ _10554_/A _10161_/B vssd1 vssd1 vccd1 vccd1 _10161_/X sky130_fd_sc_hd__or2_1
Xhold5296 _12031_/X vssd1 vssd1 vccd1 vccd1 _17167_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4551 _11758_/Y vssd1 vssd1 vccd1 vccd1 _17076_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4562 _12214_/X vssd1 vssd1 vccd1 vccd1 _17228_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4573 _16609_/Q vssd1 vssd1 vccd1 vccd1 hold4573/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4584 _12238_/X vssd1 vssd1 vccd1 vccd1 _17236_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4595 _10258_/X vssd1 vssd1 vccd1 vccd1 _16576_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3850 _16807_/Q vssd1 vssd1 vccd1 vccd1 hold3850/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3861 _09655_/X vssd1 vssd1 vccd1 vccd1 _16375_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10092_ _10560_/A _10092_/B vssd1 vssd1 vccd1 vccd1 _10092_/X sky130_fd_sc_hd__or2_1
XFILLER_0_22_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3872 _16743_/Q vssd1 vssd1 vccd1 vccd1 hold3872/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3883 _10366_/X vssd1 vssd1 vccd1 vccd1 _16612_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3894 _17415_/Q vssd1 vssd1 vccd1 vccd1 hold3894/X sky130_fd_sc_hd__dlygate4sd3_1
X_13920_ _14529_/A hold1413/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13921_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_233_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13851_ hold4495/X _13791_/A _13850_/X vssd1 vssd1 vccd1 vccd1 _13851_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_236_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12802_ hold1248/X hold3210/X _12838_/S vssd1 vssd1 vccd1 vccd1 _12802_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16570_ _18213_/CLK _16570_/D vssd1 vssd1 vccd1 vccd1 _16570_/Q sky130_fd_sc_hd__dfxtp_1
X_13782_ _13791_/A _13782_/B vssd1 vssd1 vccd1 vccd1 _13782_/X sky130_fd_sc_hd__or2_1
X_10994_ hold3167/X hold4911/X _11186_/C vssd1 vssd1 vccd1 vccd1 _10995_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ hold1237/X _17422_/Q _12811_/S vssd1 vssd1 vccd1 vccd1 _12733_/X sky130_fd_sc_hd__mux2_1
X_15521_ _15521_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15521_/X sky130_fd_sc_hd__or2_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15452_ _15489_/A _15452_/B _15452_/C _15452_/D vssd1 vssd1 vccd1 vccd1 _15452_/X
+ sky130_fd_sc_hd__or4_2
X_18240_ _18240_/CLK _18240_/D vssd1 vssd1 vccd1 vccd1 _18240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ hold2565/X hold3145/X _12850_/S vssd1 vssd1 vccd1 vccd1 _12664_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14403_ _14457_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14403_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11615_ hold2553/X hold4083/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11616_/B sky130_fd_sc_hd__mux2_1
X_18171_ _18177_/CLK _18171_/D vssd1 vssd1 vccd1 vccd1 _18171_/Q sky130_fd_sc_hd__dfxtp_1
X_15383_ _15481_/A1 _15375_/X _15382_/X _15481_/B1 hold5933/A vssd1 vssd1 vccd1 vccd1
+ _15383_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_136_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12595_ hold1552/X _17376_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12595_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_53_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14334_ _15229_/A _14334_/B vssd1 vssd1 vccd1 vccd1 _14334_/X sky130_fd_sc_hd__or2_1
X_17122_ _17187_/CLK _17122_/D vssd1 vssd1 vccd1 vccd1 _17122_/Q sky130_fd_sc_hd__dfxtp_1
X_11546_ hold2147/X _17006_/Q _11738_/C vssd1 vssd1 vccd1 vccd1 _11547_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17053_ _17901_/CLK _17053_/D vssd1 vssd1 vccd1 vccd1 _17053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14265_ hold2088/X _14272_/B _14264_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _14265_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11477_ hold1201/X _16983_/Q _11765_/C vssd1 vssd1 vccd1 vccd1 _11478_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16004_ _18411_/CLK _16004_/D vssd1 vssd1 vccd1 vccd1 hold478/A sky130_fd_sc_hd__dfxtp_1
X_13216_ _13209_/X _13215_/X _13296_/B1 vssd1 vssd1 vccd1 vccd1 _17545_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_208_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10428_ _10524_/A _10428_/B vssd1 vssd1 vccd1 vccd1 _10428_/X sky130_fd_sc_hd__or2_1
X_14196_ _15215_/A _14198_/B vssd1 vssd1 vccd1 vccd1 _14196_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _13146_/X _16911_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13147_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10359_ _10551_/A _10359_/B vssd1 vssd1 vccd1 vccd1 _10359_/X sky130_fd_sc_hd__or2_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13078_ _13078_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13078_/X sky130_fd_sc_hd__or2_1
X_17955_ _18051_/CLK _17955_/D vssd1 vssd1 vccd1 vccd1 _17955_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12029_ hold2338/X hold5129/X _12317_/C vssd1 vssd1 vccd1 vccd1 _12030_/B sky130_fd_sc_hd__mux2_1
X_16906_ _18432_/CLK _16906_/D vssd1 vssd1 vccd1 vccd1 _16906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17886_ _17886_/CLK _17886_/D vssd1 vssd1 vccd1 vccd1 _17886_/Q sky130_fd_sc_hd__dfxtp_1
X_16837_ _18072_/CLK _16837_/D vssd1 vssd1 vccd1 vccd1 _16837_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_343_wb_clk_i clkbuf_6_42_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17653_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_233_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16768_ _17971_/CLK _16768_/D vssd1 vssd1 vccd1 vccd1 _16768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15719_ _17157_/CLK _15719_/D vssd1 vssd1 vccd1 vccd1 _15719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16699_ _18115_/CLK _16699_/D vssd1 vssd1 vccd1 vccd1 _16699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09240_ _12786_/A _09240_/B vssd1 vssd1 vccd1 vccd1 _16231_/D sky130_fd_sc_hd__and2_1
X_18438_ _18438_/CLK _18438_/D vssd1 vssd1 vccd1 vccd1 _18438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_1371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09171_ hold2633/X _09177_/A2 _09170_/X _12924_/A vssd1 vssd1 vccd1 vccd1 _09171_/X
+ sky130_fd_sc_hd__o211a_1
X_18369_ _18369_/CLK hold843/X vssd1 vssd1 vccd1 vccd1 _18369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08122_ _14413_/A hold2582/X hold108/X vssd1 vssd1 vccd1 vccd1 _08123_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08053_ hold1716/X _08097_/A2 _08052_/X _08167_/A vssd1 vssd1 vccd1 vccd1 _08053_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3102 _18278_/Q vssd1 vssd1 vccd1 vccd1 hold3102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3113 _14305_/X vssd1 vssd1 vccd1 vccd1 _17952_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3124 _15699_/Q vssd1 vssd1 vccd1 vccd1 hold3124/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3135 _17384_/Q vssd1 vssd1 vccd1 vccd1 hold3135/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2401 _08239_/X vssd1 vssd1 vccd1 vccd1 _15754_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3146 _17394_/Q vssd1 vssd1 vccd1 vccd1 hold3146/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2412 _18352_/Q vssd1 vssd1 vccd1 vccd1 hold2412/X sky130_fd_sc_hd__dlygate4sd3_1
X_08955_ hold23/X _16095_/Q _08997_/S vssd1 vssd1 vccd1 vccd1 hold211/A sky130_fd_sc_hd__mux2_1
XTAP_5319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3157 _12734_/X vssd1 vssd1 vccd1 vccd1 _12735_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2423 _15164_/X vssd1 vssd1 vccd1 vccd1 _18365_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3168 _14456_/X vssd1 vssd1 vccd1 vccd1 _18025_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3179 _12746_/X vssd1 vssd1 vccd1 vccd1 _12747_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2434 _08034_/X vssd1 vssd1 vccd1 vccd1 _15658_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1700 _18135_/Q vssd1 vssd1 vccd1 vccd1 hold1700/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2445 _15645_/Q vssd1 vssd1 vccd1 vccd1 hold2445/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07906_ _15529_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07906_/X sky130_fd_sc_hd__or2_1
Xhold1711 _15497_/X vssd1 vssd1 vccd1 vccd1 _15498_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2456 _13985_/X vssd1 vssd1 vccd1 vccd1 _17799_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1722 _18398_/Q vssd1 vssd1 vccd1 vccd1 hold1722/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08886_ hold452/X hold806/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08887_/B sky130_fd_sc_hd__mux2_1
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2467 _08265_/X vssd1 vssd1 vccd1 vccd1 _15767_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1733 _14669_/X vssd1 vssd1 vccd1 vccd1 _18127_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2478 _15814_/Q vssd1 vssd1 vccd1 vccd1 hold2478/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1744 _15751_/Q vssd1 vssd1 vccd1 vccd1 hold1744/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2489 _17855_/Q vssd1 vssd1 vccd1 vccd1 hold2489/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1755 _14823_/X vssd1 vssd1 vccd1 vccd1 _18201_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1766 _18154_/Q vssd1 vssd1 vccd1 vccd1 hold1766/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07837_ _15515_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07837_/X sky130_fd_sc_hd__or2_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_1372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1777 _17981_/Q vssd1 vssd1 vccd1 vccd1 hold1777/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1788 _13967_/X vssd1 vssd1 vccd1 vccd1 _17790_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1799 _18037_/Q vssd1 vssd1 vccd1 vccd1 hold1799/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09507_ _09987_/A _09507_/B vssd1 vssd1 vccd1 vccd1 _09507_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09438_ _16305_/Q _09438_/B vssd1 vssd1 vccd1 vccd1 _09438_/X sky130_fd_sc_hd__or2_1
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09369_ _09386_/B _09369_/B _09369_/C _09369_/D vssd1 vssd1 vccd1 vccd1 _09369_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_240_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ _12234_/A _11400_/B vssd1 vssd1 vccd1 vccd1 _11400_/X sky130_fd_sc_hd__or2_1
XFILLER_0_227_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12380_ _12380_/A _12380_/B vssd1 vssd1 vccd1 vccd1 _12405_/S sky130_fd_sc_hd__or2_2
XFILLER_0_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_70 hold597/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_81 _15145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11331_ _11622_/A _11331_/B vssd1 vssd1 vccd1 vccd1 _11331_/X sky130_fd_sc_hd__or2_1
XANTENNA_92 hold5946/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14050_ _14443_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14050_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11262_ _11556_/A _11262_/B vssd1 vssd1 vccd1 vccd1 _11262_/X sky130_fd_sc_hd__or2_1
XFILLER_0_238_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13001_ hold4760/X _13000_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _13001_/X sky130_fd_sc_hd__mux2_1
Xhold5060 _16817_/Q vssd1 vssd1 vccd1 vccd1 hold5060/X sky130_fd_sc_hd__dlygate4sd3_1
X_10213_ hold3907/X _10631_/B _10212_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10213_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5071 _10999_/X vssd1 vssd1 vccd1 vccd1 _16823_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5082 _16981_/Q vssd1 vssd1 vccd1 vccd1 hold5082/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5093 _10234_/X vssd1 vssd1 vccd1 vccd1 _16568_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11193_ hold4531/X _11103_/A _11192_/X vssd1 vssd1 vccd1 vccd1 _11193_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4370 _17116_/Q vssd1 vssd1 vccd1 vccd1 hold4370/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10144_ hold3999/X _10649_/B _10143_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10144_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4381 _16727_/Q vssd1 vssd1 vccd1 vccd1 hold4381/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4392 _11791_/Y vssd1 vssd1 vccd1 vccd1 _17087_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3680 _16471_/Q vssd1 vssd1 vccd1 vccd1 hold3680/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17740_ _17740_/CLK _17740_/D vssd1 vssd1 vccd1 vccd1 _17740_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3691 _10369_/X vssd1 vssd1 vccd1 vccd1 _16613_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10075_ _10603_/A _10075_/B vssd1 vssd1 vccd1 vccd1 _16515_/D sky130_fd_sc_hd__nor2_1
X_14952_ _14952_/A _14952_/B vssd1 vssd1 vccd1 vccd1 _14952_/Y sky130_fd_sc_hd__nand2_1
XTAP_5864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2990 _14061_/X vssd1 vssd1 vccd1 vccd1 _17835_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13903_ _13903_/A _13903_/B vssd1 vssd1 vccd1 vccd1 _17759_/D sky130_fd_sc_hd__and2_1
X_17671_ _17703_/CLK _17671_/D vssd1 vssd1 vccd1 vccd1 _17671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14883_ hold1060/X hold332/X _14882_/Y _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14883_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16622_ _18180_/CLK _16622_/D vssd1 vssd1 vccd1 vccd1 _16622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13834_ _13864_/A _13834_/B vssd1 vssd1 vccd1 vccd1 _13834_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16553_ _18206_/CLK _16553_/D vssd1 vssd1 vccd1 vccd1 _16553_/Q sky130_fd_sc_hd__dfxtp_1
X_13765_ hold5438/X _13883_/B _13764_/X _13765_/C1 vssd1 vssd1 vccd1 vccd1 _13765_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10977_ _11649_/A _10977_/B vssd1 vssd1 vccd1 vccd1 _10977_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15504_ _15506_/A hold424/X vssd1 vssd1 vccd1 vccd1 hold425/A sky130_fd_sc_hd__and2_1
XFILLER_0_127_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12716_ hold3894/X _12715_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12717_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16484_ _18399_/CLK _16484_/D vssd1 vssd1 vccd1 vccd1 _16484_/Q sky130_fd_sc_hd__dfxtp_1
X_13696_ hold5605/X _13877_/B _13695_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13696_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18223_ _18223_/CLK _18223_/D vssd1 vssd1 vccd1 vccd1 _18223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15435_ hold154/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15435_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12647_ hold3343/X _12646_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12647_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_150_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15366_ _17340_/Q _15486_/B1 _15485_/B1 hold264/X vssd1 vssd1 vccd1 vccd1 _15366_/X
+ sky130_fd_sc_hd__a22o_1
X_18154_ _18154_/CLK _18154_/D vssd1 vssd1 vccd1 vccd1 _18154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12578_ hold3399/X _12577_/X _12971_/S vssd1 vssd1 vccd1 vccd1 _12579_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17105_ _17900_/CLK _17105_/D vssd1 vssd1 vccd1 vccd1 _17105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14317_ hold1875/X _14333_/A2 _14316_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _14317_/X
+ sky130_fd_sc_hd__o211a_1
X_11529_ _12210_/A _11529_/B vssd1 vssd1 vccd1 vccd1 _11529_/X sky130_fd_sc_hd__or2_1
X_15297_ hold571/X _15487_/A2 _15484_/B1 hold695/X _15296_/X vssd1 vssd1 vccd1 vccd1
+ _15302_/B sky130_fd_sc_hd__a221o_1
X_18085_ _18213_/CLK _18085_/D vssd1 vssd1 vccd1 vccd1 _18085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold307 hold307/A vssd1 vssd1 vccd1 vccd1 hold307/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold318 hold43/X vssd1 vssd1 vccd1 vccd1 input28/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14248_ _14517_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14248_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold329 hold404/X vssd1 vssd1 vccd1 vccd1 hold405/A sky130_fd_sc_hd__buf_4
X_17036_ _17884_/CLK _17036_/D vssd1 vssd1 vccd1 vccd1 _17036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14179_ hold1321/X _14202_/B _14178_/X _14462_/C1 vssd1 vssd1 vccd1 vccd1 _14179_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout809 fanout816/X vssd1 vssd1 vccd1 vccd1 _15070_/A sky130_fd_sc_hd__buf_4
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_225_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08740_ _15491_/A _08740_/B vssd1 vssd1 vccd1 vccd1 _15990_/D sky130_fd_sc_hd__and2_1
Xhold1007 hold520/X vssd1 vssd1 vccd1 vccd1 hold1007/X sky130_fd_sc_hd__buf_4
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1018 _14907_/X vssd1 vssd1 vccd1 vccd1 _18241_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17938_ _17997_/CLK _17938_/D vssd1 vssd1 vccd1 vccd1 _17938_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1029 _18132_/Q vssd1 vssd1 vccd1 vccd1 hold1029/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08671_ hold684/X hold718/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold719/A sky130_fd_sc_hd__mux2_1
XFILLER_0_212_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17869_ _17901_/CLK _17869_/D vssd1 vssd1 vccd1 vccd1 _17869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09223_ hold1929/X _09214_/B _09222_/X _12837_/A vssd1 vssd1 vccd1 vccd1 _09223_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09154_ _15537_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09154_/X sky130_fd_sc_hd__or2_1
XFILLER_0_185_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08105_ _15494_/A _08105_/B vssd1 vssd1 vccd1 vccd1 _15691_/D sky130_fd_sc_hd__and2_1
XFILLER_0_86_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09085_ hold3070/X _09102_/B _09084_/X _12984_/A vssd1 vssd1 vccd1 vccd1 _09085_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08036_ hold2173/X _08033_/B _08035_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _08036_/X
+ sky130_fd_sc_hd__o211a_1
Xhold830 hold830/A vssd1 vssd1 vccd1 vccd1 hold830/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold841 hold990/X vssd1 vssd1 vccd1 vccd1 hold991/A sky130_fd_sc_hd__buf_6
XFILLER_0_229_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold852 hold852/A vssd1 vssd1 vccd1 vccd1 hold852/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold863 hold863/A vssd1 vssd1 vccd1 vccd1 hold863/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 hold874/A vssd1 vssd1 vccd1 vccd1 hold874/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold885 hold885/A vssd1 vssd1 vccd1 vccd1 hold885/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 hold896/A vssd1 vssd1 vccd1 vccd1 hold896/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_239_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_265_wb_clk_i clkbuf_6_56_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17929_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09987_ _09987_/A _09987_/B vssd1 vssd1 vccd1 vccd1 _09987_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2220 _18343_/Q vssd1 vssd1 vccd1 vccd1 hold2220/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2231 _18078_/Q vssd1 vssd1 vccd1 vccd1 hold2231/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08938_ _15344_/A hold717/X vssd1 vssd1 vccd1 vccd1 _16086_/D sky130_fd_sc_hd__and2_1
XTAP_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2242 _14568_/X vssd1 vssd1 vccd1 vccd1 hold2242/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2253 _07811_/X vssd1 vssd1 vccd1 vccd1 hold2253/X sky130_fd_sc_hd__buf_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2264 hold2270/X vssd1 vssd1 vccd1 vccd1 hold2264/X sky130_fd_sc_hd__clkbuf_2
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1530 _16311_/Q vssd1 vssd1 vccd1 vccd1 _09456_/B sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2275 _07807_/X vssd1 vssd1 vccd1 vccd1 hold2275/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1541 hold1541/A vssd1 vssd1 vccd1 vccd1 input65/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2286 _08430_/X vssd1 vssd1 vccd1 vccd1 _15845_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08869_ _12380_/B _12445_/B vssd1 vssd1 vccd1 vccd1 _08910_/S sky130_fd_sc_hd__or2_2
Xhold2297 _18300_/Q vssd1 vssd1 vccd1 vccd1 hold2297/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1552 _16274_/Q vssd1 vssd1 vccd1 vccd1 hold1552/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1563 _07887_/X vssd1 vssd1 vccd1 vccd1 _15587_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1574 _15588_/Q vssd1 vssd1 vccd1 vccd1 hold1574/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10900_ hold4911/X _11186_/B _10899_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _10900_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1585 _15790_/Q vssd1 vssd1 vccd1 vccd1 hold1585/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11880_ _12159_/A _11880_/B vssd1 vssd1 vccd1 vccd1 _11880_/X sky130_fd_sc_hd__or2_1
Xhold1596 _17859_/Q vssd1 vssd1 vccd1 vccd1 hold1596/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10831_ hold5448/X _11213_/B _10830_/X _14342_/A vssd1 vssd1 vccd1 vccd1 _10831_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13550_ hold1066/X hold5231/X _13871_/C vssd1 vssd1 vccd1 vccd1 _13551_/B sky130_fd_sc_hd__mux2_1
X_10762_ hold4095/X _11144_/B _10761_/X _14364_/A vssd1 vssd1 vccd1 vccd1 _10762_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12501_ hold82/A _12509_/A2 _12501_/A3 _12500_/X _15364_/A vssd1 vssd1 vccd1 vccd1
+ hold21/A sky130_fd_sc_hd__o311a_1
XFILLER_0_183_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13481_ hold1564/X _17614_/Q _13481_/S vssd1 vssd1 vccd1 vccd1 _13482_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_48_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10693_ hold4575/X _11171_/B _10692_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _10693_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15220_ hold1165/X _15219_/B _15219_/Y _15030_/A vssd1 vssd1 vccd1 vccd1 _15220_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12432_ _15324_/A _12432_/B vssd1 vssd1 vccd1 vccd1 _17309_/D sky130_fd_sc_hd__and2_1
XFILLER_0_129_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15151_ _15205_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15151_/X sky130_fd_sc_hd__or2_1
XFILLER_0_152_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12363_ hold5717/X _12267_/A _12362_/X vssd1 vssd1 vccd1 vccd1 _12363_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14102_ hold820/A _14104_/B vssd1 vssd1 vccd1 vccd1 hold709/A sky130_fd_sc_hd__or2_1
XFILLER_0_200_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11314_ hold4097/X _12335_/B _11313_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _11314_/X
+ sky130_fd_sc_hd__o211a_1
X_15082_ hold3171/X hold340/X _15081_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _15082_/X
+ sky130_fd_sc_hd__o211a_1
X_12294_ hold4373/X _12198_/A _12293_/X vssd1 vssd1 vccd1 vccd1 _12294_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_240_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14033_ hold1550/X _14038_/B _14032_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _14033_/X
+ sky130_fd_sc_hd__o211a_1
X_11245_ hold5525/X _11726_/B _11244_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _11245_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11176_ _12331_/A _11176_/B vssd1 vssd1 vccd1 vccd1 _11176_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_38_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10127_ hold2886/X hold3488/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10128_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_175_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15984_ _18308_/CLK _15984_/D vssd1 vssd1 vccd1 vccd1 hold389/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17723_ _17723_/CLK _17723_/D vssd1 vssd1 vccd1 vccd1 _17723_/Q sky130_fd_sc_hd__dfxtp_1
X_14935_ hold1576/X _14946_/B _14934_/X _15146_/C1 vssd1 vssd1 vccd1 vccd1 _14935_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10058_ _16510_/Q _10634_/B _10634_/C vssd1 vssd1 vccd1 vccd1 _10058_/X sky130_fd_sc_hd__and3_1
XFILLER_0_234_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17654_ _17686_/CLK _17654_/D vssd1 vssd1 vccd1 vccd1 _17654_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14866_ _15205_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14866_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16605_ _18227_/CLK _16605_/D vssd1 vssd1 vccd1 vccd1 _16605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13817_ _13817_/A _13817_/B _13817_/C vssd1 vssd1 vccd1 vccd1 _13817_/X sky130_fd_sc_hd__and3_1
XFILLER_0_58_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17585_ _17745_/CLK _17585_/D vssd1 vssd1 vccd1 vccd1 _17585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14797_ hold2920/X _14828_/B _14796_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14797_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_69_wb_clk_i clkbuf_6_19_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16319_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16536_ _17960_/CLK _16536_/D vssd1 vssd1 vccd1 vccd1 _16536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13748_ hold2234/X _17703_/Q _13748_/S vssd1 vssd1 vccd1 vccd1 _13749_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16467_ _18380_/CLK _16467_/D vssd1 vssd1 vccd1 vccd1 _16467_/Q sky130_fd_sc_hd__dfxtp_1
X_13679_ hold1404/X hold5285/X _13865_/C vssd1 vssd1 vccd1 vccd1 _13680_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_214_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18206_ _18206_/CLK _18206_/D vssd1 vssd1 vccd1 vccd1 _18206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15418_ hold560/X _15448_/A2 _09362_/C _17345_/Q vssd1 vssd1 vccd1 vccd1 _15418_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16398_ _18375_/CLK _16398_/D vssd1 vssd1 vccd1 vccd1 _16398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18137_ _18181_/CLK _18137_/D vssd1 vssd1 vccd1 vccd1 _18137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15349_ hold799/X _09365_/B _09392_/C hold500/X _15348_/X vssd1 vssd1 vccd1 vccd1
+ _15352_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_13_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_1360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5807 _16498_/Q vssd1 vssd1 vccd1 vccd1 hold5807/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5818 _09922_/X vssd1 vssd1 vccd1 vccd1 _16464_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5829 _16452_/Q vssd1 vssd1 vccd1 vccd1 hold5829/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 hold334/X vssd1 vssd1 vccd1 vccd1 hold335/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 hold115/A vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__clkbuf_16
Xhold126 hold126/A vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
X_18068_ _18070_/CLK _18068_/D vssd1 vssd1 vccd1 vccd1 _18068_/Q sky130_fd_sc_hd__dfxtp_1
Xhold137 hold137/A vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold148 hold148/A vssd1 vssd1 vccd1 vccd1 hold148/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold159 hold159/A vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ hold4735/X _10004_/B _09909_/X _15042_/A vssd1 vssd1 vccd1 vccd1 _09910_/X
+ sky130_fd_sc_hd__o211a_1
X_17019_ _17771_/CLK _17019_/D vssd1 vssd1 vccd1 vccd1 _17019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout606 _09364_/Y vssd1 vssd1 vccd1 vccd1 _09392_/D sky130_fd_sc_hd__buf_8
X_09841_ hold4711/X _10031_/B _09840_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09841_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout617 _09356_/Y vssd1 vssd1 vccd1 vccd1 _09392_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout628 hold355/X vssd1 vssd1 vccd1 vccd1 _08504_/A sky130_fd_sc_hd__clkbuf_8
Xfanout639 _12849_/A vssd1 vssd1 vccd1 vccd1 _12837_/A sky130_fd_sc_hd__buf_4
XFILLER_0_237_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09772_ hold3660/X _10052_/B _09771_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _09772_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ hold495/X _15983_/Q _08723_/S vssd1 vssd1 vccd1 vccd1 hold496/A sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_213_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_234_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08654_ _15364_/A hold456/X vssd1 vssd1 vccd1 vccd1 _15949_/D sky130_fd_sc_hd__and2_1
XFILLER_0_55_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08585_ _08851_/A _08585_/B vssd1 vssd1 vccd1 vccd1 _15916_/D sky130_fd_sc_hd__and2_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_234_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09206_ _09313_/A _09206_/B vssd1 vssd1 vccd1 vccd1 _09206_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09137_ hold1130/X _09177_/A2 _09136_/X _12855_/A vssd1 vssd1 vccd1 vccd1 _09137_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09068_ hold927/X _09118_/B vssd1 vssd1 vccd1 vccd1 _09068_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_446_wb_clk_i clkbuf_6_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17127_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_103_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08019_ _15533_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08019_/X sky130_fd_sc_hd__or2_1
Xhold660 hold660/A vssd1 vssd1 vccd1 vccd1 hold660/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold671 hold73/X vssd1 vssd1 vccd1 vccd1 input36/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold682 hold682/A vssd1 vssd1 vccd1 vccd1 input30/A sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ hold1799/X _16834_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _11031_/B sky130_fd_sc_hd__mux2_1
Xhold693 hold693/A vssd1 vssd1 vccd1 vccd1 hold693/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2050 _14711_/X vssd1 vssd1 vccd1 vccd1 _18147_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2061 _09117_/X vssd1 vssd1 vccd1 vccd1 _16173_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2072 _14097_/X vssd1 vssd1 vccd1 vccd1 _17853_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _12987_/A _12981_/B vssd1 vssd1 vccd1 vccd1 _17503_/D sky130_fd_sc_hd__and2_1
Xhold2083 _17997_/Q vssd1 vssd1 vccd1 vccd1 hold2083/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_231_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2094 _17931_/Q vssd1 vssd1 vccd1 vccd1 hold2094/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1360 _17936_/Q vssd1 vssd1 vccd1 vccd1 hold1360/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14720_ _14952_/A _14720_/B vssd1 vssd1 vccd1 vccd1 _14720_/Y sky130_fd_sc_hd__nand2_1
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1371 _08271_/X vssd1 vssd1 vccd1 vccd1 _15770_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ hold3702/X _12356_/B _11931_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _11932_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1382 _15624_/Q vssd1 vssd1 vccd1 vccd1 hold1382/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1393 _17857_/Q vssd1 vssd1 vccd1 vccd1 hold1393/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14651_ hold1455/X _14666_/B _14650_/X _15218_/C1 vssd1 vssd1 vccd1 vccd1 _14651_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ hold4011/X _12365_/B _11862_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _11863_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ hold1592/X hold4056/X _11213_/C vssd1 vssd1 vccd1 vccd1 _10815_/B sky130_fd_sc_hd__mux2_1
X_13602_ _13794_/A _13602_/B vssd1 vssd1 vccd1 vccd1 _13602_/X sky130_fd_sc_hd__or2_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17370_ _18013_/CLK _17370_/D vssd1 vssd1 vccd1 vccd1 _17370_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14582_ _15191_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14582_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11794_ _12337_/A _11794_/B vssd1 vssd1 vccd1 vccd1 _11794_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_28_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16321_ _16323_/CLK _16321_/D vssd1 vssd1 vccd1 vccd1 _16321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10745_ hold1420/X hold4278/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10746_/B sky130_fd_sc_hd__mux2_1
X_13533_ _13734_/A _13533_/B vssd1 vssd1 vccd1 vccd1 _13533_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16252_ _17754_/CLK _16252_/D vssd1 vssd1 vccd1 vccd1 hold973/A sky130_fd_sc_hd__dfxtp_1
X_13464_ _13581_/A _13464_/B vssd1 vssd1 vccd1 vccd1 _13464_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10676_ hold2199/X hold3479/X _11162_/C vssd1 vssd1 vccd1 vccd1 _10677_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15203_ _15203_/A _15227_/B vssd1 vssd1 vccd1 vccd1 _15203_/X sky130_fd_sc_hd__or2_1
X_12415_ hold254/X hold540/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12416_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13395_ _13758_/A _13395_/B vssd1 vssd1 vccd1 vccd1 _13395_/X sky130_fd_sc_hd__or2_1
X_16183_ _17468_/CLK _16183_/D vssd1 vssd1 vccd1 vccd1 _16183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15134_ hold2037/X _15165_/B _15133_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _15134_/X
+ sky130_fd_sc_hd__o211a_1
X_12346_ _13888_/A _12346_/B vssd1 vssd1 vccd1 vccd1 _12346_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_187_wb_clk_i clkbuf_6_52_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18346_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_116_wb_clk_i clkbuf_6_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16125_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15065_ _15227_/A hold2536/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15066_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12277_ hold5171/X _12374_/B _12276_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _12277_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14016_ hold933/X _14042_/B vssd1 vssd1 vccd1 vccd1 _14016_/X sky130_fd_sc_hd__or2_1
X_11228_ hold1813/X _16900_/Q _11717_/C vssd1 vssd1 vccd1 vccd1 _11229_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_226_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11159_ _16877_/Q _11162_/B _11162_/C vssd1 vssd1 vccd1 vccd1 _11159_/X sky130_fd_sc_hd__and3_1
XTAP_6181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15967_ _18409_/CLK _15967_/D vssd1 vssd1 vccd1 vccd1 hold608/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17706_ _17738_/CLK _17706_/D vssd1 vssd1 vccd1 vccd1 _17706_/Q sky130_fd_sc_hd__dfxtp_1
X_14918_ _15187_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14918_/X sky130_fd_sc_hd__or2_1
XFILLER_0_188_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_236_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15898_ _17523_/CLK _15898_/D vssd1 vssd1 vccd1 vccd1 hold454/A sky130_fd_sc_hd__dfxtp_1
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17637_ _17733_/CLK _17637_/D vssd1 vssd1 vccd1 vccd1 _17637_/Q sky130_fd_sc_hd__dfxtp_1
X_14849_ hold2051/X hold332/X _14848_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14849_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_231_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08370_ _15539_/A hold1263/X hold115/X vssd1 vssd1 vccd1 vccd1 _08371_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_74_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17568_ _17728_/CLK _17568_/D vssd1 vssd1 vccd1 vccd1 _17568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16519_ _18174_/CLK _16519_/D vssd1 vssd1 vccd1 vccd1 _16519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17499_ _17499_/CLK _17499_/D vssd1 vssd1 vccd1 vccd1 _17499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5604 _13792_/X vssd1 vssd1 vccd1 vccd1 _17717_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5615 _11332_/X vssd1 vssd1 vccd1 vccd1 _16934_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5626 _16874_/Q vssd1 vssd1 vccd1 vccd1 hold5626/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5637 _16997_/Q vssd1 vssd1 vccd1 vccd1 hold5637/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5648 _10783_/X vssd1 vssd1 vccd1 vccd1 _16751_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4903 _17190_/Q vssd1 vssd1 vccd1 vccd1 hold4903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4914 _12154_/X vssd1 vssd1 vccd1 vccd1 _17208_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5659 _16967_/Q vssd1 vssd1 vccd1 vccd1 hold5659/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4925 _16852_/Q vssd1 vssd1 vccd1 vccd1 hold4925/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_223_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4936 _10873_/X vssd1 vssd1 vccd1 vccd1 _16781_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4947 _17014_/Q vssd1 vssd1 vccd1 vccd1 hold4947/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4958 _11080_/X vssd1 vssd1 vccd1 vccd1 _16850_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4969 _12127_/X vssd1 vssd1 vccd1 vccd1 _17199_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout403 _14393_/Y vssd1 vssd1 vccd1 vccd1 _14446_/A2 sky130_fd_sc_hd__buf_8
Xfanout414 _14162_/Y vssd1 vssd1 vccd1 vccd1 _14202_/B sky130_fd_sc_hd__buf_6
XFILLER_0_39_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout425 _13946_/Y vssd1 vssd1 vccd1 vccd1 _13995_/A2 sky130_fd_sc_hd__buf_8
Xfanout436 _13721_/S vssd1 vssd1 vccd1 vccd1 _13817_/C sky130_fd_sc_hd__buf_6
XFILLER_0_195_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09824_ hold2950/X hold4891/X _11171_/C vssd1 vssd1 vccd1 vccd1 _09825_/B sky130_fd_sc_hd__mux2_1
Xfanout447 _11717_/C vssd1 vssd1 vccd1 vccd1 _12299_/C sky130_fd_sc_hd__clkbuf_8
Xfanout458 fanout485/X vssd1 vssd1 vccd1 vccd1 _11168_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout469 fanout485/X vssd1 vssd1 vccd1 vccd1 _13877_/C sky130_fd_sc_hd__clkbuf_4
X_09755_ hold1941/X hold4687/X _10031_/C vssd1 vssd1 vccd1 vccd1 _09756_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_226_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08706_ _15254_/A _08706_/B vssd1 vssd1 vccd1 vccd1 _15974_/D sky130_fd_sc_hd__and2_1
XFILLER_0_119_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09686_ hold2856/X hold3662/X _10985_/S vssd1 vssd1 vccd1 vccd1 _09687_/B sky130_fd_sc_hd__mux2_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ hold215/X hold769/X _08657_/S vssd1 vssd1 vccd1 vccd1 _08638_/B sky130_fd_sc_hd__mux2_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_234_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08568_ hold245/X hold547/X _08592_/S vssd1 vssd1 vccd1 vccd1 _08569_/B sky130_fd_sc_hd__mux2_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08499_ hold1188/X _08486_/B _08498_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _08499_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10530_ _10530_/A _10530_/B vssd1 vssd1 vccd1 vccd1 _10530_/X sky130_fd_sc_hd__or2_1
XFILLER_0_147_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10461_ _10986_/A _10461_/B vssd1 vssd1 vccd1 vccd1 _10461_/X sky130_fd_sc_hd__or2_1
X_12200_ hold1602/X hold4797/X _13811_/C vssd1 vssd1 vccd1 vccd1 _12201_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_280_wb_clk_i clkbuf_6_50_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18208_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13180_ hold4341/X _13179_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13180_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10392_ _10524_/A _10392_/B vssd1 vssd1 vccd1 vccd1 _10392_/X sky130_fd_sc_hd__or2_1
XFILLER_0_206_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12131_ hold1354/X hold5430/X _12362_/C vssd1 vssd1 vccd1 vccd1 _12132_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_102_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12062_ hold1590/X _17178_/Q _13463_/S vssd1 vssd1 vccd1 vccd1 _12063_/B sky130_fd_sc_hd__mux2_1
Xhold490 hold490/A vssd1 vssd1 vccd1 vccd1 hold490/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11013_ _11109_/A _11013_/B vssd1 vssd1 vccd1 vccd1 _11013_/X sky130_fd_sc_hd__or2_1
XFILLER_0_99_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16870_ _17913_/CLK _16870_/D vssd1 vssd1 vccd1 vccd1 _16870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_216_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15821_ _17732_/CLK hold117/X vssd1 vssd1 vccd1 vccd1 _15821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _17745_/CLK _15752_/D vssd1 vssd1 vccd1 vccd1 _15752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12964_ hold2002/X _17499_/Q _12970_/S vssd1 vssd1 vccd1 vccd1 _12964_/X sky130_fd_sc_hd__mux2_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1190 la_data_in[0] vssd1 vssd1 vccd1 vccd1 hold925/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14703_ hold2659/X _14718_/B _14702_/X _14769_/C1 vssd1 vssd1 vccd1 vccd1 _14703_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ hold2705/X _17129_/Q _12299_/C vssd1 vssd1 vccd1 vccd1 _11916_/B sky130_fd_sc_hd__mux2_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ _17281_/CLK _15683_/D vssd1 vssd1 vccd1 vccd1 _15683_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ hold3021/X _17476_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12895_/X sky130_fd_sc_hd__mux2_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17422_ _17690_/CLK _17422_/D vssd1 vssd1 vccd1 vccd1 _17422_/Q sky130_fd_sc_hd__dfxtp_1
X_14634_ _15189_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14634_/X sky130_fd_sc_hd__or2_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ hold941/X hold4290/X _12332_/C vssd1 vssd1 vccd1 vccd1 _11847_/B sky130_fd_sc_hd__mux2_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17353_ _17516_/CLK _17353_/D vssd1 vssd1 vccd1 vccd1 _17353_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565_ _15189_/A _14557_/Y hold2280/X _15218_/C1 vssd1 vssd1 vccd1 vccd1 _14565_/X
+ sky130_fd_sc_hd__o211a_1
X_11777_ _17083_/Q _12317_/B _12317_/C vssd1 vssd1 vccd1 vccd1 _11777_/X sky130_fd_sc_hd__and3_1
XFILLER_0_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16304_ _18408_/CLK _16304_/D vssd1 vssd1 vccd1 vccd1 _16304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13516_ hold5787/X _13808_/B _13515_/X _12738_/A vssd1 vssd1 vccd1 vccd1 _13516_/X
+ sky130_fd_sc_hd__o211a_1
X_10728_ _11661_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _10728_/X sky130_fd_sc_hd__or2_1
X_17284_ _17284_/CLK _17284_/D vssd1 vssd1 vccd1 vccd1 hold726/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_368_wb_clk_i clkbuf_6_34_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17707_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14496_ hold878/X _14487_/B _14495_/X _15506_/A vssd1 vssd1 vccd1 vccd1 hold879/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16235_ _17430_/CLK _16235_/D vssd1 vssd1 vccd1 vccd1 _16235_/Q sky130_fd_sc_hd__dfxtp_1
X_13447_ hold4559/X _13829_/B _13446_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13447_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10659_ _11637_/A _10659_/B vssd1 vssd1 vccd1 vccd1 _10659_/X sky130_fd_sc_hd__or2_1
XFILLER_0_113_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16166_ _17513_/CLK _16166_/D vssd1 vssd1 vccd1 vccd1 _16166_/Q sky130_fd_sc_hd__dfxtp_1
X_13378_ hold5519/X _13847_/B _13377_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13378_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15117_ _15225_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15117_/X sky130_fd_sc_hd__or2_1
X_12329_ _17267_/Q _12329_/B _12329_/C vssd1 vssd1 vccd1 vccd1 _12329_/X sky130_fd_sc_hd__and3_1
XFILLER_0_220_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16097_ _16129_/CLK _16097_/D vssd1 vssd1 vccd1 vccd1 _16097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3509 _11145_/Y vssd1 vssd1 vccd1 vccd1 _11146_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15048_ _15048_/A _15048_/B vssd1 vssd1 vccd1 vccd1 _18309_/D sky130_fd_sc_hd__and2_1
XFILLER_0_142_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2808 _08292_/X vssd1 vssd1 vccd1 vccd1 _15779_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2819 _18371_/Q vssd1 vssd1 vccd1 vccd1 hold2819/X sky130_fd_sc_hd__dlygate4sd3_1
X_07870_ hold2402/X _07869_/B _07869_/Y _08153_/A vssd1 vssd1 vccd1 vccd1 _07870_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_218_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16999_ _17882_/CLK _16999_/D vssd1 vssd1 vccd1 vccd1 _16999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09540_ _09933_/A _09540_/B vssd1 vssd1 vccd1 vccd1 _09540_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_84_wb_clk_i clkbuf_6_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17493_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_183_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_wb_clk_i clkbuf_6_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17471_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_231_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09471_ hold733/X _09471_/B vssd1 vssd1 vccd1 vccd1 _09473_/C sky130_fd_sc_hd__or2_1
Xclkbuf_6_41_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_41_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_176_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08422_ hold1548/X _08442_/A2 _08421_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _08422_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08353_ _12750_/A _08353_/B vssd1 vssd1 vccd1 vccd1 _15808_/D sky130_fd_sc_hd__and2_1
XFILLER_0_164_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08284_ _08504_/A hold338/X vssd1 vssd1 vccd1 vccd1 _08335_/B sky130_fd_sc_hd__or2_4
XFILLER_0_15_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6102 la_data_in[30] vssd1 vssd1 vccd1 vccd1 hold350/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold6113 _16323_/Q vssd1 vssd1 vccd1 vccd1 hold6113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6124 _16518_/Q vssd1 vssd1 vccd1 vccd1 hold6124/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6135 la_data_in[7] vssd1 vssd1 vccd1 vccd1 hold929/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5401 _11602_/X vssd1 vssd1 vccd1 vccd1 _17024_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5412 _17715_/Q vssd1 vssd1 vccd1 vccd1 hold5412/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5423 _10534_/X vssd1 vssd1 vccd1 vccd1 _16668_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5434 _16938_/Q vssd1 vssd1 vccd1 vccd1 hold5434/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4700 _11905_/X vssd1 vssd1 vccd1 vccd1 _17125_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5445 _11542_/X vssd1 vssd1 vccd1 vccd1 _17004_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4711 _16469_/Q vssd1 vssd1 vccd1 vccd1 hold4711/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5456 _17230_/Q vssd1 vssd1 vccd1 vccd1 hold5456/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5467 _13393_/X vssd1 vssd1 vccd1 vccd1 _17584_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4722 _17107_/Q vssd1 vssd1 vccd1 vccd1 hold4722/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4733 _17729_/Q vssd1 vssd1 vccd1 vccd1 hold4733/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5478 _17735_/Q vssd1 vssd1 vccd1 vccd1 hold5478/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4744 _13798_/X vssd1 vssd1 vccd1 vccd1 _17719_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5489 _11074_/X vssd1 vssd1 vccd1 vccd1 _16848_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4755 _09937_/X vssd1 vssd1 vccd1 vccd1 _16469_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4766 _16899_/Q vssd1 vssd1 vccd1 vccd1 hold4766/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout200 fanout210/X vssd1 vssd1 vccd1 vccd1 _11786_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4777 _16362_/Q vssd1 vssd1 vccd1 vccd1 hold4777/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout211 _11144_/B vssd1 vssd1 vccd1 vccd1 _11153_/B sky130_fd_sc_hd__buf_4
Xhold4788 _11920_/X vssd1 vssd1 vccd1 vccd1 _17130_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout222 _09494_/X vssd1 vssd1 vccd1 vccd1 _10013_/B sky130_fd_sc_hd__clkbuf_8
Xfanout233 _10634_/B vssd1 vssd1 vccd1 vccd1 _10604_/B sky130_fd_sc_hd__clkbuf_4
Xhold4799 _16741_/Q vssd1 vssd1 vccd1 vccd1 hold4799/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout244 _10637_/B vssd1 vssd1 vccd1 vccd1 _10619_/B sky130_fd_sc_hd__buf_4
Xfanout255 _13794_/A vssd1 vssd1 vccd1 vccd1 _13737_/A sky130_fd_sc_hd__buf_4
XFILLER_0_214_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout266 _11553_/A vssd1 vssd1 vccd1 vccd1 _12285_/A sky130_fd_sc_hd__buf_4
XFILLER_0_201_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09807_ _11067_/A _09807_/B vssd1 vssd1 vccd1 vccd1 _09807_/X sky130_fd_sc_hd__or2_1
Xfanout277 _12159_/A vssd1 vssd1 vccd1 vccd1 _12255_/A sky130_fd_sc_hd__buf_4
Xfanout288 fanout299/X vssd1 vssd1 vccd1 vccd1 _11667_/A sky130_fd_sc_hd__clkbuf_4
Xfanout299 wire337/A vssd1 vssd1 vccd1 vccd1 fanout299/X sky130_fd_sc_hd__buf_12
X_07999_ hold911/X _08045_/B vssd1 vssd1 vccd1 vccd1 _07999_/X sky130_fd_sc_hd__or2_1
XFILLER_0_241_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09738_ _09948_/A _09738_/B vssd1 vssd1 vccd1 vccd1 _09738_/X sky130_fd_sc_hd__or2_1
XFILLER_0_213_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09669_ _09957_/A _09669_/B vssd1 vssd1 vccd1 vccd1 _09669_/X sky130_fd_sc_hd__or2_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _12174_/A _11700_/B vssd1 vssd1 vccd1 vccd1 _11700_/X sky130_fd_sc_hd__or2_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12680_ hold3379/X _12679_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12681_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_194_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11631_ _11631_/A _11631_/B vssd1 vssd1 vccd1 vccd1 _11631_/X sky130_fd_sc_hd__or2_1
XFILLER_0_155_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14350_ _14350_/A _14350_/B vssd1 vssd1 vccd1 vccd1 _17974_/D sky130_fd_sc_hd__and2_1
XFILLER_0_68_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11562_ _11658_/A _11562_/B vssd1 vssd1 vccd1 vccd1 _11562_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_461_wb_clk_i clkbuf_6_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17753_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10513_ hold3765/X _10631_/B _10512_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10513_/X
+ sky130_fd_sc_hd__o211a_1
X_13301_ _13300_/X hold4245/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13301_/X sky130_fd_sc_hd__mux2_1
X_14281_ hold2777/X _14272_/B _14280_/X _14526_/C1 vssd1 vssd1 vccd1 vccd1 _14281_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11493_ _12219_/A _11493_/B vssd1 vssd1 vccd1 vccd1 _11493_/X sky130_fd_sc_hd__or2_1
X_13232_ _13225_/X _13231_/X _13296_/B1 vssd1 vssd1 vccd1 vccd1 _17547_/D sky130_fd_sc_hd__o21a_1
X_16020_ _16120_/CLK _16020_/D vssd1 vssd1 vccd1 vccd1 hold431/A sky130_fd_sc_hd__dfxtp_1
X_10444_ hold3878/X _10598_/B _10443_/X _14895_/C1 vssd1 vssd1 vccd1 vccd1 _10444_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13163_ _13162_/X hold4430/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13163_/X sky130_fd_sc_hd__mux2_1
X_10375_ hold3775/X _10589_/B _10374_/X _14769_/C1 vssd1 vssd1 vccd1 vccd1 _10375_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12114_ _12210_/A _12114_/B vssd1 vssd1 vccd1 vccd1 _12114_/X sky130_fd_sc_hd__or2_1
X_13094_ _13094_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13094_/X sky130_fd_sc_hd__or2_1
X_17971_ _17971_/CLK _17971_/D vssd1 vssd1 vccd1 vccd1 _17971_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5990 _16902_/Q vssd1 vssd1 vccd1 vccd1 hold5990/X sky130_fd_sc_hd__dlygate4sd3_1
X_12045_ _12255_/A _12045_/B vssd1 vssd1 vccd1 vccd1 _12045_/X sky130_fd_sc_hd__or2_1
X_16922_ _17834_/CLK _16922_/D vssd1 vssd1 vccd1 vccd1 _16922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_236_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_217_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16853_ _18056_/CLK _16853_/D vssd1 vssd1 vccd1 vccd1 _16853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15804_ _17620_/CLK _15804_/D vssd1 vssd1 vccd1 vccd1 _15804_/Q sky130_fd_sc_hd__dfxtp_1
X_16784_ _18019_/CLK _16784_/D vssd1 vssd1 vccd1 vccd1 _16784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13996_ _14443_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13996_/X sky130_fd_sc_hd__or2_1
X_15735_ _17740_/CLK _15735_/D vssd1 vssd1 vccd1 vccd1 _15735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12947_ hold4441/X _12946_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12948_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18454_ _18455_/CLK _18454_/D vssd1 vssd1 vccd1 vccd1 _18454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15666_ _17222_/CLK _15666_/D vssd1 vssd1 vccd1 vccd1 _15666_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ hold3361/X _12877_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12879_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_185_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17405_ _18457_/CLK _17405_/D vssd1 vssd1 vccd1 vccd1 _17405_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ hold2141/X _14612_/B _14616_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14617_/X
+ sky130_fd_sc_hd__o211a_1
X_18385_ _18385_/CLK _18385_/D vssd1 vssd1 vccd1 vccd1 _18385_/Q sky130_fd_sc_hd__dfxtp_1
X_11829_ _13797_/A _11829_/B vssd1 vssd1 vccd1 vccd1 _11829_/X sky130_fd_sc_hd__or2_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15597_ _17277_/CLK _15597_/D vssd1 vssd1 vccd1 vccd1 _15597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17336_ _17336_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 _17336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14548_ hold2546/X _14541_/B _14547_/X _14346_/A vssd1 vssd1 vccd1 vccd1 _14548_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_131_wb_clk_i clkbuf_6_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17322_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_181_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17267_ _17901_/CLK _17267_/D vssd1 vssd1 vccd1 vccd1 _17267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14479_ _14604_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14479_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16218_ _18443_/CLK _16218_/D vssd1 vssd1 vccd1 vccd1 _16218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17198_ _17900_/CLK _17198_/D vssd1 vssd1 vccd1 vccd1 _17198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4007 _16685_/Q vssd1 vssd1 vccd1 vccd1 hold4007/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16149_ _17486_/CLK _16149_/D vssd1 vssd1 vccd1 vccd1 _16149_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4018 _16944_/Q vssd1 vssd1 vccd1 vccd1 hold4018/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4029 _12836_/X vssd1 vssd1 vccd1 vccd1 _12837_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3306 _17468_/Q vssd1 vssd1 vccd1 vccd1 hold3306/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3317 _12896_/X vssd1 vssd1 vccd1 vccd1 _12897_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3328 _16567_/Q vssd1 vssd1 vccd1 vccd1 hold3328/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ hold245/X _16103_/Q _08997_/S vssd1 vssd1 vccd1 vccd1 hold246/A sky130_fd_sc_hd__mux2_1
Xhold3339 _16623_/Q vssd1 vssd1 vccd1 vccd1 hold3339/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2605 _18341_/Q vssd1 vssd1 vccd1 vccd1 hold2605/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2616 _15573_/Q vssd1 vssd1 vccd1 vccd1 hold2616/X sky130_fd_sc_hd__dlygate4sd3_1
X_07922_ _15545_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _07922_/Y sky130_fd_sc_hd__nand2_1
Xhold19 hold79/X vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2627 _17785_/Q vssd1 vssd1 vccd1 vccd1 hold2627/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2638 _14673_/X vssd1 vssd1 vccd1 vccd1 _18129_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1904 _15142_/X vssd1 vssd1 vccd1 vccd1 _18354_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2649 _07975_/X vssd1 vssd1 vccd1 vccd1 _15630_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1915 _17938_/Q vssd1 vssd1 vccd1 vccd1 hold1915/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07853_ _15531_/A _07871_/B vssd1 vssd1 vccd1 vccd1 _07853_/X sky130_fd_sc_hd__or2_1
Xhold1926 _14857_/X vssd1 vssd1 vccd1 vccd1 _18217_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_223_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1937 _18456_/Q vssd1 vssd1 vccd1 vccd1 hold1937/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1948 _14575_/X vssd1 vssd1 vccd1 vccd1 _18081_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1959 _14969_/X vssd1 vssd1 vccd1 vccd1 _18270_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07784_ _07784_/A vssd1 vssd1 vccd1 vccd1 _14556_/A sky130_fd_sc_hd__inv_2
XFILLER_0_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09523_ hold3564/X _10025_/B _09522_/X _15473_/A vssd1 vssd1 vccd1 vccd1 _09523_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_1351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09454_ _09455_/B _09478_/B _09454_/C vssd1 vssd1 vccd1 vccd1 _16311_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_176_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08405_ _15519_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08405_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_219_wb_clk_i clkbuf_6_61_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18177_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09385_ hold5941/A _09342_/B _09342_/Y _09384_/X _15314_/A vssd1 vssd1 vccd1 vccd1
+ _09385_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_136_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08336_ hold1054/X _08336_/A2 _08335_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _08336_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_188_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08267_ hold2406/X _08268_/B _08266_/Y _09272_/A vssd1 vssd1 vccd1 vccd1 _08267_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08198_ hold1307/X _08213_/B _08197_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _08198_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5220 _11011_/X vssd1 vssd1 vccd1 vccd1 _16827_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_1356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5231 _17637_/Q vssd1 vssd1 vccd1 vccd1 hold5231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5242 _10948_/X vssd1 vssd1 vccd1 vccd1 _16806_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5253 _17041_/Q vssd1 vssd1 vccd1 vccd1 hold5253/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5264 _13417_/X vssd1 vssd1 vccd1 vccd1 _17592_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4530 _17485_/Q vssd1 vssd1 vccd1 vccd1 hold4530/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5275 _17283_/Q vssd1 vssd1 vccd1 vccd1 hold5275/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10160_ hold2141/X hold3459/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10161_/B sky130_fd_sc_hd__mux2_1
Xhold5286 _13585_/X vssd1 vssd1 vccd1 vccd1 _17648_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4541 _17666_/Q vssd1 vssd1 vccd1 vccd1 hold4541/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4552 _17360_/Q vssd1 vssd1 vccd1 vccd1 hold4552/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5297 _16708_/Q vssd1 vssd1 vccd1 vccd1 hold5297/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4563 _17236_/Q vssd1 vssd1 vccd1 vccd1 hold4563/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4574 _10261_/X vssd1 vssd1 vccd1 vccd1 _16577_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3840 _16563_/Q vssd1 vssd1 vccd1 vccd1 hold3840/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4585 _17181_/Q vssd1 vssd1 vccd1 vccd1 hold4585/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10091_ hold2241/X _16521_/Q _10475_/S vssd1 vssd1 vccd1 vccd1 _10092_/B sky130_fd_sc_hd__mux2_1
Xhold3851 _10855_/X vssd1 vssd1 vccd1 vccd1 _16775_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4596 _17156_/Q vssd1 vssd1 vccd1 vccd1 hold4596/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3862 _16683_/Q vssd1 vssd1 vccd1 vccd1 hold3862/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3873 _10663_/X vssd1 vssd1 vccd1 vccd1 _16711_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_238_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3884 _16588_/Q vssd1 vssd1 vccd1 vccd1 hold3884/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3895 _16675_/Q vssd1 vssd1 vccd1 vccd1 hold3895/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_236_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13850_ _17737_/Q _13880_/B _13880_/C vssd1 vssd1 vccd1 vccd1 _13850_/X sky130_fd_sc_hd__and3_1
XFILLER_0_92_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_230_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12801_ _12804_/A _12801_/B vssd1 vssd1 vccd1 vccd1 _17443_/D sky130_fd_sc_hd__and2_1
XFILLER_0_199_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10993_ hold3980/X _10616_/B _10992_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _10993_/X
+ sky130_fd_sc_hd__o211a_1
X_13781_ hold2398/X hold5555/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13782_/B sky130_fd_sc_hd__mux2_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15520_ hold1087/X _15560_/A2 _15519_/X _12873_/A vssd1 vssd1 vccd1 vccd1 _15520_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _12753_/A _12732_/B vssd1 vssd1 vccd1 vccd1 _17420_/D sky130_fd_sc_hd__and2_1
XFILLER_0_167_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15451_ hold410/X _09392_/D _15484_/B1 hold587/X _15446_/X vssd1 vssd1 vccd1 vccd1
+ _15452_/D sky130_fd_sc_hd__a221o_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _12873_/A _12663_/B vssd1 vssd1 vccd1 vccd1 _17397_/D sky130_fd_sc_hd__and2_1
XFILLER_0_195_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ hold3169/X _14446_/A2 _14401_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _14402_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18170_ _18170_/CLK _18170_/D vssd1 vssd1 vccd1 vccd1 _18170_/Q sky130_fd_sc_hd__dfxtp_1
X_11614_ hold5199/X _12317_/B _11613_/X _14211_/C1 vssd1 vssd1 vccd1 vccd1 _11614_/X
+ sky130_fd_sc_hd__o211a_1
X_15382_ _15480_/A _15382_/B _15382_/C _15382_/D vssd1 vssd1 vccd1 vccd1 _15382_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_154_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12594_ _12597_/A _12594_/B vssd1 vssd1 vccd1 vccd1 _17374_/D sky130_fd_sc_hd__and2_1
XFILLER_0_136_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17121_ _17153_/CLK _17121_/D vssd1 vssd1 vccd1 vccd1 _17121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14333_ hold1448/X _14333_/A2 _14332_/X _14372_/A vssd1 vssd1 vccd1 vccd1 _14333_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11545_ hold5577/X _11744_/B _11544_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _11545_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17052_ _17900_/CLK _17052_/D vssd1 vssd1 vccd1 vccd1 _17052_/Q sky130_fd_sc_hd__dfxtp_1
X_14264_ _14604_/A _14282_/B vssd1 vssd1 vccd1 vccd1 _14264_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11476_ hold4947/X _11195_/B _11475_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _11476_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16003_ _16086_/CLK _16003_/D vssd1 vssd1 vccd1 vccd1 hold343/A sky130_fd_sc_hd__dfxtp_1
X_13215_ _13311_/A1 _13213_/X _13214_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13215_/X
+ sky130_fd_sc_hd__o211a_1
X_10427_ hold1978/X _16633_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10428_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14195_ hold1484/X _14198_/B _14194_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _14195_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10358_ hold2836/X _16610_/Q _10646_/C vssd1 vssd1 vccd1 vccd1 _10359_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13146_ _17569_/Q _17103_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13146_/X sky130_fd_sc_hd__mux2_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13077_ _13076_/X hold3893/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13077_/X sky130_fd_sc_hd__mux2_1
X_17954_ _17985_/CLK _17954_/D vssd1 vssd1 vccd1 vccd1 _17954_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ hold2679/X hold3240/X _10385_/S vssd1 vssd1 vccd1 vccd1 _10290_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12028_ hold4061/X _12323_/B _12027_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _12028_/X
+ sky130_fd_sc_hd__o211a_1
X_16905_ _18432_/CLK _16905_/D vssd1 vssd1 vccd1 vccd1 _16905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17885_ _17885_/CLK _17885_/D vssd1 vssd1 vccd1 vccd1 _17885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16836_ _18039_/CLK _16836_/D vssd1 vssd1 vccd1 vccd1 _16836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_232_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_232_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16767_ _18194_/CLK _16767_/D vssd1 vssd1 vccd1 vccd1 _16767_/Q sky130_fd_sc_hd__dfxtp_1
X_13979_ hold2131/X _13986_/B _13978_/X _14462_/C1 vssd1 vssd1 vccd1 vccd1 _13979_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_221_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15718_ _17093_/CLK _15718_/D vssd1 vssd1 vccd1 vccd1 _15718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_383_wb_clk_i clkbuf_6_33_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17202_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16698_ _18192_/CLK _16698_/D vssd1 vssd1 vccd1 vccd1 _16698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18437_ _18437_/CLK _18437_/D vssd1 vssd1 vccd1 vccd1 _18437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15649_ _17194_/CLK _15649_/D vssd1 vssd1 vccd1 vccd1 _15649_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_312_wb_clk_i clkbuf_6_45_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18064_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_115_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09170_ _15553_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09170_/X sky130_fd_sc_hd__or2_1
X_18368_ _18368_/CLK _18368_/D vssd1 vssd1 vccd1 vccd1 _18368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08121_ _13931_/A _08121_/B vssd1 vssd1 vccd1 vccd1 _15699_/D sky130_fd_sc_hd__and2_1
X_17319_ _17319_/CLK hold159/X vssd1 vssd1 vccd1 vccd1 _17319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18299_ _18363_/CLK _18299_/D vssd1 vssd1 vccd1 vccd1 _18299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08052_ _14166_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08052_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3103 _14985_/X vssd1 vssd1 vccd1 vccd1 _18278_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3114 _17815_/Q vssd1 vssd1 vccd1 vccd1 hold3114/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3125 _17401_/Q vssd1 vssd1 vccd1 vccd1 hold3125/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3136 _17450_/Q vssd1 vssd1 vccd1 vccd1 hold3136/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2402 _15580_/Q vssd1 vssd1 vccd1 vccd1 hold2402/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3147 _17473_/Q vssd1 vssd1 vccd1 vccd1 hold3147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2413 _15138_/X vssd1 vssd1 vccd1 vccd1 _18352_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08954_ _08954_/A hold674/X vssd1 vssd1 vccd1 vccd1 _16094_/D sky130_fd_sc_hd__and2_1
Xhold3158 _17396_/Q vssd1 vssd1 vccd1 vccd1 hold3158/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2424 _18289_/Q vssd1 vssd1 vccd1 vccd1 hold2424/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3169 _17999_/Q vssd1 vssd1 vccd1 vccd1 hold3169/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2435 _17937_/Q vssd1 vssd1 vccd1 vccd1 hold2435/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1701 _14687_/X vssd1 vssd1 vccd1 vccd1 _18135_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2446 _08008_/X vssd1 vssd1 vccd1 vccd1 _15645_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07905_ hold2840/X _07924_/B _07904_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _07905_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1712 _18157_/Q vssd1 vssd1 vccd1 vccd1 hold1712/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2457 _18262_/Q vssd1 vssd1 vccd1 vccd1 hold2457/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1723 _15232_/X vssd1 vssd1 vccd1 vccd1 _18398_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08885_ _15274_/A hold881/X vssd1 vssd1 vccd1 vccd1 _16060_/D sky130_fd_sc_hd__and2_1
Xhold2468 _16168_/Q vssd1 vssd1 vccd1 vccd1 hold2468/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1734 _18109_/Q vssd1 vssd1 vccd1 vccd1 hold1734/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2479 _16194_/Q vssd1 vssd1 vccd1 vccd1 hold2479/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1745 _08233_/X vssd1 vssd1 vccd1 vccd1 _15751_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1756 la_data_in[3] vssd1 vssd1 vccd1 vccd1 hold1756/X sky130_fd_sc_hd__dlygate4sd3_1
X_07836_ hold2912/X _07865_/B _07835_/X _14211_/C1 vssd1 vssd1 vccd1 vccd1 _07836_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1767 _14725_/X vssd1 vssd1 vccd1 vccd1 _18154_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1778 _14363_/X vssd1 vssd1 vccd1 vccd1 _14364_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1789 _18336_/Q vssd1 vssd1 vccd1 vccd1 hold1789/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_1384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09506_ hold1913/X _16326_/Q _09992_/C vssd1 vssd1 vccd1 vccd1 _09507_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_78_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09437_ _07804_/A _09483_/A _09440_/B _09436_/X vssd1 vssd1 vccd1 vccd1 _09437_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09368_ _09386_/B _09369_/B _09369_/C _09369_/D vssd1 vssd1 vccd1 vccd1 _09368_/Y
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_19_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08319_ _15543_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08319_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_90_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09299_ _14980_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09299_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_60 hold363/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_71 hold597/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_82 _15145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11330_ hold1628/X _16934_/Q _12305_/C vssd1 vssd1 vccd1 vccd1 _11331_/B sky130_fd_sc_hd__mux2_1
XANTENNA_93 hold5944/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11261_ hold2291/X hold3520/X _11654_/S vssd1 vssd1 vccd1 vccd1 _11262_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5050 _17206_/Q vssd1 vssd1 vccd1 vccd1 hold5050/X sky130_fd_sc_hd__dlygate4sd3_1
X_10212_ _10536_/A _10212_/B vssd1 vssd1 vccd1 vccd1 _10212_/X sky130_fd_sc_hd__or2_1
X_13000_ hold1639/X _17348_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _13000_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5061 _10885_/X vssd1 vssd1 vccd1 vccd1 _16785_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5072 _16795_/Q vssd1 vssd1 vccd1 vccd1 hold5072/X sky130_fd_sc_hd__dlygate4sd3_1
X_11192_ _16888_/Q _11213_/B _11213_/C vssd1 vssd1 vccd1 vccd1 _11192_/X sky130_fd_sc_hd__and3_1
XFILLER_0_203_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5083 _11377_/X vssd1 vssd1 vccd1 vccd1 _16949_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5094 _16326_/Q vssd1 vssd1 vccd1 vccd1 _13078_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4360 _15403_/X vssd1 vssd1 vccd1 vccd1 _15404_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10143_ _10554_/A _10143_/B vssd1 vssd1 vccd1 vccd1 _10143_/X sky130_fd_sc_hd__or2_1
Xhold4371 _12357_/Y vssd1 vssd1 vccd1 vccd1 _12358_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4382 _11190_/Y vssd1 vssd1 vccd1 vccd1 _11191_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4393 _16918_/Q vssd1 vssd1 vccd1 vccd1 hold4393/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3670 _16594_/Q vssd1 vssd1 vccd1 vccd1 hold3670/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3681 _09847_/X vssd1 vssd1 vccd1 vccd1 _16439_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14951_ hold2457/X _14946_/B _14950_/Y _15030_/A vssd1 vssd1 vccd1 vccd1 _14951_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10074_ _13310_/A _10476_/A _10073_/X vssd1 vssd1 vccd1 vccd1 _10074_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3692 _16557_/Q vssd1 vssd1 vccd1 vccd1 hold3692/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13902_ _14457_/A hold2291/X hold297/X vssd1 vssd1 vccd1 vccd1 _13903_/B sky130_fd_sc_hd__mux2_1
XTAP_5887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2980 _08402_/X vssd1 vssd1 vccd1 vccd1 _15831_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17670_ _17734_/CLK _17670_/D vssd1 vssd1 vccd1 vccd1 _17670_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2991 _18123_/Q vssd1 vssd1 vccd1 vccd1 hold2991/X sky130_fd_sc_hd__dlygate4sd3_1
X_14882_ _14952_/A hold332/X vssd1 vssd1 vccd1 vccd1 _14882_/Y sky130_fd_sc_hd__nand2_1
X_16621_ _18087_/CLK _16621_/D vssd1 vssd1 vccd1 vccd1 _16621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13833_ _17571_/Q _13737_/A _13832_/X vssd1 vssd1 vccd1 vccd1 _13833_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_230_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16552_ _18265_/CLK _16552_/D vssd1 vssd1 vccd1 vccd1 _16552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13764_ _13788_/A _13764_/B vssd1 vssd1 vccd1 vccd1 _13764_/X sky130_fd_sc_hd__or2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ hold3023/X hold4167/X _11738_/C vssd1 vssd1 vccd1 vccd1 _10977_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_174_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15503_ hold423/X _18431_/Q _15505_/S vssd1 vssd1 vccd1 vccd1 hold424/A sky130_fd_sc_hd__mux2_1
X_12715_ hold2935/X hold3783/X _12766_/S vssd1 vssd1 vccd1 vccd1 _12715_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16483_ _18396_/CLK _16483_/D vssd1 vssd1 vccd1 vccd1 _16483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13695_ _13791_/A _13695_/B vssd1 vssd1 vccd1 vccd1 _13695_/X sky130_fd_sc_hd__or2_1
XFILLER_0_210_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18222_ _18222_/CLK _18222_/D vssd1 vssd1 vccd1 vccd1 _18222_/Q sky130_fd_sc_hd__dfxtp_1
X_15434_ _15434_/A _15434_/B vssd1 vssd1 vccd1 vccd1 _18419_/D sky130_fd_sc_hd__and2_1
X_12646_ hold1453/X _17393_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12646_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18153_ _18211_/CLK _18153_/D vssd1 vssd1 vccd1 vccd1 _18153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15365_ _15365_/A _15483_/B vssd1 vssd1 vccd1 vccd1 _15365_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12577_ hold2145/X hold3389/X _12985_/S vssd1 vssd1 vccd1 vccd1 _12577_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17104_ _17229_/CLK _17104_/D vssd1 vssd1 vccd1 vccd1 _17104_/Q sky130_fd_sc_hd__dfxtp_1
X_14316_ _15103_/A _14334_/B vssd1 vssd1 vccd1 vccd1 _14316_/X sky130_fd_sc_hd__or2_1
X_18084_ _18188_/CLK _18084_/D vssd1 vssd1 vccd1 vccd1 _18084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11528_ hold2218/X hold4173/X _11717_/C vssd1 vssd1 vccd1 vccd1 _11529_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_80_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15296_ _17333_/Q _09362_/C _15485_/B1 hold569/X vssd1 vssd1 vccd1 vccd1 _15296_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold308 hold308/A vssd1 vssd1 vccd1 vccd1 hold308/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold319 input28/X vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__buf_1
XFILLER_0_150_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17035_ _17883_/CLK _17035_/D vssd1 vssd1 vccd1 vccd1 _17035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14247_ hold2731/X _14268_/B _14246_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _14247_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11459_ hold2418/X _16977_/Q _11654_/S vssd1 vssd1 vccd1 vccd1 _11460_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14178_ _14517_/A _14204_/B vssd1 vssd1 vccd1 vccd1 _14178_/X sky130_fd_sc_hd__or2_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _13129_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13129_/X sky130_fd_sc_hd__and2_1
XFILLER_0_239_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_238_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1008 hold1008/A vssd1 vssd1 vccd1 vccd1 _15531_/A sky130_fd_sc_hd__buf_8
XFILLER_0_225_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17937_ _18028_/CLK _17937_/D vssd1 vssd1 vccd1 vccd1 _17937_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1019 hold6106/X vssd1 vssd1 vccd1 vccd1 hold913/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08670_ _15434_/A hold190/X vssd1 vssd1 vccd1 vccd1 _15956_/D sky130_fd_sc_hd__and2_1
X_17868_ _17868_/CLK _17868_/D vssd1 vssd1 vccd1 vccd1 _17868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16819_ _18321_/CLK _16819_/D vssd1 vssd1 vccd1 vccd1 _16819_/Q sky130_fd_sc_hd__dfxtp_1
X_17799_ _17799_/CLK _17799_/D vssd1 vssd1 vccd1 vccd1 _17799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09222_ hold992/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09222_/X sky130_fd_sc_hd__or2_1
XFILLER_0_185_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09153_ hold2193/X _09164_/B _09152_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _09153_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08104_ _14164_/A hold1726/X hold108/X vssd1 vssd1 vccd1 vccd1 _08104_/X sky130_fd_sc_hd__mux2_1
X_09084_ _15199_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09084_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08035_ _15549_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08035_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold820 hold820/A vssd1 vssd1 vccd1 vccd1 hold820/X sky130_fd_sc_hd__buf_6
XFILLER_0_82_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold831 hold831/A vssd1 vssd1 vccd1 vccd1 hold831/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 hold842/A vssd1 vssd1 vccd1 vccd1 hold842/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold853 hold853/A vssd1 vssd1 vccd1 vccd1 hold853/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_229_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold864 hold864/A vssd1 vssd1 vccd1 vccd1 hold864/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold875 hold875/A vssd1 vssd1 vccd1 vccd1 hold875/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold886 hold886/A vssd1 vssd1 vccd1 vccd1 hold886/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold897 hold897/A vssd1 vssd1 vccd1 vccd1 hold897/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09986_ hold1803/X hold5008/X _09992_/C vssd1 vssd1 vccd1 vccd1 _09987_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_228_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2210 _14005_/X vssd1 vssd1 vccd1 vccd1 _17808_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2221 _15118_/X vssd1 vssd1 vccd1 vccd1 _18343_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2232 _14566_/X vssd1 vssd1 vccd1 vccd1 hold2232/X sky130_fd_sc_hd__dlygate4sd3_1
X_08937_ hold618/X hold716/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold717/A sky130_fd_sc_hd__mux2_1
Xhold2243 _14569_/X vssd1 vssd1 vccd1 vccd1 _18079_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_6_0_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
Xhold2254 _07812_/Y vssd1 vssd1 vccd1 vccd1 hold2254/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1520 _14677_/X vssd1 vssd1 vccd1 vccd1 _18131_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2265 hold2271/X vssd1 vssd1 vccd1 vccd1 _12626_/S sky130_fd_sc_hd__buf_4
Xhold1531 _09415_/X vssd1 vssd1 vccd1 vccd1 _16293_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2276 _07808_/X vssd1 vssd1 vccd1 vccd1 _17752_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2287 _18093_/Q vssd1 vssd1 vccd1 vccd1 hold2287/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1542 input65/X vssd1 vssd1 vccd1 vccd1 hold1542/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08868_ _17520_/Q _08868_/B _13056_/C vssd1 vssd1 vccd1 vccd1 _08868_/X sky130_fd_sc_hd__or3b_4
XFILLER_0_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1553 _09328_/X vssd1 vssd1 vccd1 vccd1 _16274_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2298 _15656_/Q vssd1 vssd1 vccd1 vccd1 hold2298/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1564 _15851_/Q vssd1 vssd1 vccd1 vccd1 hold1564/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1575 _07889_/X vssd1 vssd1 vccd1 vccd1 _15588_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_234_wb_clk_i clkbuf_6_62_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18192_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07819_ _15559_/A _15231_/A vssd1 vssd1 vccd1 vccd1 _09495_/C sky130_fd_sc_hd__nand2_1
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1586 _08314_/X vssd1 vssd1 vccd1 vccd1 _15790_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1597 _14111_/X vssd1 vssd1 vccd1 vccd1 _17859_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08799_ hold618/X hold803/X _08801_/S vssd1 vssd1 vccd1 vccd1 hold804/A sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_212_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10830_ _11103_/A _10830_/B vssd1 vssd1 vccd1 vccd1 _10830_/X sky130_fd_sc_hd__or2_1
XFILLER_0_197_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10761_ _11049_/A _10761_/B vssd1 vssd1 vccd1 vccd1 _10761_/X sky130_fd_sc_hd__or2_1
XFILLER_0_177_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12500_ _17343_/Q _12506_/B vssd1 vssd1 vccd1 vccd1 _12500_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10692_ _11010_/A _10692_/B vssd1 vssd1 vccd1 vccd1 _10692_/X sky130_fd_sc_hd__or2_1
X_13480_ hold3888/X _13795_/A2 _13479_/X _13729_/C1 vssd1 vssd1 vccd1 vccd1 _13480_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12431_ hold438/X hold460/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12432_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15150_ hold6071/X _15165_/B hold1108/X _15212_/C1 vssd1 vssd1 vccd1 vccd1 _15150_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12362_ _17278_/Q _12362_/B _12362_/C vssd1 vssd1 vccd1 vccd1 _12362_/X sky130_fd_sc_hd__and3_1
X_14101_ hold2489/X _14107_/A2 _14100_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _14101_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11313_ _12240_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11313_/X sky130_fd_sc_hd__or2_1
X_15081_ _15189_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15081_/X sky130_fd_sc_hd__or2_1
X_12293_ _17255_/Q _12293_/B _12293_/C vssd1 vssd1 vccd1 vccd1 _12293_/X sky130_fd_sc_hd__and3_1
XFILLER_0_200_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14032_ _15539_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14032_/X sky130_fd_sc_hd__or2_1
X_11244_ _11631_/A _11244_/B vssd1 vssd1 vccd1 vccd1 _11244_/X sky130_fd_sc_hd__or2_1
XFILLER_0_200_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ hold3483/X _11100_/A _11174_/X vssd1 vssd1 vccd1 vccd1 _11175_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4190 _15293_/X vssd1 vssd1 vccd1 vccd1 _15294_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10126_ hold4521/X _10604_/B _10125_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _10126_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15983_ _17345_/CLK _15983_/D vssd1 vssd1 vccd1 vccd1 _15983_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17722_ _17722_/CLK _17722_/D vssd1 vssd1 vccd1 vccd1 _17722_/Q sky130_fd_sc_hd__dfxtp_1
X_14934_ _15203_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14934_/X sky130_fd_sc_hd__or2_1
X_10057_ _10603_/A _10057_/B vssd1 vssd1 vccd1 vccd1 _16509_/D sky130_fd_sc_hd__nor2_1
XTAP_5673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ _17653_/CLK _17653_/D vssd1 vssd1 vccd1 vccd1 _17653_/Q sky130_fd_sc_hd__dfxtp_1
X_14865_ hold2940/X _14880_/B _14864_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14865_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16604_ _18168_/CLK _16604_/D vssd1 vssd1 vccd1 vccd1 _16604_/Q sky130_fd_sc_hd__dfxtp_1
X_13816_ _13819_/A _13816_/B vssd1 vssd1 vccd1 vccd1 _13816_/Y sky130_fd_sc_hd__nor2_1
X_17584_ _17584_/CLK _17584_/D vssd1 vssd1 vccd1 vccd1 _17584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14796_ _15189_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14796_/X sky130_fd_sc_hd__or2_1
XFILLER_0_58_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16535_ _18125_/CLK _16535_/D vssd1 vssd1 vccd1 vccd1 _16535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13747_ hold5553/X _13847_/B _13746_/X _13765_/C1 vssd1 vssd1 vccd1 vccd1 _13747_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10959_ _11631_/A _10959_/B vssd1 vssd1 vccd1 vccd1 _10959_/X sky130_fd_sc_hd__or2_1
XFILLER_0_169_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16466_ _18315_/CLK _16466_/D vssd1 vssd1 vccd1 vccd1 _16466_/Q sky130_fd_sc_hd__dfxtp_1
X_13678_ hold5396/X _13871_/B _13677_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _13678_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18205_ _18205_/CLK _18205_/D vssd1 vssd1 vccd1 vccd1 _18205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15417_ _16094_/Q _09392_/B _15488_/A2 hold515/X vssd1 vssd1 vccd1 vccd1 _15417_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12629_ hold3137/X _12628_/X _12851_/S vssd1 vssd1 vccd1 vccd1 _12629_/X sky130_fd_sc_hd__mux2_1
X_16397_ _18342_/CLK _16397_/D vssd1 vssd1 vccd1 vccd1 _16397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18136_ _18156_/CLK _18136_/D vssd1 vssd1 vccd1 vccd1 _18136_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_38_wb_clk_i clkbuf_6_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17161_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15348_ hold867/X _09386_/A _15441_/A2 hold749/X vssd1 vssd1 vccd1 vccd1 _15348_/X
+ sky130_fd_sc_hd__a22o_1
Xhold5808 _09928_/X vssd1 vssd1 vccd1 vccd1 _16466_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_1372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5819 _17629_/Q vssd1 vssd1 vccd1 vccd1 hold5819/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18067_ _18067_/CLK _18067_/D vssd1 vssd1 vccd1 vccd1 _18067_/Q sky130_fd_sc_hd__dfxtp_1
Xhold105 hold336/X vssd1 vssd1 vccd1 vccd1 hold337/A sky130_fd_sc_hd__clkbuf_8
X_15279_ hold558/X _15485_/A2 _15488_/A2 hold461/X _15278_/X vssd1 vssd1 vccd1 vccd1
+ _15282_/C sky130_fd_sc_hd__a221o_1
Xhold116 hold116/A vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 hold127/A vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold138 hold138/A vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 hold217/X vssd1 vssd1 vccd1 vccd1 hold218/A sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ _17898_/CLK _17018_/D vssd1 vssd1 vccd1 vccd1 _17018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09840_ _09948_/A _09840_/B vssd1 vssd1 vccd1 vccd1 _09840_/X sky130_fd_sc_hd__or2_1
Xfanout607 _09364_/Y vssd1 vssd1 vccd1 vccd1 _15441_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_106_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout618 _09357_/A vssd1 vssd1 vccd1 vccd1 _15487_/A2 sky130_fd_sc_hd__buf_6
Xfanout629 hold354/X vssd1 vssd1 vccd1 vccd1 hold355/A sky130_fd_sc_hd__buf_1
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09771_ _09957_/A _09771_/B vssd1 vssd1 vccd1 vccd1 _09771_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _12416_/A hold530/X vssd1 vssd1 vccd1 vccd1 _15982_/D sky130_fd_sc_hd__and2_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_234_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08653_ hold82/X hold455/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold456/A sky130_fd_sc_hd__mux2_1
XFILLER_0_233_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08584_ hold315/X hold763/X _08592_/S vssd1 vssd1 vccd1 vccd1 _08585_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09205_ hold2673/X _09214_/B _09204_/X _12753_/A vssd1 vssd1 vccd1 vccd1 _09205_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09136_ _15519_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09136_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09067_ _15182_/A hold363/X vssd1 vssd1 vccd1 vccd1 _09098_/B sky130_fd_sc_hd__or2_2
XFILLER_0_5_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08018_ hold1303/X _08029_/B _08017_/X _12103_/C1 vssd1 vssd1 vccd1 vccd1 _08018_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold650 hold650/A vssd1 vssd1 vccd1 vccd1 hold650/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold661 hold661/A vssd1 vssd1 vccd1 vccd1 hold661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 input36/X vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 input30/X vssd1 vssd1 vccd1 vccd1 hold683/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 hold694/A vssd1 vssd1 vccd1 vccd1 hold694/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09969_ _09978_/A _09969_/B vssd1 vssd1 vccd1 vccd1 _09969_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_415_wb_clk_i clkbuf_6_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17910_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2040 _13949_/X vssd1 vssd1 vccd1 vccd1 _17781_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2051 _18213_/Q vssd1 vssd1 vccd1 vccd1 hold2051/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2062 _17820_/Q vssd1 vssd1 vccd1 vccd1 hold2062/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2073 _18128_/Q vssd1 vssd1 vccd1 vccd1 hold2073/X sky130_fd_sc_hd__dlygate4sd3_1
X_12980_ hold3624/X _12979_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12980_/X sky130_fd_sc_hd__mux2_1
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2084 _14398_/X vssd1 vssd1 vccd1 vccd1 _17997_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2095 _14261_/X vssd1 vssd1 vccd1 vccd1 _17931_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1350 _18442_/Q vssd1 vssd1 vccd1 vccd1 hold1350/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1361 _14271_/X vssd1 vssd1 vccd1 vccd1 _17936_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1372 _15840_/Q vssd1 vssd1 vccd1 vccd1 hold1372/X sky130_fd_sc_hd__dlygate4sd3_1
X_11931_ _13482_/A _11931_/B vssd1 vssd1 vccd1 vccd1 _11931_/X sky130_fd_sc_hd__or2_1
XFILLER_0_197_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1383 _07963_/X vssd1 vssd1 vccd1 vccd1 _15624_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1394 _14105_/X vssd1 vssd1 vccd1 vccd1 _17857_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14650_ _15205_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14650_/X sky130_fd_sc_hd__or2_1
XFILLER_0_135_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _12273_/A _11862_/B vssd1 vssd1 vccd1 vccd1 _11862_/X sky130_fd_sc_hd__or2_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13601_ hold1203/X _17654_/Q _13766_/S vssd1 vssd1 vccd1 vccd1 _13602_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_95_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10813_ hold5335/X _11195_/B _10812_/X _14462_/C1 vssd1 vssd1 vccd1 vccd1 _10813_/X
+ sky130_fd_sc_hd__o211a_1
X_14581_ hold3163/X _14612_/B _14580_/X _14697_/C1 vssd1 vssd1 vccd1 vccd1 _14581_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ hold4427/X _11697_/A _11792_/X vssd1 vssd1 vccd1 vccd1 _11793_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16320_ _16323_/CLK _16320_/D vssd1 vssd1 vccd1 vccd1 _16320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13532_ hold1081/X _17631_/Q _13829_/C vssd1 vssd1 vccd1 vccd1 _13533_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_138_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10744_ hold4117/X _11789_/B _10743_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _10744_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16251_ _17430_/CLK _16251_/D vssd1 vssd1 vccd1 vccd1 hold980/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13463_ hold2285/X hold4077/X _13463_/S vssd1 vssd1 vccd1 vccd1 _13464_/B sky130_fd_sc_hd__mux2_1
X_10675_ hold4666/X _11153_/B _10674_/X _14552_/C1 vssd1 vssd1 vccd1 vccd1 _10675_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15202_ hold3087/X _15221_/B _15201_/X _15202_/C1 vssd1 vssd1 vccd1 vccd1 _15202_/X
+ sky130_fd_sc_hd__o211a_1
X_12414_ _15274_/A hold801/X vssd1 vssd1 vccd1 vccd1 _17300_/D sky130_fd_sc_hd__and2_1
XFILLER_0_207_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16182_ _17468_/CLK _16182_/D vssd1 vssd1 vccd1 vccd1 _16182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13394_ hold1340/X hold4424/X _13874_/C vssd1 vssd1 vccd1 vccd1 _13395_/B sky130_fd_sc_hd__mux2_1
X_15133_ _15187_/A _15157_/B vssd1 vssd1 vccd1 vccd1 _15133_/X sky130_fd_sc_hd__or2_1
X_12345_ hold3453/X _12273_/A _12344_/X vssd1 vssd1 vccd1 vccd1 _12345_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15064_ _15064_/A _15064_/B vssd1 vssd1 vccd1 vccd1 _18317_/D sky130_fd_sc_hd__and2_1
X_12276_ _13749_/A _12276_/B vssd1 vssd1 vccd1 vccd1 _12276_/X sky130_fd_sc_hd__or2_1
XFILLER_0_142_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14015_ hold2873/X _14038_/B _14014_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _14015_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_1278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11227_ _12337_/A _11227_/B vssd1 vssd1 vccd1 vccd1 _11227_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_235_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_156_wb_clk_i clkbuf_6_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17321_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11158_ _11158_/A _11158_/B vssd1 vssd1 vccd1 vccd1 _16876_/D sky130_fd_sc_hd__nor2_1
XTAP_6171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10109_ hold2491/X _16527_/Q _10625_/C vssd1 vssd1 vccd1 vccd1 _10110_/B sky130_fd_sc_hd__mux2_1
X_15966_ _17328_/CLK _15966_/D vssd1 vssd1 vccd1 vccd1 hold689/A sky130_fd_sc_hd__dfxtp_1
X_11089_ hold3942/X _11225_/B _11088_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _11089_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14917_ hold1881/X _14952_/B _14916_/X _15042_/A vssd1 vssd1 vccd1 vccd1 _14917_/X
+ sky130_fd_sc_hd__o211a_1
X_17705_ _17705_/CLK _17705_/D vssd1 vssd1 vccd1 vccd1 _17705_/Q sky130_fd_sc_hd__dfxtp_1
X_15897_ _17345_/CLK _15897_/D vssd1 vssd1 vccd1 vccd1 _15897_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_31_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_31_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14848_ _15187_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14848_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17636_ _17732_/CLK _17636_/D vssd1 vssd1 vccd1 vccd1 _17636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17567_ _17599_/CLK _17567_/D vssd1 vssd1 vccd1 vccd1 _17567_/Q sky130_fd_sc_hd__dfxtp_1
X_14779_ hold2161/X _14774_/B _14778_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14779_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16518_ _18214_/CLK _16518_/D vssd1 vssd1 vccd1 vccd1 _16518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17498_ _17499_/CLK _17498_/D vssd1 vssd1 vccd1 vccd1 _17498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16449_ _18394_/CLK _16449_/D vssd1 vssd1 vccd1 vccd1 _16449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18119_ _18149_/CLK _18119_/D vssd1 vssd1 vccd1 vccd1 _18119_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5605 _17717_/Q vssd1 vssd1 vccd1 vccd1 hold5605/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5616 _16658_/Q vssd1 vssd1 vccd1 vccd1 hold5616/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5627 _11056_/X vssd1 vssd1 vccd1 vccd1 _16842_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5638 _11425_/X vssd1 vssd1 vccd1 vccd1 _16965_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4904 _12004_/X vssd1 vssd1 vccd1 vccd1 _17158_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5649 _16968_/Q vssd1 vssd1 vccd1 vccd1 hold5649/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4915 _17208_/Q vssd1 vssd1 vccd1 vccd1 hold4915/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4926 _10990_/X vssd1 vssd1 vccd1 vccd1 _16820_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4937 _17255_/Q vssd1 vssd1 vccd1 vccd1 hold4937/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4948 _11476_/X vssd1 vssd1 vccd1 vccd1 _16982_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4959 _16824_/Q vssd1 vssd1 vccd1 vccd1 hold4959/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout404 _14340_/X vssd1 vssd1 vccd1 vccd1 _14381_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout415 _14140_/B vssd1 vssd1 vccd1 vccd1 _14160_/B sky130_fd_sc_hd__buf_8
XFILLER_0_201_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout426 _13946_/Y vssd1 vssd1 vccd1 vccd1 _13986_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_238_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09823_ hold4622/X _10013_/B _09822_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _09823_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout437 _13721_/S vssd1 vssd1 vccd1 vccd1 _13811_/C sky130_fd_sc_hd__buf_6
XFILLER_0_201_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout448 _11717_/C vssd1 vssd1 vccd1 vccd1 _12305_/C sky130_fd_sc_hd__buf_6
Xfanout459 _13868_/C vssd1 vssd1 vccd1 vccd1 _13871_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_226_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_214_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09754_ hold3755/X _11204_/B _09753_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _09754_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08705_ hold5/X hold471/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08706_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09685_ hold3864/X _10571_/B _09684_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _09685_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _15344_/A _08636_/B vssd1 vssd1 vccd1 vccd1 _15940_/D sky130_fd_sc_hd__and2_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08567_ _15364_/A _08567_/B vssd1 vssd1 vccd1 vccd1 _15907_/D sky130_fd_sc_hd__and2_1
XFILLER_0_232_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08498_ _14443_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08498_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ hold2376/X hold3882/X _11186_/C vssd1 vssd1 vccd1 vccd1 _10461_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_190_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09119_ hold1639/X _09106_/B _09118_/X _15244_/A vssd1 vssd1 vccd1 vccd1 _09119_/X
+ sky130_fd_sc_hd__o211a_1
X_10391_ hold1781/X _16621_/Q _10595_/C vssd1 vssd1 vccd1 vccd1 _10392_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_165_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12130_ hold4893/X _12353_/B _12129_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _12130_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12061_ hold5745/X _12362_/B _12060_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _12061_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold480 hold480/A vssd1 vssd1 vccd1 vccd1 hold480/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold491 hold491/A vssd1 vssd1 vccd1 vccd1 hold491/X sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ hold2962/X hold4955/X _11204_/C vssd1 vssd1 vccd1 vccd1 _11013_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_216_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15820_ _17731_/CLK hold222/X vssd1 vssd1 vccd1 vccd1 _15820_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15751_ _17702_/CLK _15751_/D vssd1 vssd1 vccd1 vccd1 _15751_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12963_ _14358_/A _12963_/B vssd1 vssd1 vccd1 vccd1 _17497_/D sky130_fd_sc_hd__and2_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1180 hold6109/X vssd1 vssd1 vccd1 vccd1 hold690/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _14988_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14702_/X sky130_fd_sc_hd__or2_1
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1191 hold925/X vssd1 vssd1 vccd1 vccd1 input37/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11914_ hold4654/X _13811_/B _11913_/X _08363_/A vssd1 vssd1 vccd1 vccd1 _11914_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15682_ _17906_/CLK _15682_/D vssd1 vssd1 vccd1 vccd1 _15682_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12894_ _12894_/A _12894_/B vssd1 vssd1 vccd1 vccd1 _17474_/D sky130_fd_sc_hd__and2_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _17661_/CLK _17421_/D vssd1 vssd1 vccd1 vccd1 _17421_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14633_ hold1734/X _14664_/B _14632_/X _14769_/C1 vssd1 vssd1 vccd1 vccd1 _14633_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11845_ hold5509/X _12329_/B _11844_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11845_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _17516_/CLK _17352_/D vssd1 vssd1 vccd1 vccd1 _17352_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _15492_/A _14573_/B hold2279/X vssd1 vssd1 vccd1 vccd1 _14564_/X sky130_fd_sc_hd__a21o_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _12337_/A _11776_/B vssd1 vssd1 vccd1 vccd1 _11776_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_83_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16303_ _17291_/CLK hold715/X vssd1 vssd1 vccd1 vccd1 _16303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13515_ _13719_/A _13515_/B vssd1 vssd1 vccd1 vccd1 _13515_/X sky130_fd_sc_hd__or2_1
X_17283_ _17735_/CLK _17283_/D vssd1 vssd1 vccd1 vccd1 _17283_/Q sky130_fd_sc_hd__dfxtp_1
X_10727_ hold1360/X hold4399/X _11660_/S vssd1 vssd1 vccd1 vccd1 _10728_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_126_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14495_ hold820/X _14499_/B vssd1 vssd1 vccd1 vccd1 _14495_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16234_ _17754_/CLK _16234_/D vssd1 vssd1 vccd1 vccd1 _16234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13446_ _13734_/A _13446_/B vssd1 vssd1 vccd1 vccd1 _13446_/X sky130_fd_sc_hd__or2_1
X_10658_ hold2149/X hold4079/X _11732_/C vssd1 vssd1 vccd1 vccd1 _10659_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16165_ _17513_/CLK _16165_/D vssd1 vssd1 vccd1 vccd1 _16165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13377_ _13752_/A _13377_/B vssd1 vssd1 vccd1 vccd1 _13377_/X sky130_fd_sc_hd__or2_1
X_10589_ _10589_/A _10589_/B _10640_/C vssd1 vssd1 vccd1 vccd1 _10589_/X sky130_fd_sc_hd__and3_1
XFILLER_0_152_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15116_ hold1624/X hold341/X _15115_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _15116_/X
+ sky130_fd_sc_hd__o211a_1
X_12328_ _13873_/A _12328_/B vssd1 vssd1 vccd1 vccd1 _12328_/Y sky130_fd_sc_hd__nor2_1
X_16096_ _18419_/CLK _16096_/D vssd1 vssd1 vccd1 vccd1 _16096_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_337_wb_clk_i clkbuf_6_43_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17281_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_220_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15047_ _09313_/A hold1262/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15048_/B sky130_fd_sc_hd__mux2_1
X_12259_ hold4843/X _12353_/B _12258_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _12259_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2809 _16224_/Q vssd1 vssd1 vccd1 vccd1 hold2809/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16998_ _17846_/CLK _16998_/D vssd1 vssd1 vccd1 vccd1 _16998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15949_ _18425_/CLK _15949_/D vssd1 vssd1 vccd1 vccd1 hold455/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09470_ _09471_/B _09478_/B _09470_/C vssd1 vssd1 vccd1 vccd1 _16317_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_176_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08421_ _14529_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08421_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17619_ _17620_/CLK _17619_/D vssd1 vssd1 vccd1 vccd1 _17619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_wb_clk_i clkbuf_6_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17985_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08352_ _15521_/A hold2615/X hold115/X vssd1 vssd1 vccd1 vccd1 _08353_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_157_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08283_ _08504_/A hold338/X vssd1 vssd1 vccd1 vccd1 _08283_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_46_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6103 _17523_/Q vssd1 vssd1 vccd1 vccd1 hold6103/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6114 data_in[14] vssd1 vssd1 vccd1 vccd1 hold604/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6125 _16313_/Q vssd1 vssd1 vccd1 vccd1 hold6125/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5402 _17742_/Q vssd1 vssd1 vccd1 vccd1 hold5402/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5413 _13690_/X vssd1 vssd1 vccd1 vccd1 _17683_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5424 _16696_/Q vssd1 vssd1 vccd1 vccd1 hold5424/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5435 _11248_/X vssd1 vssd1 vccd1 vccd1 _16906_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4701 _16867_/Q vssd1 vssd1 vccd1 vccd1 hold4701/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5446 _16746_/Q vssd1 vssd1 vccd1 vccd1 hold5446/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4712 _09841_/X vssd1 vssd1 vccd1 vccd1 _16437_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5457 _12124_/X vssd1 vssd1 vccd1 vccd1 _17198_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5468 _17237_/Q vssd1 vssd1 vccd1 vccd1 hold5468/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4723 _12330_/Y vssd1 vssd1 vccd1 vccd1 _12331_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4734 _13732_/X vssd1 vssd1 vccd1 vccd1 _17697_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5479 _13750_/X vssd1 vssd1 vccd1 vccd1 _17703_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4745 _17094_/Q vssd1 vssd1 vccd1 vccd1 hold4745/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4756 _17692_/Q vssd1 vssd1 vccd1 vccd1 hold4756/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4767 _11131_/X vssd1 vssd1 vccd1 vccd1 _16867_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout201 _11210_/B vssd1 vssd1 vccd1 vccd1 _11753_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4778 _09520_/X vssd1 vssd1 vccd1 vccd1 _16330_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout212 _10013_/B vssd1 vssd1 vccd1 vccd1 _11144_/B sky130_fd_sc_hd__buf_4
XFILLER_0_26_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout223 _10070_/B vssd1 vssd1 vccd1 vccd1 _11204_/B sky130_fd_sc_hd__buf_4
Xhold4789 _16994_/Q vssd1 vssd1 vccd1 vccd1 hold4789/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout234 _10067_/B vssd1 vssd1 vccd1 vccd1 _10046_/B sky130_fd_sc_hd__buf_4
XFILLER_0_201_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout245 _10637_/B vssd1 vssd1 vccd1 vccd1 _10631_/B sky130_fd_sc_hd__buf_4
XFILLER_0_5_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout256 _12216_/A vssd1 vssd1 vccd1 vccd1 _13794_/A sky130_fd_sc_hd__buf_4
X_09806_ hold2631/X _16426_/Q _11162_/C vssd1 vssd1 vccd1 vccd1 _09807_/B sky130_fd_sc_hd__mux2_1
Xfanout267 _11553_/A vssd1 vssd1 vccd1 vccd1 _12219_/A sky130_fd_sc_hd__buf_4
Xfanout278 fanout299/X vssd1 vssd1 vccd1 vccd1 _12159_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_214_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout289 _11100_/A vssd1 vssd1 vccd1 vccd1 _11658_/A sky130_fd_sc_hd__buf_4
X_07998_ hold1837/X _08033_/B _07997_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _07998_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_213_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09737_ hold1179/X hold3602/X _10031_/C vssd1 vssd1 vccd1 vccd1 _09738_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09668_ hold3051/X _16380_/Q _10040_/C vssd1 vssd1 vccd1 vccd1 _09669_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ hold23/X hold302/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08620_/B sky130_fd_sc_hd__mux2_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09599_ hold1958/X _16357_/Q _10025_/C vssd1 vssd1 vccd1 vccd1 _09600_/B sky130_fd_sc_hd__mux2_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11630_ hold884/X hold5440/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11631_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11561_ hold1596/X _17011_/Q _11753_/C vssd1 vssd1 vccd1 vccd1 _11562_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_181_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13300_ hold4414/X _13299_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13300_/X sky130_fd_sc_hd__mux2_1
X_10512_ _10536_/A _10512_/B vssd1 vssd1 vccd1 vccd1 _10512_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14280_ _15229_/A _14282_/B vssd1 vssd1 vccd1 vccd1 _14280_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11492_ hold2884/X hold4101/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11493_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_61_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13231_ _13311_/A1 _13229_/X _13230_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13231_/X
+ sky130_fd_sc_hd__o211a_1
X_10443_ _10563_/A _10443_/B vssd1 vssd1 vccd1 vccd1 _10443_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13162_ _17571_/Q _17105_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13162_/X sky130_fd_sc_hd__mux2_1
X_10374_ _10530_/A _10374_/B vssd1 vssd1 vccd1 vccd1 _10374_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_430_wb_clk_i clkbuf_6_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17599_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_62_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12113_ hold2618/X hold5543/X _12299_/C vssd1 vssd1 vccd1 vccd1 _12114_/B sky130_fd_sc_hd__mux2_1
Xhold5980 _16321_/Q vssd1 vssd1 vccd1 vccd1 _09483_/B sky130_fd_sc_hd__dlygate4sd3_1
X_13093_ _13092_/X hold3428/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13093_/X sky130_fd_sc_hd__mux2_1
X_17970_ _18194_/CLK _17970_/D vssd1 vssd1 vccd1 vccd1 _17970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5991 _16908_/Q vssd1 vssd1 vccd1 vccd1 hold5991/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12044_ hold1173/X _17172_/Q _13463_/S vssd1 vssd1 vccd1 vccd1 _12045_/B sky130_fd_sc_hd__mux2_1
X_16921_ _17865_/CLK _16921_/D vssd1 vssd1 vccd1 vccd1 _16921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16852_ _18063_/CLK _16852_/D vssd1 vssd1 vccd1 vccd1 _16852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout790 fanout791/X vssd1 vssd1 vccd1 vccd1 _14350_/A sky130_fd_sc_hd__buf_2
X_15803_ _17639_/CLK _15803_/D vssd1 vssd1 vccd1 vccd1 _15803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16783_ _18050_/CLK _16783_/D vssd1 vssd1 vccd1 vccd1 _16783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13995_ hold1457/X _13995_/A2 _13994_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _13995_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15734_ _17705_/CLK _15734_/D vssd1 vssd1 vccd1 vccd1 _15734_/Q sky130_fd_sc_hd__dfxtp_1
X_12946_ hold1260/X hold4015/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12946_/X sky130_fd_sc_hd__mux2_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15665_ _17157_/CLK _15665_/D vssd1 vssd1 vccd1 vccd1 _15665_/Q sky130_fd_sc_hd__dfxtp_1
X_18453_ _18453_/CLK _18453_/D vssd1 vssd1 vccd1 vccd1 _18453_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ hold3010/X hold3152/X _12916_/S vssd1 vssd1 vccd1 vccd1 _12877_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14616_ _15225_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14616_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17404_ _18457_/CLK _17404_/D vssd1 vssd1 vccd1 vccd1 _17404_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18384_ _18384_/CLK _18384_/D vssd1 vssd1 vccd1 vccd1 _18384_/Q sky130_fd_sc_hd__dfxtp_1
X_11828_ hold1305/X hold3470/X _13796_/S vssd1 vssd1 vccd1 vccd1 _11829_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_56_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15596_ _17244_/CLK _15596_/D vssd1 vssd1 vccd1 vccd1 _15596_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _17335_/CLK hold33/X vssd1 vssd1 vccd1 vccd1 _17335_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14547_ _14726_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14547_/X sky130_fd_sc_hd__or2_1
X_11759_ _17077_/Q _11765_/B _11765_/C vssd1 vssd1 vccd1 vccd1 _11759_/X sky130_fd_sc_hd__and3_1
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17266_ _17266_/CLK _17266_/D vssd1 vssd1 vccd1 vccd1 _17266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14478_ hold1407/X _14481_/B _14477_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _14478_/X
+ sky130_fd_sc_hd__o211a_1
X_16217_ _17724_/CLK _16217_/D vssd1 vssd1 vccd1 vccd1 _16217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13429_ hold4813/X _13811_/B _13428_/X _08363_/A vssd1 vssd1 vccd1 vccd1 _13429_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17197_ _17261_/CLK _17197_/D vssd1 vssd1 vccd1 vccd1 _17197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16148_ _17345_/CLK _16148_/D vssd1 vssd1 vccd1 vccd1 hold387/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4008 _10489_/X vssd1 vssd1 vccd1 vccd1 _16653_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_171_wb_clk_i clkbuf_6_48_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18030_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4019 _11266_/X vssd1 vssd1 vccd1 vccd1 _16912_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08970_ _15364_/A hold255/X vssd1 vssd1 vccd1 vccd1 _16102_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_100_wb_clk_i clkbuf_6_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16058_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16079_ _17291_/CLK _16079_/D vssd1 vssd1 vccd1 vccd1 hold782/A sky130_fd_sc_hd__dfxtp_1
Xhold3307 _12875_/X vssd1 vssd1 vccd1 vccd1 _12876_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3318 _17462_/Q vssd1 vssd1 vccd1 vccd1 hold3318/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3329 _10135_/X vssd1 vssd1 vccd1 vccd1 _16535_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2606 _15114_/X vssd1 vssd1 vccd1 vccd1 _18341_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07921_ hold2599/X _07924_/B _07920_/Y _15494_/A vssd1 vssd1 vccd1 vccd1 _07921_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2617 _07856_/X vssd1 vssd1 vccd1 vccd1 _15573_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2628 _13957_/X vssd1 vssd1 vccd1 vccd1 _17785_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2639 _17803_/Q vssd1 vssd1 vccd1 vccd1 hold2639/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1905 _18107_/Q vssd1 vssd1 vccd1 vccd1 hold1905/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1916 _14275_/X vssd1 vssd1 vccd1 vccd1 _17938_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07852_ hold2539/X _07869_/B _07851_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _07852_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1927 _17996_/Q vssd1 vssd1 vccd1 vccd1 hold1927/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1938 _15556_/X vssd1 vssd1 vccd1 vccd1 _18456_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1949 _18389_/Q vssd1 vssd1 vccd1 vccd1 hold1949/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput1 input1/A vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
X_07783_ hold384/X vssd1 vssd1 vccd1 vccd1 _07783_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_155_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09522_ _09912_/A _09522_/B vssd1 vssd1 vccd1 vccd1 _09522_/X sky130_fd_sc_hd__or2_1
XFILLER_0_211_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_231_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09453_ _09456_/B _09456_/C _09456_/D vssd1 vssd1 vccd1 vccd1 _09455_/B sky130_fd_sc_hd__and3_1
XFILLER_0_188_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08404_ hold2388/X _08442_/A2 _08403_/X _08361_/A vssd1 vssd1 vccd1 vccd1 _08404_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09384_ hold475/X _15474_/B _09383_/X _07809_/B vssd1 vssd1 vccd1 vccd1 _09384_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08335_ _14732_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08335_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08266_ _15545_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08266_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_166_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_259_wb_clk_i clkbuf_6_58_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17971_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08197_ _15531_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08197_/X sky130_fd_sc_hd__or2_1
XFILLER_0_166_1395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5210 _11005_/X vssd1 vssd1 vccd1 vccd1 _16825_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5221 _17019_/Q vssd1 vssd1 vccd1 vccd1 hold5221/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5232 _13456_/X vssd1 vssd1 vccd1 vccd1 _17605_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5243 _16750_/Q vssd1 vssd1 vccd1 vccd1 hold5243/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5254 _11557_/X vssd1 vssd1 vccd1 vccd1 _17009_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4520 _12533_/X vssd1 vssd1 vccd1 vccd1 _12534_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5265 _17732_/Q vssd1 vssd1 vccd1 vccd1 hold5265/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4531 _16728_/Q vssd1 vssd1 vccd1 vccd1 hold4531/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5276 _12283_/X vssd1 vssd1 vccd1 vccd1 _17251_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5287 _17739_/Q vssd1 vssd1 vccd1 vccd1 hold5287/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4542 _13543_/X vssd1 vssd1 vccd1 vccd1 _17634_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4553 _12551_/X vssd1 vssd1 vccd1 vccd1 _12552_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5298 _11134_/X vssd1 vssd1 vccd1 vccd1 _16868_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4564 _12142_/X vssd1 vssd1 vccd1 vccd1 _17204_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3830 _16669_/Q vssd1 vssd1 vccd1 vccd1 hold3830/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4575 _16753_/Q vssd1 vssd1 vccd1 vccd1 hold4575/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3841 _10123_/X vssd1 vssd1 vccd1 vccd1 _16531_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10090_ hold3616/X _10568_/B _10089_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _16520_/D
+ sky130_fd_sc_hd__o211a_1
Xhold4586 _11977_/X vssd1 vssd1 vccd1 vccd1 _17149_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3852 _16695_/Q vssd1 vssd1 vccd1 vccd1 hold3852/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4597 _11902_/X vssd1 vssd1 vccd1 vccd1 _17124_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3863 _10483_/X vssd1 vssd1 vccd1 vccd1 _16651_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3874 _16549_/Q vssd1 vssd1 vccd1 vccd1 hold3874/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3885 _10198_/X vssd1 vssd1 vccd1 vccd1 _16556_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3896 _10459_/X vssd1 vssd1 vccd1 vccd1 _16643_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_215_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12800_ hold3350/X _12799_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12800_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13780_ hold5416/X _13883_/B _13779_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _13780_/X
+ sky130_fd_sc_hd__o211a_1
X_10992_ _11121_/A _10992_/B vssd1 vssd1 vccd1 vccd1 _10992_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ hold3165/X _12730_/X _12749_/S vssd1 vssd1 vccd1 vccd1 _12731_/X sky130_fd_sc_hd__mux2_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ hold757/X _15485_/A2 _15485_/B1 hold876/X _15448_/X vssd1 vssd1 vccd1 vccd1
+ _15452_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_84_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ hold3133/X _12661_/X _12851_/S vssd1 vssd1 vccd1 vccd1 _12662_/X sky130_fd_sc_hd__mux2_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14401_ _15189_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14401_/X sky130_fd_sc_hd__or2_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _12285_/A _11613_/B vssd1 vssd1 vccd1 vccd1 _11613_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15381_ _16302_/Q _09362_/A _09392_/B hold796/X _15380_/X vssd1 vssd1 vccd1 vccd1
+ _15382_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_0_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12593_ hold3118/X _12592_/X _12905_/S vssd1 vssd1 vccd1 vccd1 _12593_/X sky130_fd_sc_hd__mux2_1
X_17120_ _17271_/CLK _17120_/D vssd1 vssd1 vccd1 vccd1 _17120_/Q sky130_fd_sc_hd__dfxtp_1
X_14332_ _15173_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14332_/X sky130_fd_sc_hd__or2_1
XFILLER_0_167_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11544_ _11649_/A _11544_/B vssd1 vssd1 vccd1 vccd1 _11544_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17051_ _17771_/CLK _17051_/D vssd1 vssd1 vccd1 vccd1 _17051_/Q sky130_fd_sc_hd__dfxtp_1
X_14263_ hold2004/X _14272_/B _14262_/X _14526_/C1 vssd1 vssd1 vccd1 vccd1 _14263_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11475_ _11661_/A _11475_/B vssd1 vssd1 vccd1 vccd1 _11475_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16002_ _18409_/CLK _16002_/D vssd1 vssd1 vccd1 vccd1 hold563/A sky130_fd_sc_hd__dfxtp_1
X_13214_ _13214_/A _13294_/B vssd1 vssd1 vccd1 vccd1 _13214_/X sky130_fd_sc_hd__or2_1
X_10426_ hold5420/X _11213_/B _10425_/X _14342_/A vssd1 vssd1 vccd1 vccd1 _10426_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14194_ _14194_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14194_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13145_ _13145_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13145_/X sky130_fd_sc_hd__and2_1
X_10357_ hold4620/X _10646_/B _10356_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10357_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ _18030_/CLK _17953_/D vssd1 vssd1 vccd1 vccd1 _17953_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ hold4079/X _13075_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13076_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_237_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10288_ hold5048/X _10070_/B _10287_/X _15160_/C1 vssd1 vssd1 vccd1 vccd1 _10288_/X
+ sky130_fd_sc_hd__o211a_1
X_12027_ _13482_/A _12027_/B vssd1 vssd1 vccd1 vccd1 _12027_/X sky130_fd_sc_hd__or2_1
X_16904_ _17161_/CLK _16904_/D vssd1 vssd1 vccd1 vccd1 _16904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17884_ _17884_/CLK hold581/X vssd1 vssd1 vccd1 vccd1 _17884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_217_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16835_ _18070_/CLK _16835_/D vssd1 vssd1 vccd1 vccd1 _16835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16766_ _18028_/CLK _16766_/D vssd1 vssd1 vccd1 vccd1 _16766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13978_ _14604_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13978_/X sky130_fd_sc_hd__or2_1
XFILLER_0_215_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12929_ hold4445/X _12928_/X _12929_/S vssd1 vssd1 vccd1 vccd1 _12929_/X sky130_fd_sc_hd__mux2_1
X_15717_ _17093_/CLK _15717_/D vssd1 vssd1 vccd1 vccd1 _15717_/Q sky130_fd_sc_hd__dfxtp_1
X_16697_ _18223_/CLK _16697_/D vssd1 vssd1 vccd1 vccd1 _16697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18436_ _18438_/CLK _18436_/D vssd1 vssd1 vccd1 vccd1 _18436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15648_ _17628_/CLK _15648_/D vssd1 vssd1 vccd1 vccd1 _15648_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18367_ _18399_/CLK _18367_/D vssd1 vssd1 vccd1 vccd1 _18367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15579_ _17144_/CLK _15579_/D vssd1 vssd1 vccd1 vccd1 _15579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08120_ _15525_/A hold3124/X hold108/X vssd1 vssd1 vccd1 vccd1 _08121_/B sky130_fd_sc_hd__mux2_1
X_17318_ _17318_/CLK hold39/X vssd1 vssd1 vccd1 vccd1 _17318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_352_wb_clk_i clkbuf_6_40_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17748_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18298_ _18298_/CLK _18298_/D vssd1 vssd1 vccd1 vccd1 _18298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08051_ hold2077/X _08097_/A2 _08050_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _08051_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_189_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17249_ _17279_/CLK _17249_/D vssd1 vssd1 vccd1 vccd1 _17249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3104 _17926_/Q vssd1 vssd1 vccd1 vccd1 hold3104/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3115 _14019_/X vssd1 vssd1 vccd1 vccd1 _17815_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3126 _12674_/X vssd1 vssd1 vccd1 vccd1 _12675_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08953_ hold673/X _16094_/Q _08997_/S vssd1 vssd1 vccd1 vccd1 hold674/A sky130_fd_sc_hd__mux2_1
Xhold3137 _17386_/Q vssd1 vssd1 vccd1 vccd1 hold3137/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2403 _07870_/X vssd1 vssd1 vccd1 vccd1 _15580_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3148 _12890_/X vssd1 vssd1 vccd1 vccd1 _12891_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2414 _15647_/Q vssd1 vssd1 vccd1 vccd1 hold2414/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3159 _17474_/Q vssd1 vssd1 vccd1 vccd1 hold3159/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2425 _15007_/X vssd1 vssd1 vccd1 vccd1 _18289_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07904_ _14413_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07904_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2436 _14273_/X vssd1 vssd1 vccd1 vccd1 _17937_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1702 _16163_/Q vssd1 vssd1 vccd1 vccd1 hold1702/X sky130_fd_sc_hd__dlygate4sd3_1
X_08884_ hold679/X hold880/X _08930_/S vssd1 vssd1 vccd1 vccd1 hold881/A sky130_fd_sc_hd__mux2_1
Xhold2447 _16167_/Q vssd1 vssd1 vccd1 vccd1 hold2447/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1713 _14731_/X vssd1 vssd1 vccd1 vccd1 _18157_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2458 _14951_/X vssd1 vssd1 vccd1 vccd1 _18262_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1724 _18105_/Q vssd1 vssd1 vccd1 vccd1 hold1724/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2469 _09107_/X vssd1 vssd1 vccd1 vccd1 _16168_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1735 _14633_/X vssd1 vssd1 vccd1 vccd1 _18109_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1746 _17916_/Q vssd1 vssd1 vccd1 vccd1 hold1746/X sky130_fd_sc_hd__dlygate4sd3_1
X_07835_ _15513_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07835_/X sky130_fd_sc_hd__or2_1
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1757 hold1757/A vssd1 vssd1 vccd1 vccd1 input62/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1768 _16309_/Q vssd1 vssd1 vccd1 vccd1 _09447_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1779 _18240_/Q vssd1 vssd1 vccd1 vccd1 hold1779/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09505_ hold3716/X _10004_/B _09504_/X _08954_/A vssd1 vssd1 vccd1 vccd1 _09505_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09436_ _09438_/B _16304_/Q vssd1 vssd1 vccd1 vccd1 _09436_/X sky130_fd_sc_hd__or2_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _09367_/A _09386_/D vssd1 vssd1 vccd1 vccd1 _09369_/D sky130_fd_sc_hd__or2_1
XFILLER_0_35_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08318_ hold2669/X _08323_/B _08317_/Y _08361_/A vssd1 vssd1 vccd1 vccd1 _08318_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09298_ hold1121/X _09325_/B _09297_/X _12924_/A vssd1 vssd1 vccd1 vccd1 _09298_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_50 _15537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_61 hold363/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_72 hold597/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_83 _15145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ hold2848/X _08268_/B _08248_/X _13675_/C1 vssd1 vssd1 vccd1 vccd1 _08249_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_94 hold5952/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11260_ hold5390/X _11165_/B _11259_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _11260_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5040 _16892_/Q vssd1 vssd1 vccd1 vccd1 hold5040/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10211_ hold2918/X hold3816/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10212_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5051 _12052_/X vssd1 vssd1 vccd1 vccd1 _17174_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5062 _17197_/Q vssd1 vssd1 vccd1 vccd1 hold5062/X sky130_fd_sc_hd__dlygate4sd3_1
X_11191_ _11218_/A _11191_/B vssd1 vssd1 vccd1 vccd1 _11191_/Y sky130_fd_sc_hd__nor2_1
Xhold5073 _10819_/X vssd1 vssd1 vccd1 vccd1 _16763_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5084 _17655_/Q vssd1 vssd1 vccd1 vccd1 hold5084/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4350 _16724_/Q vssd1 vssd1 vccd1 vccd1 hold4350/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5095 _16896_/Q vssd1 vssd1 vccd1 vccd1 hold5095/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10142_ hold1984/X hold3503/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10143_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4361 _17098_/Q vssd1 vssd1 vccd1 vccd1 hold4361/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4372 _12358_/Y vssd1 vssd1 vccd1 vccd1 _17276_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4383 _11191_/Y vssd1 vssd1 vccd1 vccd1 _16887_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4394 _11763_/Y vssd1 vssd1 vccd1 vccd1 _11764_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3660 _16446_/Q vssd1 vssd1 vccd1 vccd1 hold3660/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14950_ _15165_/A _14952_/B vssd1 vssd1 vccd1 vccd1 _14950_/Y sky130_fd_sc_hd__nand2_1
XTAP_5833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10073_ _16515_/Q _10568_/B _10475_/S vssd1 vssd1 vccd1 vccd1 _10073_/X sky130_fd_sc_hd__and3_1
Xhold3671 _10216_/X vssd1 vssd1 vccd1 vccd1 _16562_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3682 _16380_/Q vssd1 vssd1 vccd1 vccd1 hold3682/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3693 _10105_/X vssd1 vssd1 vccd1 vccd1 _16525_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2970 _14309_/X vssd1 vssd1 vccd1 vccd1 _17954_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13901_ _13901_/A _13901_/B vssd1 vssd1 vccd1 vccd1 _17758_/D sky130_fd_sc_hd__and2_1
X_14881_ hold2620/X _14880_/B _14880_/Y _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14881_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2981 _18057_/Q vssd1 vssd1 vccd1 vccd1 hold2981/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2992 _14661_/X vssd1 vssd1 vccd1 vccd1 _18123_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_230_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16620_ _18146_/CLK _16620_/D vssd1 vssd1 vccd1 vccd1 _16620_/Q sky130_fd_sc_hd__dfxtp_1
X_13832_ _13832_/A _13862_/B _13862_/C vssd1 vssd1 vccd1 vccd1 _13832_/X sky130_fd_sc_hd__and3_1
XFILLER_0_199_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16551_ _18172_/CLK _16551_/D vssd1 vssd1 vccd1 vccd1 _16551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13763_ hold2017/X _17708_/Q _13883_/C vssd1 vssd1 vccd1 vccd1 _13764_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_69_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10975_ hold5205/X _11165_/B _10974_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _10975_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12714_ _12810_/A _12714_/B vssd1 vssd1 vccd1 vccd1 _17414_/D sky130_fd_sc_hd__and2_1
X_15502_ _15502_/A _15502_/B vssd1 vssd1 vccd1 vccd1 _18430_/D sky130_fd_sc_hd__and2_1
X_16482_ _18395_/CLK _16482_/D vssd1 vssd1 vccd1 vccd1 _16482_/Q sky130_fd_sc_hd__dfxtp_1
X_13694_ hold2893/X hold4129/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13695_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18221_ _18221_/CLK _18221_/D vssd1 vssd1 vccd1 vccd1 _18221_/Q sky130_fd_sc_hd__dfxtp_1
X_15433_ _15481_/A1 _15425_/X _15432_/X _15481_/B1 _18419_/Q vssd1 vssd1 vccd1 vccd1
+ _15433_/X sky130_fd_sc_hd__a32o_1
X_12645_ _12837_/A _12645_/B vssd1 vssd1 vccd1 vccd1 _17391_/D sky130_fd_sc_hd__and2_1
XFILLER_0_210_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15364_ _15364_/A _15364_/B vssd1 vssd1 vccd1 vccd1 _18412_/D sky130_fd_sc_hd__and2_1
XFILLER_0_182_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18152_ _18162_/CLK _18152_/D vssd1 vssd1 vccd1 vccd1 _18152_/Q sky130_fd_sc_hd__dfxtp_1
X_12576_ _14358_/A _12576_/B vssd1 vssd1 vccd1 vccd1 _17368_/D sky130_fd_sc_hd__and2_1
XFILLER_0_124_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17103_ _17167_/CLK _17103_/D vssd1 vssd1 vccd1 vccd1 _17103_/Q sky130_fd_sc_hd__dfxtp_1
X_14315_ hold1501/X _14326_/B _14314_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _14315_/X
+ sky130_fd_sc_hd__o211a_1
X_18083_ _18203_/CLK _18083_/D vssd1 vssd1 vccd1 vccd1 _18083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11527_ hold5703/X _12299_/B _11526_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _11527_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_230_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15295_ hold412/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15295_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17034_ _17850_/CLK _17034_/D vssd1 vssd1 vccd1 vccd1 _17034_/Q sky130_fd_sc_hd__dfxtp_1
X_14246_ _14980_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14246_/X sky130_fd_sc_hd__or2_1
Xhold309 hold309/A vssd1 vssd1 vccd1 vccd1 hold309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11458_ hold5148/X _11741_/B _11457_/X _14211_/C1 vssd1 vssd1 vccd1 vccd1 _11458_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10409_ hold1998/X hold3781/X _10595_/C vssd1 vssd1 vccd1 vccd1 _10410_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14177_ hold3061/X _14198_/B _14176_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _14177_/X
+ sky130_fd_sc_hd__o211a_1
X_11389_ hold4156/X _11771_/B _11388_/X _14131_/C1 vssd1 vssd1 vccd1 vccd1 _11389_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_221_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _13121_/X _13127_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17534_/D sky130_fd_sc_hd__o21a_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _13058_/X _16900_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13059_/X sky130_fd_sc_hd__mux2_1
X_17936_ _17936_/CLK _17936_/D vssd1 vssd1 vccd1 vccd1 _17936_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1009 _08126_/X vssd1 vssd1 vccd1 vccd1 _08127_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17867_ _17867_/CLK _17867_/D vssd1 vssd1 vccd1 vccd1 _17867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16818_ _18021_/CLK _16818_/D vssd1 vssd1 vccd1 vccd1 _16818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17798_ _17936_/CLK _17798_/D vssd1 vssd1 vccd1 vccd1 _17798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16749_ _18016_/CLK _16749_/D vssd1 vssd1 vccd1 vccd1 _16749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09221_ hold1923/X _09214_/B _09220_/X _12837_/A vssd1 vssd1 vccd1 vccd1 _09221_/X
+ sky130_fd_sc_hd__o211a_1
X_18419_ _18419_/CLK _18419_/D vssd1 vssd1 vccd1 vccd1 _18419_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09152_ _15535_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09152_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08103_ hold355/X hold307/X vssd1 vssd1 vccd1 vccd1 hold107/A sky130_fd_sc_hd__nand2b_1
X_09083_ hold1260/X _09106_/B _09082_/X _12987_/A vssd1 vssd1 vccd1 vccd1 _09083_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08034_ hold2433/X _08033_/B _08033_/Y _08143_/A vssd1 vssd1 vccd1 vccd1 _08034_/X
+ sky130_fd_sc_hd__o211a_1
Xinput70 input70/A vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_1
XFILLER_0_13_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold810 hold810/A vssd1 vssd1 vccd1 vccd1 hold810/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold821 hold821/A vssd1 vssd1 vccd1 vccd1 hold821/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold832 hold832/A vssd1 vssd1 vccd1 vccd1 hold832/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 hold843/A vssd1 vssd1 vccd1 vccd1 hold843/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold854 hold854/A vssd1 vssd1 vccd1 vccd1 hold854/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold865 hold865/A vssd1 vssd1 vccd1 vccd1 hold865/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold876 hold876/A vssd1 vssd1 vccd1 vccd1 hold876/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 hold887/A vssd1 vssd1 vccd1 vccd1 hold887/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 becStatus[0] vssd1 vssd1 vccd1 vccd1 input1/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09985_ _13070_/A _10004_/B _09984_/X _15042_/A vssd1 vssd1 vccd1 vccd1 _09985_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2200 _14237_/X vssd1 vssd1 vccd1 vccd1 _17919_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2211 _18363_/Q vssd1 vssd1 vccd1 vccd1 hold2211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08936_ _12416_/A hold721/X vssd1 vssd1 vccd1 vccd1 _16085_/D sky130_fd_sc_hd__and2_1
XTAP_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2222 _18432_/Q vssd1 vssd1 vccd1 vccd1 hold2222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2233 _14567_/X vssd1 vssd1 vccd1 vccd1 _18078_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2244 _17841_/Q vssd1 vssd1 vccd1 vccd1 hold2244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1510 _15078_/X vssd1 vssd1 vccd1 vccd1 _18323_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2255 _07825_/X vssd1 vssd1 vccd1 vccd1 _17751_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1521 _16292_/Q vssd1 vssd1 vccd1 vccd1 _09412_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2266 _12620_/X vssd1 vssd1 vccd1 vccd1 _12621_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08867_ _12410_/A hold698/X vssd1 vssd1 vccd1 vccd1 _16052_/D sky130_fd_sc_hd__and2_1
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1532 _15724_/Q vssd1 vssd1 vccd1 vccd1 hold1532/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2277 _17385_/Q vssd1 vssd1 vccd1 vccd1 hold2277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2288 _14599_/X vssd1 vssd1 vccd1 vccd1 _18093_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1543 _14927_/X vssd1 vssd1 vccd1 vccd1 _18250_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1554 _15581_/Q vssd1 vssd1 vccd1 vccd1 hold1554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2299 _08030_/X vssd1 vssd1 vccd1 vccd1 _15656_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1565 _08442_/X vssd1 vssd1 vccd1 vccd1 _15851_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1576 _18254_/Q vssd1 vssd1 vccd1 vccd1 hold1576/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07818_ hold444/A hold337/A hold509/A hold405/A vssd1 vssd1 vccd1 vccd1 _14735_/A
+ sky130_fd_sc_hd__or4bb_4
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08798_ _15491_/A hold748/X vssd1 vssd1 vccd1 vccd1 _16018_/D sky130_fd_sc_hd__and2_1
XFILLER_0_212_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1587 _17984_/Q vssd1 vssd1 vccd1 vccd1 hold1587/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1598 _18183_/Q vssd1 vssd1 vccd1 vccd1 hold1598/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_8_wb_clk_i clkbuf_6_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18443_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10760_ hold2175/X hold3828/X _11144_/C vssd1 vssd1 vccd1 vccd1 _10761_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_94_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_274_wb_clk_i clkbuf_6_51_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18150_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09419_ _07785_/Y hold5993/X _15274_/A _09418_/X vssd1 vssd1 vccd1 vccd1 _09419_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_203_wb_clk_i clkbuf_6_55_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18384_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_192_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10691_ hold2731/X hold4251/X _11171_/C vssd1 vssd1 vccd1 vccd1 _10692_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12430_ _15254_/A _12430_/B vssd1 vssd1 vccd1 vccd1 _17308_/D sky130_fd_sc_hd__and2_1
XFILLER_0_35_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12361_ _13873_/A _12361_/B vssd1 vssd1 vccd1 vccd1 _12361_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_133_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14100_ _15553_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14100_/X sky130_fd_sc_hd__or2_1
X_11312_ hold1486/X _16928_/Q _11774_/C vssd1 vssd1 vccd1 vccd1 _11313_/B sky130_fd_sc_hd__mux2_1
X_15080_ hold2137/X hold341/X _15079_/X _15146_/C1 vssd1 vssd1 vccd1 vccd1 _15080_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12292_ hold4745/X _12308_/B _12291_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _12292_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14031_ hold2121/X _14038_/B _14030_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _14031_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_240_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11243_ _18431_/Q hold3538/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11244_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11174_ _16882_/Q _11210_/B _11210_/C vssd1 vssd1 vccd1 vccd1 _11174_/X sky130_fd_sc_hd__and3_1
XTAP_6331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4180 _11530_/X vssd1 vssd1 vccd1 vccd1 _17000_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4191 hold5945/X vssd1 vssd1 vccd1 vccd1 hold5946/A sky130_fd_sc_hd__buf_4
X_10125_ _10413_/A _10125_/B vssd1 vssd1 vccd1 vccd1 _10125_/X sky130_fd_sc_hd__or2_1
XTAP_6364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15982_ _17301_/CLK _15982_/D vssd1 vssd1 vccd1 vccd1 hold529/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3490 _16725_/Q vssd1 vssd1 vccd1 vccd1 hold3490/X sky130_fd_sc_hd__buf_1
XTAP_5663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17721_ _17721_/CLK _17721_/D vssd1 vssd1 vccd1 vccd1 _17721_/Q sky130_fd_sc_hd__dfxtp_1
X_10056_ _13262_/A _10482_/A _10055_/X vssd1 vssd1 vccd1 vccd1 _10056_/Y sky130_fd_sc_hd__a21oi_1
X_14933_ hold3065/X _14952_/B _14932_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _14933_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_21_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_21_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_216_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ _17716_/CLK _17652_/D vssd1 vssd1 vccd1 vccd1 _17652_/Q sky130_fd_sc_hd__dfxtp_1
X_14864_ _14988_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14864_/X sky130_fd_sc_hd__or2_1
XFILLER_0_188_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16603_ _18225_/CLK _16603_/D vssd1 vssd1 vccd1 vccd1 _16603_/Q sky130_fd_sc_hd__dfxtp_1
X_13815_ hold5726/X _13722_/A _13814_/X vssd1 vssd1 vccd1 vccd1 _13815_/Y sky130_fd_sc_hd__a21oi_1
X_14795_ hold2064/X _14826_/B _14794_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14795_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17583_ _17608_/CLK _17583_/D vssd1 vssd1 vccd1 vccd1 _17583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16534_ _18124_/CLK _16534_/D vssd1 vssd1 vccd1 vccd1 _16534_/Q sky130_fd_sc_hd__dfxtp_1
X_13746_ _13752_/A _13746_/B vssd1 vssd1 vccd1 vccd1 _13746_/X sky130_fd_sc_hd__or2_1
X_10958_ hold2975/X hold4143/X _11726_/C vssd1 vssd1 vccd1 vccd1 _10959_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16465_ _18378_/CLK _16465_/D vssd1 vssd1 vccd1 vccd1 _16465_/Q sky130_fd_sc_hd__dfxtp_1
X_13677_ _13776_/A _13677_/B vssd1 vssd1 vccd1 vccd1 _13677_/X sky130_fd_sc_hd__or2_1
X_10889_ hold1406/X hold4945/X _11171_/C vssd1 vssd1 vccd1 vccd1 _10890_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_128_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18204_ _18236_/CLK _18204_/D vssd1 vssd1 vccd1 vccd1 _18204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15416_ _17317_/Q _09357_/A _09392_/A hold501/X vssd1 vssd1 vccd1 vccd1 _15416_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12628_ hold1087/X _17387_/Q _12850_/S vssd1 vssd1 vccd1 vccd1 _12628_/X sky130_fd_sc_hd__mux2_1
X_16396_ _18349_/CLK _16396_/D vssd1 vssd1 vccd1 vccd1 _16396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15347_ hold864/X _09357_/A _09386_/D hold735/X _15346_/X vssd1 vssd1 vccd1 vccd1
+ _15352_/B sky130_fd_sc_hd__a221o_1
X_18135_ _18232_/CLK _18135_/D vssd1 vssd1 vccd1 vccd1 _18135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12559_ hold3055/X _17364_/Q _12925_/S vssd1 vssd1 vccd1 vccd1 _12559_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_227_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5809 _17725_/Q vssd1 vssd1 vccd1 vccd1 hold5809/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15278_ hold769/X _15484_/A2 _09392_/D hold805/X vssd1 vssd1 vccd1 vccd1 _15278_/X
+ sky130_fd_sc_hd__a22o_1
X_18066_ _18066_/CLK _18066_/D vssd1 vssd1 vccd1 vccd1 _18066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold106 hold306/X vssd1 vssd1 vccd1 vccd1 hold307/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold117 hold117/A vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 data_in[2] vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 hold139/A vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ hold1746/X _14216_/Y _14228_/X _14354_/A vssd1 vssd1 vccd1 vccd1 _14229_/X
+ sky130_fd_sc_hd__o211a_1
X_17017_ _17865_/CLK _17017_/D vssd1 vssd1 vccd1 vccd1 _17017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_78_wb_clk_i clkbuf_6_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17512_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_6_60_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_60_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout608 _15488_/A2 vssd1 vssd1 vccd1 vccd1 _09392_/C sky130_fd_sc_hd__buf_6
Xfanout619 _09354_/Y vssd1 vssd1 vccd1 vccd1 _09357_/A sky130_fd_sc_hd__buf_6
XFILLER_0_238_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09770_ hold1031/X hold3228/X _10040_/C vssd1 vssd1 vccd1 vccd1 _09771_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08721_ hold87/X hold529/X _08721_/S vssd1 vssd1 vccd1 vccd1 hold530/A sky130_fd_sc_hd__mux2_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17919_ _18307_/CLK _17919_/D vssd1 vssd1 vccd1 vccd1 _17919_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08652_ _12412_/A _08652_/B vssd1 vssd1 vccd1 vccd1 _15948_/D sky130_fd_sc_hd__and2_1
XFILLER_0_90_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08583_ _15324_/A _08583_/B vssd1 vssd1 vccd1 vccd1 _15915_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09204_ _15533_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09204_/X sky130_fd_sc_hd__or2_1
XFILLER_0_45_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09135_ hold2371/X _09177_/A2 _09134_/X _12864_/A vssd1 vssd1 vccd1 vccd1 _09135_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09066_ _15182_/A hold363/X vssd1 vssd1 vccd1 vccd1 _09066_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08017_ _15531_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08017_/X sky130_fd_sc_hd__or2_1
Xhold640 hold640/A vssd1 vssd1 vccd1 vccd1 hold640/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold651 hold651/A vssd1 vssd1 vccd1 vccd1 hold651/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 hold662/A vssd1 vssd1 vccd1 vccd1 hold662/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 hold74/X vssd1 vssd1 vccd1 vccd1 hold673/X sky130_fd_sc_hd__buf_4
Xhold684 hold684/A vssd1 vssd1 vccd1 vccd1 hold684/X sky130_fd_sc_hd__buf_4
Xhold695 hold695/A vssd1 vssd1 vccd1 vccd1 hold695/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ hold2306/X _16480_/Q _10067_/C vssd1 vssd1 vccd1 vccd1 _09969_/B sky130_fd_sc_hd__mux2_1
Xhold2030 _14131_/X vssd1 vssd1 vccd1 vccd1 _17869_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2041 _15880_/Q vssd1 vssd1 vccd1 vccd1 hold2041/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_08919_ _09047_/A _08919_/B vssd1 vssd1 vccd1 vccd1 _16077_/D sky130_fd_sc_hd__and2_1
Xhold2052 _14849_/X vssd1 vssd1 vccd1 vccd1 _18213_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2063 _14029_/X vssd1 vssd1 vccd1 vccd1 _17820_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09899_ _18370_/Q _16457_/Q _10964_/S vssd1 vssd1 vccd1 vccd1 _09900_/B sky130_fd_sc_hd__mux2_1
Xhold2074 _14671_/X vssd1 vssd1 vccd1 vccd1 _18128_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2085 _18238_/Q vssd1 vssd1 vccd1 vccd1 hold2085/X sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1340 _15874_/Q vssd1 vssd1 vccd1 vccd1 hold1340/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2096 _18206_/Q vssd1 vssd1 vccd1 vccd1 hold2096/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1351 _15528_/X vssd1 vssd1 vccd1 vccd1 _18442_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11930_ hold2662/X _17134_/Q _12227_/S vssd1 vssd1 vccd1 vccd1 _11931_/B sky130_fd_sc_hd__mux2_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1362 _17899_/Q vssd1 vssd1 vccd1 vccd1 hold1362/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1373 _08420_/X vssd1 vssd1 vccd1 vccd1 _15840_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_455_wb_clk_i clkbuf_6_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17427_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1384 _16288_/Q vssd1 vssd1 vccd1 vccd1 _09404_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1395 _15855_/Q vssd1 vssd1 vccd1 vccd1 hold1395/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11861_ hold2622/X _17111_/Q _12371_/C vssd1 vssd1 vccd1 vccd1 _11862_/B sky130_fd_sc_hd__mux2_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ hold4129/X _13880_/B _13599_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13600_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _11661_/A _10812_/B vssd1 vssd1 vccd1 vccd1 _10812_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14580_ _15189_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14580_/X sky130_fd_sc_hd__or2_1
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _17088_/Q _11792_/B _12335_/C vssd1 vssd1 vccd1 vccd1 _11792_/X sky130_fd_sc_hd__and3_1
XFILLER_0_95_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13531_ hold4689/X _13829_/B _13530_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13531_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10743_ _11694_/A _10743_/B vssd1 vssd1 vccd1 vccd1 _10743_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16250_ _17429_/CLK _16250_/D vssd1 vssd1 vccd1 vccd1 _16250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13462_ hold5643/X _13880_/B _13461_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _13462_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10674_ _11136_/A _10674_/B vssd1 vssd1 vccd1 vccd1 _10674_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15201_ _15201_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15201_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12413_ hold185/X hold800/X _12441_/S vssd1 vssd1 vccd1 vccd1 hold801/A sky130_fd_sc_hd__mux2_1
XFILLER_0_51_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16181_ _17464_/CLK _16181_/D vssd1 vssd1 vccd1 vccd1 _16181_/Q sky130_fd_sc_hd__dfxtp_1
X_13393_ hold5466/X _13871_/B _13392_/X _13675_/C1 vssd1 vssd1 vccd1 vccd1 _13393_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15132_ hold1479/X _15165_/B _15131_/X _15048_/A vssd1 vssd1 vccd1 vccd1 _15132_/X
+ sky130_fd_sc_hd__o211a_1
X_12344_ _17272_/Q _12374_/B _12371_/C vssd1 vssd1 vccd1 vccd1 _12344_/X sky130_fd_sc_hd__and3_1
XFILLER_0_50_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15063_ _15225_/A hold1470/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15064_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12275_ hold1554/X _17249_/Q _13748_/S vssd1 vssd1 vccd1 vccd1 _12276_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14014_ _15521_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14014_/X sky130_fd_sc_hd__or2_1
X_11226_ hold4278/X _11670_/A _11225_/X vssd1 vssd1 vccd1 vccd1 _11226_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11157_ hold3479/X _11067_/A _11156_/X vssd1 vssd1 vccd1 vccd1 _11157_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10108_ hold4475/X _10628_/B _10107_/X _14863_/C1 vssd1 vssd1 vccd1 vccd1 _10108_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15965_ _17284_/CLK _15965_/D vssd1 vssd1 vccd1 vccd1 hold414/A sky130_fd_sc_hd__dfxtp_1
X_11088_ _11088_/A _11088_/B vssd1 vssd1 vccd1 vccd1 _11088_/X sky130_fd_sc_hd__or2_1
XTAP_5471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17704_ _17740_/CLK _17704_/D vssd1 vssd1 vccd1 vccd1 _17704_/Q sky130_fd_sc_hd__dfxtp_1
X_10039_ _10603_/A _10039_/B vssd1 vssd1 vccd1 vccd1 _10039_/Y sky130_fd_sc_hd__nor2_1
XTAP_5493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14916_ _15185_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14916_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_196_wb_clk_i clkbuf_6_53_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18382_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15896_ _16147_/CLK _15896_/D vssd1 vssd1 vccd1 vccd1 _15896_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17635_ _17731_/CLK _17635_/D vssd1 vssd1 vccd1 vccd1 _17635_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_125_wb_clk_i clkbuf_6_22_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18412_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14847_ hold2025/X _14880_/B _14846_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14847_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_216_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17566_ _17718_/CLK _17566_/D vssd1 vssd1 vccd1 vccd1 _17566_/Q sky130_fd_sc_hd__dfxtp_1
X_14778_ _15225_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14778_/X sky130_fd_sc_hd__or2_1
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16517_ _18235_/CLK _16517_/D vssd1 vssd1 vccd1 vccd1 _16517_/Q sky130_fd_sc_hd__dfxtp_1
X_13729_ _13823_/A _13795_/A2 _13728_/X _13729_/C1 vssd1 vssd1 vccd1 vccd1 _13729_/X
+ sky130_fd_sc_hd__o211a_1
X_17497_ _17499_/CLK _17497_/D vssd1 vssd1 vccd1 vccd1 _17497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16448_ _16480_/CLK _16448_/D vssd1 vssd1 vccd1 vccd1 _16448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16379_ _18346_/CLK _16379_/D vssd1 vssd1 vccd1 vccd1 _16379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18118_ _18150_/CLK _18118_/D vssd1 vssd1 vccd1 vccd1 _18118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5606 _13696_/X vssd1 vssd1 vccd1 vccd1 _17685_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5617 _10408_/X vssd1 vssd1 vccd1 vccd1 _16626_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5628 _17671_/Q vssd1 vssd1 vccd1 vccd1 hold5628/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5639 _16941_/Q vssd1 vssd1 vccd1 vccd1 hold5639/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4905 _16748_/Q vssd1 vssd1 vccd1 vccd1 hold4905/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18049_ _18049_/CLK _18049_/D vssd1 vssd1 vccd1 vccd1 _18049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4916 _12058_/X vssd1 vssd1 vccd1 vccd1 _17176_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4927 _17179_/Q vssd1 vssd1 vccd1 vccd1 hold4927/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4938 _12199_/X vssd1 vssd1 vccd1 vccd1 _17223_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4949 _16790_/Q vssd1 vssd1 vccd1 vccd1 hold4949/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout405 _14340_/X vssd1 vssd1 vccd1 vccd1 _14391_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_240_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout416 _14108_/Y vssd1 vssd1 vccd1 vccd1 _14148_/B sky130_fd_sc_hd__buf_8
X_09822_ _09933_/A _09822_/B vssd1 vssd1 vccd1 vccd1 _09822_/X sky130_fd_sc_hd__or2_1
Xfanout427 hold296/X vssd1 vssd1 vccd1 vccd1 hold297/A sky130_fd_sc_hd__clkbuf_2
Xfanout438 _13721_/S vssd1 vssd1 vccd1 vccd1 _12293_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_225_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout449 fanout485/X vssd1 vssd1 vccd1 vccd1 _11717_/C sky130_fd_sc_hd__clkbuf_8
X_09753_ _11109_/A _09753_/B vssd1 vssd1 vccd1 vccd1 _09753_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08704_ _12416_/A _08704_/B vssd1 vssd1 vccd1 vccd1 _15973_/D sky130_fd_sc_hd__and2_1
XFILLER_0_240_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09684_ _10560_/A _09684_/B vssd1 vssd1 vccd1 vccd1 _09684_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08635_ hold245/X hold539/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08636_/B sky130_fd_sc_hd__mux2_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08566_ hold254/X hold694/X _08592_/S vssd1 vssd1 vccd1 vccd1 _08567_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08497_ hold1497/X _08486_/B _08496_/X _08347_/A vssd1 vssd1 vccd1 vccd1 _08497_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09118_ _15559_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09118_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10390_ hold3666/X _10625_/B _10389_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10390_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09049_ _09057_/A hold144/X vssd1 vssd1 vccd1 vccd1 _16141_/D sky130_fd_sc_hd__and2_1
XFILLER_0_27_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12060_ _12255_/A _12060_/B vssd1 vssd1 vccd1 vccd1 _12060_/X sky130_fd_sc_hd__or2_1
Xhold470 hold470/A vssd1 vssd1 vccd1 vccd1 hold470/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold481 hold481/A vssd1 vssd1 vccd1 vccd1 hold481/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold492 hold492/A vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ hold5219/X _11171_/B _11010_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _11011_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ hold3232/X _12961_/X _12971_/S vssd1 vssd1 vccd1 vccd1 _12963_/B sky130_fd_sc_hd__mux2_1
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _17733_/CLK _15750_/D vssd1 vssd1 vccd1 vccd1 _15750_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1170 _15620_/Q vssd1 vssd1 vccd1 vccd1 hold1170/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ hold2891/X _14720_/B _14700_/X _14769_/C1 vssd1 vssd1 vccd1 vccd1 _14701_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1181 hold690/X vssd1 vssd1 vccd1 vccd1 input41/A sky130_fd_sc_hd__dlygate4sd3_1
X_11913_ _13716_/A _11913_/B vssd1 vssd1 vccd1 vccd1 _11913_/X sky130_fd_sc_hd__or2_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1192 input37/X vssd1 vssd1 vccd1 vccd1 hold926/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15681_ _17843_/CLK _15681_/D vssd1 vssd1 vccd1 vccd1 _15681_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ hold3159/X _12892_/X _12905_/S vssd1 vssd1 vccd1 vccd1 _12893_/X sky130_fd_sc_hd__mux2_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17420_ _17661_/CLK _17420_/D vssd1 vssd1 vccd1 vccd1 _17420_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ hold911/X _14678_/B vssd1 vssd1 vccd1 vccd1 _14632_/X sky130_fd_sc_hd__or2_1
X_11844_ _12234_/A _11844_/B vssd1 vssd1 vccd1 vccd1 _11844_/X sky130_fd_sc_hd__or2_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14563_ hold911/X _14557_/Y _14562_/X _15218_/C1 vssd1 vssd1 vccd1 vccd1 hold912/A
+ sky130_fd_sc_hd__o211a_1
X_17351_ _17512_/CLK _17351_/D vssd1 vssd1 vccd1 vccd1 _17351_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11775_ hold3465/X _11697_/A _11774_/X vssd1 vssd1 vccd1 vccd1 _11775_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_200_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16302_ _16319_/CLK hold706/X vssd1 vssd1 vccd1 vccd1 _16302_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10726_ hold4907/X _11204_/B _10725_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _10726_/X
+ sky130_fd_sc_hd__o211a_1
X_13514_ hold3016/X hold4831/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13515_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_166_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14494_ hold1517/X _14487_/B _14493_/X _14354_/A vssd1 vssd1 vccd1 vccd1 _14494_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17282_ _17617_/CLK _17282_/D vssd1 vssd1 vccd1 vccd1 _17282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13445_ hold1045/X _17602_/Q _13829_/C vssd1 vssd1 vccd1 vccd1 _13446_/B sky130_fd_sc_hd__mux2_1
X_16233_ _17754_/CLK _16233_/D vssd1 vssd1 vccd1 vccd1 hold917/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10657_ hold4799/X _11153_/B _10656_/X _14552_/C1 vssd1 vssd1 vccd1 vccd1 _10657_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16164_ _17499_/CLK _16164_/D vssd1 vssd1 vccd1 vccd1 _16164_/Q sky130_fd_sc_hd__dfxtp_1
X_13376_ hold1760/X hold4408/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13377_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10588_ _10651_/A _10588_/B vssd1 vssd1 vccd1 vccd1 _16686_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_51_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15115_ _15169_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15115_/X sky130_fd_sc_hd__or2_1
XFILLER_0_121_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12327_ hold4290/X _13482_/A _12326_/X vssd1 vssd1 vccd1 vccd1 _12327_/Y sky130_fd_sc_hd__a21oi_1
X_16095_ _18419_/CLK _16095_/D vssd1 vssd1 vccd1 vccd1 _16095_/Q sky130_fd_sc_hd__dfxtp_1
X_15046_ _15473_/A _15046_/B vssd1 vssd1 vccd1 vccd1 _18308_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12258_ _13314_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _12258_/X sky130_fd_sc_hd__or2_1
X_11209_ _12331_/A _11209_/B vssd1 vssd1 vccd1 vccd1 _11209_/Y sky130_fd_sc_hd__nor2_1
X_12189_ _12285_/A _12189_/B vssd1 vssd1 vccd1 vccd1 _12189_/X sky130_fd_sc_hd__or2_1
XFILLER_0_208_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_377_wb_clk_i clkbuf_6_32_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17742_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_236_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16997_ _17877_/CLK _16997_/D vssd1 vssd1 vccd1 vccd1 _16997_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_306_wb_clk_i clkbuf_6_45_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17871_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_183_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15948_ _17295_/CLK _15948_/D vssd1 vssd1 vccd1 vccd1 hold867/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15879_ _17590_/CLK _15879_/D vssd1 vssd1 vccd1 vccd1 _15879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08420_ hold1372/X _08442_/A2 _08419_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _08420_/X
+ sky130_fd_sc_hd__o211a_1
X_17618_ _17653_/CLK _17618_/D vssd1 vssd1 vccd1 vccd1 _17618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08351_ _08351_/A hold964/X vssd1 vssd1 vccd1 vccd1 _15807_/D sky130_fd_sc_hd__and2_1
X_17549_ _18217_/CLK _17549_/D vssd1 vssd1 vccd1 vccd1 _17549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08282_ hold444/A hold337/X hold509/A hold405/A vssd1 vssd1 vccd1 vccd1 hold338/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_73_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_93_wb_clk_i clkbuf_6_19_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16323_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold6104 la_data_in[25] vssd1 vssd1 vccd1 vccd1 hold576/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6115 _16534_/Q vssd1 vssd1 vccd1 vccd1 hold6115/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6126 _16521_/Q vssd1 vssd1 vccd1 vccd1 hold6126/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_22_wb_clk_i clkbuf_6_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17481_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5403 _13771_/X vssd1 vssd1 vccd1 vccd1 _17710_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5414 _17738_/Q vssd1 vssd1 vccd1 vccd1 hold5414/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5425 _10522_/X vssd1 vssd1 vccd1 vccd1 _16664_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5436 _17084_/Q vssd1 vssd1 vccd1 vccd1 hold5436/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4702 _11035_/X vssd1 vssd1 vccd1 vccd1 _16835_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5447 _10672_/X vssd1 vssd1 vccd1 vccd1 _16714_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4713 _16422_/Q vssd1 vssd1 vccd1 vccd1 hold4713/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5458 _17262_/Q vssd1 vssd1 vccd1 vccd1 hold5458/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5469 _12145_/X vssd1 vssd1 vccd1 vccd1 _17205_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4724 _12331_/Y vssd1 vssd1 vccd1 vccd1 _17267_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4735 _16492_/Q vssd1 vssd1 vccd1 vccd1 hold4735/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4746 _12292_/X vssd1 vssd1 vccd1 vccd1 _17254_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4757 _13621_/X vssd1 vssd1 vccd1 vccd1 _17660_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4768 _16460_/Q vssd1 vssd1 vccd1 vccd1 hold4768/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout202 _11210_/B vssd1 vssd1 vccd1 vccd1 _11195_/B sky130_fd_sc_hd__clkbuf_8
Xhold4779 _17696_/Q vssd1 vssd1 vccd1 vccd1 hold4779/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout213 _11201_/B vssd1 vssd1 vccd1 vccd1 _11162_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout224 _10070_/B vssd1 vssd1 vccd1 vccd1 _11186_/B sky130_fd_sc_hd__buf_4
Xfanout235 _10067_/B vssd1 vssd1 vccd1 vccd1 _10568_/B sky130_fd_sc_hd__clkbuf_8
Xfanout246 _10634_/B vssd1 vssd1 vccd1 vccd1 _10637_/B sky130_fd_sc_hd__buf_4
XFILLER_0_201_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09805_ hold4720/X _10028_/B _09804_/X _15042_/A vssd1 vssd1 vccd1 vccd1 _09805_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout257 _12216_/A vssd1 vssd1 vccd1 vccd1 _13314_/A sky130_fd_sc_hd__buf_4
XFILLER_0_96_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout268 _11556_/A vssd1 vssd1 vccd1 vccd1 _11553_/A sky130_fd_sc_hd__clkbuf_4
Xfanout279 _13599_/A vssd1 vssd1 vccd1 vccd1 _13788_/A sky130_fd_sc_hd__buf_4
X_07997_ hold915/X _08045_/B vssd1 vssd1 vccd1 vccd1 _07997_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_236_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09736_ hold4839/X _11171_/B _09735_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _09736_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09667_ hold3650/X _10046_/B _09666_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09667_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08618_ _12410_/A hold860/X vssd1 vssd1 vccd1 vccd1 _15931_/D sky130_fd_sc_hd__and2_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ hold5277/X _09992_/B _09597_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _09598_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08549_ _12438_/A _08549_/B vssd1 vssd1 vccd1 vccd1 _15898_/D sky130_fd_sc_hd__and2_1
XFILLER_0_155_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11560_ hold5195/X _11753_/B _11559_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _11560_/X
+ sky130_fd_sc_hd__o211a_1
X_10511_ hold2261/X _16661_/Q _10637_/C vssd1 vssd1 vccd1 vccd1 _10512_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_181_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11491_ hold5221/X _12317_/B _11490_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11491_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13230_ _13230_/A _13294_/B vssd1 vssd1 vccd1 vccd1 _13230_/X sky130_fd_sc_hd__or2_1
X_10442_ hold1495/X _16638_/Q _10634_/C vssd1 vssd1 vccd1 vccd1 _10443_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_162_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13161_ _13161_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13161_/X sky130_fd_sc_hd__and2_1
X_10373_ hold1785/X hold3259/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10374_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12112_ hold4811/X _12293_/B _12111_/X _12822_/A vssd1 vssd1 vccd1 vccd1 _12112_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5970 _17752_/Q vssd1 vssd1 vccd1 vccd1 hold5970/X sky130_fd_sc_hd__dlygate4sd3_1
X_13092_ hold3508/X _13091_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13092_/X sky130_fd_sc_hd__mux2_2
Xhold5981 _09483_/X vssd1 vssd1 vccd1 vccd1 hold5981/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5992 _16320_/Q vssd1 vssd1 vccd1 vccd1 _09477_/A sky130_fd_sc_hd__dlygate4sd3_1
X_12043_ hold5671/X _12329_/B _12042_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _12043_/X
+ sky130_fd_sc_hd__o211a_1
X_16920_ _17871_/CLK _16920_/D vssd1 vssd1 vccd1 vccd1 _16920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_236_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_219_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16851_ _18054_/CLK _16851_/D vssd1 vssd1 vccd1 vccd1 _16851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout780 fanout791/X vssd1 vssd1 vccd1 vccd1 _13917_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout791 fanout843/X vssd1 vssd1 vccd1 vccd1 fanout791/X sky130_fd_sc_hd__buf_8
X_15802_ _17617_/CLK _15802_/D vssd1 vssd1 vccd1 vccd1 _15802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16782_ _17985_/CLK _16782_/D vssd1 vssd1 vccd1 vccd1 _16782_/Q sky130_fd_sc_hd__dfxtp_1
X_13994_ _14960_/A _13994_/B vssd1 vssd1 vccd1 vccd1 _13994_/X sky130_fd_sc_hd__or2_1
XFILLER_0_233_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15733_ _17672_/CLK _15733_/D vssd1 vssd1 vccd1 vccd1 _15733_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12945_ _12987_/A _12945_/B vssd1 vssd1 vccd1 vccd1 _17491_/D sky130_fd_sc_hd__and2_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18452_ _18452_/CLK _18452_/D vssd1 vssd1 vccd1 vccd1 _18452_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _17272_/CLK hold970/X vssd1 vssd1 vccd1 vccd1 hold969/A sky130_fd_sc_hd__dfxtp_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _12888_/A _12876_/B vssd1 vssd1 vccd1 vccd1 _17468_/D sky130_fd_sc_hd__and2_1
XFILLER_0_158_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17403_ _18457_/CLK _17403_/D vssd1 vssd1 vccd1 vccd1 _17403_/Q sky130_fd_sc_hd__dfxtp_1
X_14615_ hold1764/X _14610_/B _14614_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14615_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _18383_/CLK _18383_/D vssd1 vssd1 vccd1 vccd1 _18383_/Q sky130_fd_sc_hd__dfxtp_1
X_11827_ hold5559/X _12305_/B _11826_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _11827_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _17221_/CLK _15595_/D vssd1 vssd1 vccd1 vccd1 _15595_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _18410_/CLK hold63/X vssd1 vssd1 vccd1 vccd1 _17334_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11758_ _12331_/A _11758_/B vssd1 vssd1 vccd1 vccd1 _11758_/Y sky130_fd_sc_hd__nor2_1
X_14546_ hold1951/X _14541_/B _14545_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _14546_/X
+ sky130_fd_sc_hd__o211a_1
X_10709_ hold2623/X _16727_/Q _11183_/C vssd1 vssd1 vccd1 vccd1 _10710_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17265_ _17900_/CLK _17265_/D vssd1 vssd1 vccd1 vccd1 _17265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11689_ hold5685/X _12329_/B _11688_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _11689_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14477_ _14477_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14477_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16216_ _17724_/CLK _16216_/D vssd1 vssd1 vccd1 vccd1 _16216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13428_ _13716_/A _13428_/B vssd1 vssd1 vccd1 vccd1 _13428_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17196_ _17259_/CLK _17196_/D vssd1 vssd1 vccd1 vccd1 _17196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16147_ _16147_/CLK _16147_/D vssd1 vssd1 vccd1 vccd1 hold459/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13359_ _13776_/A _13359_/B vssd1 vssd1 vccd1 vccd1 _13359_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4009 _16650_/Q vssd1 vssd1 vccd1 vccd1 hold4009/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3308 _16631_/Q vssd1 vssd1 vccd1 vccd1 hold3308/X sky130_fd_sc_hd__dlygate4sd3_1
X_16078_ _17309_/CLK _16078_/D vssd1 vssd1 vccd1 vccd1 _16078_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3319 _12857_/X vssd1 vssd1 vccd1 vccd1 _12858_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07920_ _15543_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _07920_/Y sky130_fd_sc_hd__nand2_1
X_15029_ _15191_/A hold2297/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15030_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2607 _17867_/Q vssd1 vssd1 vccd1 vccd1 hold2607/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2618 _15631_/Q vssd1 vssd1 vccd1 vccd1 hold2618/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2629 _18014_/Q vssd1 vssd1 vccd1 vccd1 hold2629/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1906 _14629_/X vssd1 vssd1 vccd1 vccd1 _18107_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07851_ _15529_/A _07871_/B vssd1 vssd1 vccd1 vccd1 _07851_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_140_wb_clk_i clkbuf_6_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18308_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1917 _18298_/Q vssd1 vssd1 vccd1 vccd1 hold1917/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1928 _14396_/X vssd1 vssd1 vccd1 vccd1 _17996_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1939 _17920_/Q vssd1 vssd1 vccd1 vccd1 hold1939/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput2 input2/A vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07782_ hold597/X vssd1 vssd1 vccd1 vccd1 _07782_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_223_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_233_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09521_ hold1835/X _13118_/A _10025_/C vssd1 vssd1 vccd1 vccd1 _09522_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_224_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09452_ _09456_/C _09456_/D _09456_/B vssd1 vssd1 vccd1 vccd1 _09454_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08403_ _15517_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08403_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_231_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09383_ _15480_/A _09383_/B _09383_/C _09383_/D vssd1 vssd1 vccd1 vccd1 _09383_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_188_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08334_ hold1215/X _08323_/B _08333_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _08334_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08265_ hold2466/X _08268_/B _08264_/Y _13795_/C1 vssd1 vssd1 vccd1 vccd1 _08265_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08196_ hold2822/X _08213_/B _08195_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _08196_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5200 _11614_/X vssd1 vssd1 vccd1 vccd1 _17028_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5211 _17646_/Q vssd1 vssd1 vccd1 vccd1 hold5211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5222 _11491_/X vssd1 vssd1 vccd1 vccd1 _16987_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5233 _17704_/Q vssd1 vssd1 vccd1 vccd1 hold5233/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_299_wb_clk_i clkbuf_6_38_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17891_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5244 _10684_/X vssd1 vssd1 vccd1 vccd1 _16718_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4510 _09718_/X vssd1 vssd1 vccd1 vccd1 _16396_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5255 _17251_/Q vssd1 vssd1 vccd1 vccd1 hold5255/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4521 _16564_/Q vssd1 vssd1 vccd1 vccd1 hold4521/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5266 _13741_/X vssd1 vssd1 vccd1 vccd1 _17700_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5277 _16388_/Q vssd1 vssd1 vccd1 vccd1 hold5277/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4532 _11193_/Y vssd1 vssd1 vccd1 vccd1 _11194_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_228_wb_clk_i clkbuf_6_63_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18227_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_219_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4543 _16578_/Q vssd1 vssd1 vccd1 vccd1 hold4543/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5288 _13762_/X vssd1 vssd1 vccd1 vccd1 _17707_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4554 _17491_/Q vssd1 vssd1 vccd1 vccd1 hold4554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5299 _17011_/Q vssd1 vssd1 vccd1 vccd1 hold5299/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3820 _16801_/Q vssd1 vssd1 vccd1 vccd1 hold3820/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4565 _17132_/Q vssd1 vssd1 vccd1 vccd1 hold4565/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3831 _10441_/X vssd1 vssd1 vccd1 vccd1 _16637_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4576 _10693_/X vssd1 vssd1 vccd1 vccd1 _16721_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3842 _16775_/Q vssd1 vssd1 vccd1 vccd1 hold3842/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4587 _17196_/Q vssd1 vssd1 vccd1 vccd1 hold4587/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3853 _10519_/X vssd1 vssd1 vccd1 vccd1 _16663_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4598 _17506_/Q vssd1 vssd1 vccd1 vccd1 hold4598/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3864 _16417_/Q vssd1 vssd1 vccd1 vccd1 hold3864/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3875 _10081_/X vssd1 vssd1 vccd1 vccd1 _16517_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3886 _16512_/Q vssd1 vssd1 vccd1 vccd1 hold3886/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3897 _16648_/Q vssd1 vssd1 vccd1 vccd1 hold3897/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09719_ hold1621/X _16397_/Q _10031_/C vssd1 vssd1 vccd1 vccd1 _09720_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_199_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10991_ hold1688/X hold3933/X _11183_/C vssd1 vssd1 vccd1 vccd1 _10992_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _16241_/Q hold3156/X _12811_/S vssd1 vssd1 vccd1 vccd1 _12730_/X sky130_fd_sc_hd__mux2_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ hold2802/X _17398_/Q _12850_/S vssd1 vssd1 vccd1 vccd1 _12661_/X sky130_fd_sc_hd__mux2_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14400_ hold2013/X _14446_/A2 _14399_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _14400_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11612_ hold2481/X _17028_/Q _12317_/C vssd1 vssd1 vccd1 vccd1 _11613_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_203_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ hold767/X _09367_/A _09392_/A hold802/X vssd1 vssd1 vccd1 vccd1 _15380_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12592_ hold961/X _17375_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _12592_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_203_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14331_ hold1592/X _14326_/B _14330_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _14331_/X
+ sky130_fd_sc_hd__o211a_1
X_11543_ hold2071/X _17005_/Q _11738_/C vssd1 vssd1 vccd1 vccd1 _11544_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17050_ _17834_/CLK _17050_/D vssd1 vssd1 vccd1 vccd1 _17050_/Q sky130_fd_sc_hd__dfxtp_1
X_14262_ _14477_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14262_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11474_ hold2785/X hold4883/X _11660_/S vssd1 vssd1 vccd1 vccd1 _11475_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13213_ _13212_/X hold3206/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13213_/X sky130_fd_sc_hd__mux2_2
X_16001_ _18408_/CLK _16001_/D vssd1 vssd1 vccd1 vccd1 hold699/A sky130_fd_sc_hd__dfxtp_1
X_10425_ _11103_/A _10425_/B vssd1 vssd1 vccd1 vccd1 _10425_/X sky130_fd_sc_hd__or2_1
XFILLER_0_61_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14193_ hold1362/X _14198_/B _14192_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _14193_/X
+ sky130_fd_sc_hd__o211a_1
X_13144_ _13137_/X _13143_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17536_/D sky130_fd_sc_hd__o21a_1
X_10356_ _10551_/A _10356_/B vssd1 vssd1 vccd1 vccd1 _10356_/X sky130_fd_sc_hd__or2_1
XFILLER_0_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17952_ _18307_/CLK _17952_/D vssd1 vssd1 vccd1 vccd1 _17952_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ _13074_/X hold5990/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13075_/X sky130_fd_sc_hd__mux2_1
X_10287_ _11091_/A _10287_/B vssd1 vssd1 vccd1 vccd1 _10287_/X sky130_fd_sc_hd__or2_1
XFILLER_0_100_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12026_ hold1686/X hold3702/X _12227_/S vssd1 vssd1 vccd1 vccd1 _12027_/B sky130_fd_sc_hd__mux2_1
X_16903_ _17877_/CLK _16903_/D vssd1 vssd1 vccd1 vccd1 _16903_/Q sky130_fd_sc_hd__dfxtp_1
X_17883_ _17883_/CLK _17883_/D vssd1 vssd1 vccd1 vccd1 _17883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16834_ _18069_/CLK _16834_/D vssd1 vssd1 vccd1 vccd1 _16834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16765_ _17968_/CLK _16765_/D vssd1 vssd1 vccd1 vccd1 _16765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13977_ hold1783/X _13986_/B _13976_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _13977_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15716_ _17260_/CLK _15716_/D vssd1 vssd1 vccd1 vccd1 _15716_/Q sky130_fd_sc_hd__dfxtp_1
X_12928_ hold1301/X _17487_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12928_/X sky130_fd_sc_hd__mux2_1
X_16696_ _18226_/CLK _16696_/D vssd1 vssd1 vccd1 vccd1 _16696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18435_ _18437_/CLK _18435_/D vssd1 vssd1 vccd1 vccd1 _18435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15647_ _17127_/CLK _15647_/D vssd1 vssd1 vccd1 vccd1 _15647_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ hold2371/X hold3353/X _12916_/S vssd1 vssd1 vccd1 vccd1 _12859_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_189_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18366_ _18370_/CLK _18366_/D vssd1 vssd1 vccd1 vccd1 _18366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15578_ _17584_/CLK _15578_/D vssd1 vssd1 vccd1 vccd1 _15578_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17317_ _17319_/CLK hold135/X vssd1 vssd1 vccd1 vccd1 _17317_/Q sky130_fd_sc_hd__dfxtp_1
X_14529_ _14529_/A _14543_/B vssd1 vssd1 vccd1 vccd1 _14529_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18297_ _18394_/CLK _18297_/D vssd1 vssd1 vccd1 vccd1 _18297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08050_ _14164_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08050_/X sky130_fd_sc_hd__or2_1
X_17248_ _17280_/CLK _17248_/D vssd1 vssd1 vccd1 vccd1 _17248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17179_ _17590_/CLK _17179_/D vssd1 vssd1 vccd1 vccd1 _17179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_392_wb_clk_i clkbuf_6_36_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17774_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_321_wb_clk_i clkbuf_6_46_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17840_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3105 _14251_/X vssd1 vssd1 vccd1 vccd1 _17926_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3116 _15569_/Q vssd1 vssd1 vccd1 vccd1 hold3116/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3127 _17451_/Q vssd1 vssd1 vccd1 vccd1 hold3127/X sky130_fd_sc_hd__dlygate4sd3_1
X_08952_ _15244_/A _08952_/B vssd1 vssd1 vccd1 vccd1 _16093_/D sky130_fd_sc_hd__and2_1
Xhold3138 _12629_/X vssd1 vssd1 vccd1 vccd1 _12630_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2404 _17514_/Q vssd1 vssd1 vccd1 vccd1 hold2404/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3149 _17460_/Q vssd1 vssd1 vccd1 vccd1 hold3149/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2415 _08012_/X vssd1 vssd1 vccd1 vccd1 _15647_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07903_ hold3074/X _07924_/B _07902_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _07903_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2426 _15567_/Q vssd1 vssd1 vccd1 vccd1 hold2426/X sky130_fd_sc_hd__dlygate4sd3_1
X_08883_ _15324_/A _08883_/B vssd1 vssd1 vccd1 vccd1 _16059_/D sky130_fd_sc_hd__and2_1
Xhold2437 _18452_/Q vssd1 vssd1 vccd1 vccd1 hold2437/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1703 _09097_/X vssd1 vssd1 vccd1 vccd1 _16163_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2448 _09105_/X vssd1 vssd1 vccd1 vccd1 _16167_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1714 _18225_/Q vssd1 vssd1 vccd1 vccd1 hold1714/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2459 _16240_/Q vssd1 vssd1 vccd1 vccd1 hold2459/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1725 _14623_/X vssd1 vssd1 vccd1 vccd1 _18105_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07834_ hold1775/X _07865_/B _07833_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _07834_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_237_1331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1736 _17909_/Q vssd1 vssd1 vccd1 vccd1 hold1736/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1747 _14229_/X vssd1 vssd1 vccd1 vccd1 _17916_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1758 input62/X vssd1 vssd1 vccd1 vccd1 hold1758/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1769 _09411_/X vssd1 vssd1 vccd1 vccd1 _16291_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09504_ _09984_/A _09504_/B vssd1 vssd1 vccd1 vccd1 _09504_/X sky130_fd_sc_hd__or2_1
XFILLER_0_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09435_ _07785_/Y _09483_/B _09440_/B hold714/X vssd1 vssd1 vccd1 vccd1 hold715/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09366_ _09366_/A _09366_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09366_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_192_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08317_ _15541_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08317_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_40 _13260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ _15519_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09297_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_51 hold62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_62 hold384/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_73 hold597/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ _14413_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08248_/X sky130_fd_sc_hd__or2_1
XANTENNA_84 _15145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_409_wb_clk_i clkbuf_6_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17771_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_95 hold5967/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08179_ hold911/X _08225_/B vssd1 vssd1 vccd1 vccd1 _08179_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5030 _16356_/Q vssd1 vssd1 vccd1 vccd1 hold5030/X sky130_fd_sc_hd__dlygate4sd3_1
X_10210_ hold3913/X _10598_/B _10209_/X _15218_/C1 vssd1 vssd1 vccd1 vccd1 _10210_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5041 _11110_/X vssd1 vssd1 vccd1 vccd1 _16860_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5052 _16954_/Q vssd1 vssd1 vccd1 vccd1 hold5052/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11190_ hold4381/X _11121_/A _11189_/X vssd1 vssd1 vccd1 vccd1 _11190_/Y sky130_fd_sc_hd__a21oi_1
Xhold5063 _12025_/X vssd1 vssd1 vccd1 vccd1 _17165_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5074 _16864_/Q vssd1 vssd1 vccd1 vccd1 hold5074/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4340 hold6127/X vssd1 vssd1 vccd1 vccd1 hold4340/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold5085 _13510_/X vssd1 vssd1 vccd1 vccd1 _17623_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10141_ hold3779/X _10619_/B _10140_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10141_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5096 _11122_/X vssd1 vssd1 vccd1 vccd1 _16864_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4351 _11181_/Y vssd1 vssd1 vccd1 vccd1 _11182_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4362 _12303_/Y vssd1 vssd1 vccd1 vccd1 _12304_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4373 _17095_/Q vssd1 vssd1 vccd1 vccd1 hold4373/X sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_6546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4384 _16917_/Q vssd1 vssd1 vccd1 vccd1 hold4384/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3650 _16411_/Q vssd1 vssd1 vccd1 vccd1 hold3650/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4395 _11764_/Y vssd1 vssd1 vccd1 vccd1 _17078_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3661 _09772_/X vssd1 vssd1 vccd1 vccd1 _16414_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10072_ _11206_/A _10072_/B vssd1 vssd1 vccd1 vccd1 _16514_/D sky130_fd_sc_hd__nor2_1
XTAP_6579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3672 _16680_/Q vssd1 vssd1 vccd1 vccd1 hold3672/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3683 _09574_/X vssd1 vssd1 vccd1 vccd1 _16348_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3694 _16393_/Q vssd1 vssd1 vccd1 vccd1 hold3694/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_6_11_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_11_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_13900_ _15189_/A hold2890/X hold297/X vssd1 vssd1 vccd1 vccd1 _13901_/B sky130_fd_sc_hd__mux2_1
XTAP_5867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2960 _17819_/Q vssd1 vssd1 vccd1 vccd1 hold2960/X sky130_fd_sc_hd__dlygate4sd3_1
X_14880_ _15165_/A _14880_/B vssd1 vssd1 vccd1 vccd1 _14880_/Y sky130_fd_sc_hd__nand2_1
XTAP_5878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2971 _15778_/Q vssd1 vssd1 vccd1 vccd1 hold2971/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2982 _14522_/X vssd1 vssd1 vccd1 vccd1 _18057_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2993 _15564_/Q vssd1 vssd1 vccd1 vccd1 hold2993/X sky130_fd_sc_hd__dlygate4sd3_1
X_13831_ _13864_/A _13831_/B vssd1 vssd1 vccd1 vccd1 _13831_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_230_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16550_ _18164_/CLK _16550_/D vssd1 vssd1 vccd1 vccd1 _16550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13762_ hold5287/X _13856_/B _13761_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13762_/X
+ sky130_fd_sc_hd__o211a_1
X_10974_ _11655_/A _10974_/B vssd1 vssd1 vccd1 vccd1 _10974_/X sky130_fd_sc_hd__or2_1
XFILLER_0_58_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15501_ _15517_/A hold2217/X _15505_/S vssd1 vssd1 vccd1 vccd1 _15502_/B sky130_fd_sc_hd__mux2_1
X_12713_ hold3826/X _12712_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12713_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16481_ _18394_/CLK _16481_/D vssd1 vssd1 vccd1 vccd1 _16481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13693_ hold5482/X _13883_/B _13692_/X _08347_/A vssd1 vssd1 vccd1 vccd1 _13693_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18220_ _18220_/CLK _18220_/D vssd1 vssd1 vccd1 vccd1 _18220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15432_ _15480_/A _15432_/B _15432_/C _15432_/D vssd1 vssd1 vccd1 vccd1 _15432_/X
+ sky130_fd_sc_hd__or4_1
X_12644_ hold3359/X _12643_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12645_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18151_ _18197_/CLK _18151_/D vssd1 vssd1 vccd1 vccd1 _18151_/Q sky130_fd_sc_hd__dfxtp_1
X_15363_ _15490_/A1 _15355_/X _15362_/X _15490_/B1 hold5944/A vssd1 vssd1 vccd1 vccd1
+ _15363_/X sky130_fd_sc_hd__a32o_1
X_12575_ hold3235/X _12574_/X _12971_/S vssd1 vssd1 vccd1 vccd1 _12575_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17102_ _17262_/CLK _17102_/D vssd1 vssd1 vccd1 vccd1 _17102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14314_ _14529_/A _14334_/B vssd1 vssd1 vccd1 vccd1 _14314_/X sky130_fd_sc_hd__or2_1
X_18082_ _18129_/CLK _18082_/D vssd1 vssd1 vccd1 vccd1 _18082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11526_ _12210_/A _11526_/B vssd1 vssd1 vccd1 vccd1 _11526_/X sky130_fd_sc_hd__or2_1
X_15294_ _15414_/A _15294_/B vssd1 vssd1 vccd1 vccd1 _18405_/D sky130_fd_sc_hd__and2_1
XFILLER_0_145_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17033_ _17881_/CLK _17033_/D vssd1 vssd1 vccd1 vccd1 _17033_/Q sky130_fd_sc_hd__dfxtp_1
X_14245_ hold651/X _14268_/B _14244_/X _14352_/A vssd1 vssd1 vccd1 vccd1 hold652/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11457_ _11553_/A _11457_/B vssd1 vssd1 vccd1 vccd1 _11457_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10408_ hold5616/X _11213_/B _10407_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10408_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_6_50_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_50_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14176_ _14461_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14176_/X sky130_fd_sc_hd__or2_1
X_11388_ _11667_/A _11388_/B vssd1 vssd1 vccd1 vccd1 _11388_/X sky130_fd_sc_hd__or2_1
XFILLER_0_221_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ hold3280/X _10589_/B _10338_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _10339_/X
+ sky130_fd_sc_hd__o211a_1
X_13127_ _13199_/A1 _13125_/X _13126_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13127_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ _18031_/CLK _17935_/D vssd1 vssd1 vccd1 vccd1 _17935_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _17558_/Q _17092_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13058_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_237_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12009_ _13716_/A _12009_/B vssd1 vssd1 vccd1 vccd1 _12009_/X sky130_fd_sc_hd__or2_1
X_17866_ _17898_/CLK _17866_/D vssd1 vssd1 vccd1 vccd1 _17866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16817_ _18052_/CLK _16817_/D vssd1 vssd1 vccd1 vccd1 _16817_/Q sky130_fd_sc_hd__dfxtp_1
X_17797_ _17831_/CLK _17797_/D vssd1 vssd1 vccd1 vccd1 _17797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16748_ _17983_/CLK _16748_/D vssd1 vssd1 vccd1 vccd1 _16748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_1323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16679_ _18205_/CLK _16679_/D vssd1 vssd1 vccd1 vccd1 _16679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09220_ _15549_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09220_/X sky130_fd_sc_hd__or2_1
X_18418_ _18418_/CLK _18418_/D vssd1 vssd1 vccd1 vccd1 _18418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09151_ hold3037/X _09164_/B _09150_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _09151_/X
+ sky130_fd_sc_hd__o211a_1
X_18349_ _18349_/CLK _18349_/D vssd1 vssd1 vccd1 vccd1 _18349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08102_ hold405/A hold337/A hold509/A hold444/A vssd1 vssd1 vccd1 vccd1 hold306/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09082_ hold933/X _09118_/B vssd1 vssd1 vccd1 vccd1 _09082_/X sky130_fd_sc_hd__or2_1
XFILLER_0_71_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08033_ _15221_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _08033_/Y sky130_fd_sc_hd__nand2_1
Xhold800 hold800/A vssd1 vssd1 vccd1 vccd1 hold800/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput60 input60/A vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__buf_6
Xhold811 hold811/A vssd1 vssd1 vccd1 vccd1 hold811/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput71 wb_rst_i vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_1366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold822 hold822/A vssd1 vssd1 vccd1 vccd1 hold822/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 hold833/A vssd1 vssd1 vccd1 vccd1 hold833/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_12_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold844 hold844/A vssd1 vssd1 vccd1 vccd1 hold844/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 hold855/A vssd1 vssd1 vccd1 vccd1 hold855/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold866 hold866/A vssd1 vssd1 vccd1 vccd1 hold866/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold877 hold877/A vssd1 vssd1 vccd1 vccd1 hold877/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold888 hold888/A vssd1 vssd1 vccd1 vccd1 hold888/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 input1/X vssd1 vssd1 vccd1 vccd1 hold899/X sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ _09984_/A _09984_/B vssd1 vssd1 vccd1 vccd1 _09984_/X sky130_fd_sc_hd__or2_1
XFILLER_0_229_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2201 _18448_/Q vssd1 vssd1 vccd1 vccd1 hold2201/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2212 _15160_/X vssd1 vssd1 vccd1 vccd1 _18363_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08935_ hold226/X hold720/X _08991_/S vssd1 vssd1 vccd1 vccd1 hold721/A sky130_fd_sc_hd__mux2_1
Xhold2223 _18429_/Q vssd1 vssd1 vccd1 vccd1 hold2223/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2234 _15732_/Q vssd1 vssd1 vccd1 vccd1 hold2234/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2245 _14073_/X vssd1 vssd1 vccd1 vccd1 _17841_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1500 _09334_/X vssd1 vssd1 vccd1 vccd1 _16277_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1511 _17840_/Q vssd1 vssd1 vccd1 vccd1 hold1511/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2256 _17763_/Q vssd1 vssd1 vccd1 vccd1 hold2256/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1522 _09413_/X vssd1 vssd1 vccd1 vccd1 _16292_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2267 _12621_/X vssd1 vssd1 vccd1 vccd1 _17383_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08866_ hold278/X hold697/X _08866_/S vssd1 vssd1 vccd1 vccd1 hold698/A sky130_fd_sc_hd__mux2_1
Xhold1533 _08176_/X vssd1 vssd1 vccd1 vccd1 _15724_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2278 _12626_/X vssd1 vssd1 vccd1 vccd1 _12627_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1544 _15680_/Q vssd1 vssd1 vccd1 vccd1 hold1544/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2289 _16206_/Q vssd1 vssd1 vccd1 vccd1 hold2289/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1555 _07872_/X vssd1 vssd1 vccd1 vccd1 _15581_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07817_ _07817_/A _07817_/B _07817_/C _07817_/D vssd1 vssd1 vccd1 vccd1 _09366_/A
+ sky130_fd_sc_hd__or4_4
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1566 _15786_/Q vssd1 vssd1 vccd1 vccd1 hold1566/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08797_ hold226/X hold747/X _08801_/S vssd1 vssd1 vccd1 vccd1 hold748/A sky130_fd_sc_hd__mux2_1
Xhold1577 _14935_/X vssd1 vssd1 vccd1 vccd1 _18254_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1588 _17951_/Q vssd1 vssd1 vccd1 vccd1 hold1588/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1599 _14785_/X vssd1 vssd1 vccd1 vccd1 _18183_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09418_ _09438_/B _09418_/B vssd1 vssd1 vccd1 vccd1 _09418_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10690_ hold5450/X _11071_/A2 _10689_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _10690_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09349_ _09366_/A _09351_/B _09364_/B vssd1 vssd1 vccd1 vccd1 _09349_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_168_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12360_ hold5708/X _12267_/A _12359_/X vssd1 vssd1 vccd1 vccd1 _12360_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_243_wb_clk_i clkbuf_6_57_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18210_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11311_ hold4933/X _11789_/B _11310_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _11311_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12291_ _13797_/A _12291_/B vssd1 vssd1 vccd1 vccd1 _12291_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14030_ _15537_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14030_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11242_ hold5691/X _12299_/B _11241_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _11242_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11173_ _12301_/A _11173_/B vssd1 vssd1 vccd1 vccd1 _11173_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4170 _09748_/X vssd1 vssd1 vccd1 vccd1 _16406_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4181 hold5919/X vssd1 vssd1 vccd1 vccd1 hold5920/A sky130_fd_sc_hd__buf_4
X_10124_ hold2737/X _16532_/Q _10646_/C vssd1 vssd1 vccd1 vccd1 _10125_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4192 _15333_/X vssd1 vssd1 vccd1 vccd1 _15334_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15981_ _17300_/CLK _15981_/D vssd1 vssd1 vccd1 vccd1 hold634/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_234_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3480 _11157_/Y vssd1 vssd1 vccd1 vccd1 _11158_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17720_ _17720_/CLK _17720_/D vssd1 vssd1 vccd1 vccd1 _17720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10055_ _16509_/Q _10601_/B _10601_/C vssd1 vssd1 vccd1 vccd1 _10055_/X sky130_fd_sc_hd__and3_1
XTAP_5653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14932_ _15201_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14932_/X sky130_fd_sc_hd__or2_1
Xhold3491 _11184_/Y vssd1 vssd1 vccd1 vccd1 _11185_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2790 _15736_/Q vssd1 vssd1 vccd1 vccd1 hold2790/X sky130_fd_sc_hd__dlygate4sd3_1
X_17651_ _17747_/CLK _17651_/D vssd1 vssd1 vccd1 vccd1 _17651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ hold2735/X hold332/X _14862_/X _14863_/C1 vssd1 vssd1 vccd1 vccd1 _14863_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16602_ _18224_/CLK _16602_/D vssd1 vssd1 vccd1 vccd1 _16602_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13814_ _17725_/Q _13814_/B _13814_/C vssd1 vssd1 vccd1 vccd1 _13814_/X sky130_fd_sc_hd__and3_1
X_17582_ _17584_/CLK _17582_/D vssd1 vssd1 vccd1 vccd1 _17582_/Q sky130_fd_sc_hd__dfxtp_1
X_14794_ _15187_/A _14830_/B vssd1 vssd1 vccd1 vccd1 _14794_/X sky130_fd_sc_hd__or2_1
XFILLER_0_159_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16533_ _18099_/CLK _16533_/D vssd1 vssd1 vccd1 vccd1 _16533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13745_ hold1099/X _17702_/Q _13841_/C vssd1 vssd1 vccd1 vccd1 _13746_/B sky130_fd_sc_hd__mux2_1
X_10957_ hold5088/X _11153_/B _10956_/X _14354_/A vssd1 vssd1 vccd1 vccd1 _10957_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16464_ _18377_/CLK _16464_/D vssd1 vssd1 vccd1 vccd1 _16464_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13676_ hold2762/X hold3989/X _13865_/C vssd1 vssd1 vccd1 vccd1 _13677_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10888_ hold5165/X _11210_/B _10887_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _10888_/X
+ sky130_fd_sc_hd__o211a_1
X_18203_ _18203_/CLK _18203_/D vssd1 vssd1 vccd1 vccd1 _18203_/Q sky130_fd_sc_hd__dfxtp_1
X_15415_ hold458/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15415_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12627_ _12864_/A _12627_/B vssd1 vssd1 vccd1 vccd1 _17385_/D sky130_fd_sc_hd__and2_1
XPHY_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16395_ _18308_/CLK _16395_/D vssd1 vssd1 vccd1 vccd1 _16395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18134_ _18166_/CLK _18134_/D vssd1 vssd1 vccd1 vccd1 _18134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15346_ _17338_/Q _09362_/C _09362_/D hold570/X vssd1 vssd1 vccd1 vccd1 _15346_/X
+ sky130_fd_sc_hd__a22o_1
X_12558_ _12906_/A _12558_/B vssd1 vssd1 vccd1 vccd1 _17362_/D sky130_fd_sc_hd__and2_1
X_11509_ hold4941/X _11798_/B _11508_/X _14143_/C1 vssd1 vssd1 vccd1 vccd1 _11509_/X
+ sky130_fd_sc_hd__o211a_1
X_18065_ _18065_/CLK _18065_/D vssd1 vssd1 vccd1 vccd1 _18065_/Q sky130_fd_sc_hd__dfxtp_1
X_15277_ hold301/X _15487_/A2 _15484_/B1 hold118/X _15276_/X vssd1 vssd1 vccd1 vccd1
+ _15282_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_151_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12489_ hold47/X _12509_/A2 _12501_/A3 _12488_/X _15344_/A vssd1 vssd1 vccd1 vccd1
+ hold48/A sky130_fd_sc_hd__o311a_1
XFILLER_0_123_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold107 hold107/A vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__buf_1
Xhold118 hold118/A vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold129 hold37/X vssd1 vssd1 vccd1 vccd1 input27/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17016_ _17936_/CLK _17016_/D vssd1 vssd1 vccd1 vccd1 _17016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14228_ _15519_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14228_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_223_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14159_ hold1560/X _14148_/B _14158_/X _13895_/A vssd1 vssd1 vccd1 vccd1 _14159_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout609 _09363_/Y vssd1 vssd1 vccd1 vccd1 _15488_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_226_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08720_ _08851_/A hold635/X vssd1 vssd1 vccd1 vccd1 _15981_/D sky130_fd_sc_hd__and2_1
X_17918_ _18016_/CLK _17918_/D vssd1 vssd1 vccd1 vccd1 _17918_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_47_wb_clk_i clkbuf_6_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17913_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_217_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08651_ hold315/X hold867/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08652_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_234_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17849_ _17850_/CLK _17849_/D vssd1 vssd1 vccd1 vccd1 _17849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08582_ hold438/X hold470/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08583_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09203_ hold1248/X _09214_/B _09202_/X _12804_/A vssd1 vssd1 vccd1 vccd1 _09203_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09134_ _15517_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09134_/X sky130_fd_sc_hd__or2_1
XFILLER_0_72_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09065_ _14555_/C hold268/X vssd1 vssd1 vccd1 vccd1 hold362/A sky130_fd_sc_hd__or2_1
XFILLER_0_163_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08016_ hold2373/X _08029_/B _08015_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _08016_/X
+ sky130_fd_sc_hd__o211a_1
Xhold630 hold630/A vssd1 vssd1 vccd1 vccd1 hold630/X sky130_fd_sc_hd__buf_8
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold641 hold641/A vssd1 vssd1 vccd1 vccd1 hold641/X sky130_fd_sc_hd__buf_4
XFILLER_0_124_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold652 hold652/A vssd1 vssd1 vccd1 vccd1 hold652/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold663 hold663/A vssd1 vssd1 vccd1 vccd1 hold663/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 hold674/A vssd1 vssd1 vccd1 vccd1 hold674/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold685 hold685/A vssd1 vssd1 vccd1 vccd1 hold685/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold696 hold696/A vssd1 vssd1 vccd1 vccd1 hold696/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09967_ hold3541/X _10577_/B _09966_/X _15204_/C1 vssd1 vssd1 vccd1 vccd1 _09967_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2020 _14659_/X vssd1 vssd1 vccd1 vccd1 _18122_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2031 _16172_/Q vssd1 vssd1 vccd1 vccd1 hold2031/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2042 _08506_/X vssd1 vssd1 vccd1 vccd1 _15880_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08918_ hold143/X hold675/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08919_/B sky130_fd_sc_hd__mux2_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2053 _17897_/Q vssd1 vssd1 vccd1 vccd1 hold2053/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2064 _18187_/Q vssd1 vssd1 vccd1 vccd1 hold2064/X sky130_fd_sc_hd__dlygate4sd3_1
X_09898_ hold4773/X _09992_/B _09897_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _09898_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2075 _18269_/Q vssd1 vssd1 vccd1 vccd1 hold2075/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1330 _15846_/Q vssd1 vssd1 vccd1 vccd1 hold1330/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2086 _18063_/Q vssd1 vssd1 vccd1 vccd1 hold2086/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1341 _08491_/X vssd1 vssd1 vccd1 vccd1 _15874_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2097 _14833_/X vssd1 vssd1 vccd1 vccd1 _18206_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1352 _15662_/Q vssd1 vssd1 vccd1 vccd1 hold1352/X sky130_fd_sc_hd__dlygate4sd3_1
X_08849_ _12412_/A _08849_/B vssd1 vssd1 vccd1 vccd1 _16043_/D sky130_fd_sc_hd__and2_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1363 _14193_/X vssd1 vssd1 vccd1 vccd1 _17899_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1374 _18359_/Q vssd1 vssd1 vccd1 vccd1 hold1374/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1385 _09405_/X vssd1 vssd1 vccd1 vccd1 _16288_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1396 _08453_/X vssd1 vssd1 vccd1 vccd1 _15855_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ hold5769/X _12350_/B _11859_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _11860_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10811_ hold1662/X hold4135/X _11660_/S vssd1 vssd1 vccd1 vccd1 _10812_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_138_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ _12337_/A _11791_/B vssd1 vssd1 vccd1 vccd1 _11791_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_1253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13530_ _13734_/A _13530_/B vssd1 vssd1 vccd1 vccd1 _13530_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10742_ hold2777/X _16738_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _10743_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_424_wb_clk_i clkbuf_6_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17261_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10673_ hold2165/X hold4259/X _11153_/C vssd1 vssd1 vccd1 vccd1 _10674_/B sky130_fd_sc_hd__mux2_1
X_13461_ _13599_/A _13461_/B vssd1 vssd1 vccd1 vccd1 _13461_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15200_ hold3108/X _15219_/B _15199_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _15200_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12412_ _12412_/A hold771/X vssd1 vssd1 vccd1 vccd1 _17299_/D sky130_fd_sc_hd__and2_1
XFILLER_0_180_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16180_ _17464_/CLK _16180_/D vssd1 vssd1 vccd1 vccd1 _16180_/Q sky130_fd_sc_hd__dfxtp_1
X_13392_ _13773_/A _13392_/B vssd1 vssd1 vccd1 vccd1 _13392_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15131_ _15185_/A _15157_/B vssd1 vssd1 vccd1 vccd1 _15131_/X sky130_fd_sc_hd__or2_1
X_12343_ _13888_/A _12343_/B vssd1 vssd1 vccd1 vccd1 _12343_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_181_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15062_ _15062_/A _15062_/B vssd1 vssd1 vccd1 vccd1 _18316_/D sky130_fd_sc_hd__and2_1
XFILLER_0_209_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12274_ hold4921/X _13886_/B _12273_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _12274_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11225_ _16899_/Q _11225_/B _11765_/C vssd1 vssd1 vccd1 vccd1 _11225_/X sky130_fd_sc_hd__and3_1
X_14013_ hold1167/X _14038_/B _14012_/X _14211_/C1 vssd1 vssd1 vccd1 vccd1 _14013_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11156_ _16876_/Q _11201_/B _11201_/C vssd1 vssd1 vccd1 vccd1 _11156_/X sky130_fd_sc_hd__and3_1
XTAP_6140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10107_ _10515_/A _10107_/B vssd1 vssd1 vccd1 vccd1 _10107_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15964_ _17318_/CLK _15964_/D vssd1 vssd1 vccd1 vccd1 hold513/A sky130_fd_sc_hd__dfxtp_1
XTAP_5450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11087_ hold3093/X _16853_/Q _11183_/C vssd1 vssd1 vccd1 vccd1 _11088_/B sky130_fd_sc_hd__mux2_1
XTAP_6195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17703_ _17703_/CLK _17703_/D vssd1 vssd1 vccd1 vccd1 _17703_/Q sky130_fd_sc_hd__dfxtp_1
X_10038_ _13214_/A _10386_/A _10037_/X vssd1 vssd1 vccd1 vccd1 _10038_/Y sky130_fd_sc_hd__a21oi_1
X_14915_ hold1835/X _14946_/B _14914_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _14915_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15895_ _17347_/CLK _15895_/D vssd1 vssd1 vccd1 vccd1 hold659/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17634_ _17730_/CLK _17634_/D vssd1 vssd1 vccd1 vccd1 _17634_/Q sky130_fd_sc_hd__dfxtp_1
X_14846_ _15185_/A _14892_/B vssd1 vssd1 vccd1 vccd1 _14846_/X sky130_fd_sc_hd__or2_1
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17565_ _17624_/CLK _17565_/D vssd1 vssd1 vccd1 vccd1 _17565_/Q sky130_fd_sc_hd__dfxtp_1
X_14777_ hold1781/X _14774_/B _14776_/X _14853_/C1 vssd1 vssd1 vccd1 vccd1 _14777_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_1387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11989_ hold5305/X _12365_/B _11988_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _11989_/X
+ sky130_fd_sc_hd__o211a_1
X_16516_ _18106_/CLK _16516_/D vssd1 vssd1 vccd1 vccd1 _16516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13728_ _13794_/A _13728_/B vssd1 vssd1 vccd1 vccd1 _13728_/X sky130_fd_sc_hd__or2_1
X_17496_ _17500_/CLK _17496_/D vssd1 vssd1 vccd1 vccd1 _17496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_165_wb_clk_i clkbuf_6_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18399_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_190_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16447_ _18392_/CLK _16447_/D vssd1 vssd1 vccd1 vccd1 _16447_/Q sky130_fd_sc_hd__dfxtp_1
X_13659_ _13791_/A _13659_/B vssd1 vssd1 vccd1 vccd1 _13659_/X sky130_fd_sc_hd__or2_1
XFILLER_0_229_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16378_ _18361_/CLK _16378_/D vssd1 vssd1 vccd1 vccd1 _16378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18117_ _18225_/CLK _18117_/D vssd1 vssd1 vccd1 vccd1 _18117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15329_ hold471/X _15485_/A2 _15488_/A2 hold661/X _15328_/X vssd1 vssd1 vccd1 vccd1
+ _15332_/C sky130_fd_sc_hd__a221o_1
Xhold5607 _17205_/Q vssd1 vssd1 vccd1 vccd1 hold5607/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5618 _16826_/Q vssd1 vssd1 vccd1 vccd1 hold5618/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5629 _13558_/X vssd1 vssd1 vccd1 vccd1 _17639_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18048_ _18048_/CLK _18048_/D vssd1 vssd1 vccd1 vccd1 _18048_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4906 _10678_/X vssd1 vssd1 vccd1 vccd1 _16716_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4917 _17183_/Q vssd1 vssd1 vccd1 vccd1 hold4917/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4928 _11971_/X vssd1 vssd1 vccd1 vccd1 _17147_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4939 _17079_/Q vssd1 vssd1 vccd1 vccd1 hold4939/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout406 _14334_/B vssd1 vssd1 vccd1 vccd1 _14338_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_226_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09821_ hold2709/X hold4557/X _10028_/C vssd1 vssd1 vccd1 vccd1 _09822_/B sky130_fd_sc_hd__mux2_1
Xfanout417 _14108_/Y vssd1 vssd1 vccd1 vccd1 _14142_/B sky130_fd_sc_hd__buf_6
XFILLER_0_238_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout428 hold296/X vssd1 vssd1 vccd1 vccd1 _13942_/S sky130_fd_sc_hd__clkbuf_8
Xfanout439 _13721_/S vssd1 vssd1 vccd1 vccd1 _13796_/S sky130_fd_sc_hd__buf_6
XFILLER_0_158_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09752_ hold1388/X _16408_/Q _10985_/S vssd1 vssd1 vccd1 vccd1 _09753_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_225_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_236_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08703_ hold215/X hold638/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08704_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_146_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09683_ hold1917/X hold3270/X _10571_/C vssd1 vssd1 vccd1 vccd1 _09684_/B sky130_fd_sc_hd__mux2_1
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _15414_/A _08634_/B vssd1 vssd1 vccd1 vccd1 _15939_/D sky130_fd_sc_hd__and2_1
XFILLER_0_59_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _15491_/A hold746/X vssd1 vssd1 vccd1 vccd1 _15906_/D sky130_fd_sc_hd__and2_1
XFILLER_0_194_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08496_ _14960_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08496_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09117_ hold2060/X _09106_/B _09116_/X _15244_/A vssd1 vssd1 vccd1 vccd1 _09117_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09048_ hold143/X _16141_/Q _09056_/S vssd1 vssd1 vccd1 vccd1 hold144/A sky130_fd_sc_hd__mux2_1
XFILLER_0_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold460 hold460/A vssd1 vssd1 vccd1 vccd1 hold460/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold471 hold471/A vssd1 vssd1 vccd1 vccd1 hold471/X sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ _11010_/A _11010_/B vssd1 vssd1 vccd1 vccd1 _11010_/X sky130_fd_sc_hd__or2_1
Xhold482 hold482/A vssd1 vssd1 vccd1 vccd1 input49/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 hold55/X vssd1 vssd1 vccd1 vccd1 input26/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout940 hold1007/X vssd1 vssd1 vccd1 vccd1 _14596_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12961_ hold2719/X hold3212/X _12970_/S vssd1 vssd1 vccd1 vccd1 _12961_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_232_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1160 _14339_/X vssd1 vssd1 vccd1 vccd1 _17969_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14700_ _15201_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14700_/X sky130_fd_sc_hd__or2_1
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1171 _07955_/X vssd1 vssd1 vccd1 vccd1 _15620_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1182 input41/X vssd1 vssd1 vccd1 vccd1 hold691/A sky130_fd_sc_hd__buf_1
X_11912_ hold2877/X _17128_/Q _13811_/C vssd1 vssd1 vccd1 vccd1 _11913_/B sky130_fd_sc_hd__mux2_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _17270_/CLK _15680_/D vssd1 vssd1 vccd1 vccd1 _15680_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 hold926/X vssd1 vssd1 vccd1 vccd1 hold1193/X sky130_fd_sc_hd__clkbuf_16
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ hold2181/X _17475_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12892_/X sky130_fd_sc_hd__mux2_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ hold1652/X _14666_/B _14630_/X _14895_/C1 vssd1 vssd1 vccd1 vccd1 _14631_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11843_ hold2787/X hold4438/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11844_/B sky130_fd_sc_hd__mux2_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17350_ _17512_/CLK _17350_/D vssd1 vssd1 vccd1 vccd1 _17350_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _15492_/A _14573_/B _18076_/Q vssd1 vssd1 vccd1 vccd1 _14562_/X sky130_fd_sc_hd__a21o_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _17082_/Q _11798_/B _11774_/C vssd1 vssd1 vccd1 vccd1 _11774_/X sky130_fd_sc_hd__and3_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _16323_/CLK _16301_/D vssd1 vssd1 vccd1 vccd1 _16301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13513_ hold5207/X _13817_/B _13512_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _13513_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10725_ _11109_/A _10725_/B vssd1 vssd1 vccd1 vccd1 _10725_/X sky130_fd_sc_hd__or2_1
X_17281_ _17281_/CLK _17281_/D vssd1 vssd1 vccd1 vccd1 _17281_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14493_ _15173_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14493_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16232_ _17754_/CLK _16232_/D vssd1 vssd1 vccd1 vccd1 _16232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13444_ hold4642/X _13862_/B _13443_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13444_/X
+ sky130_fd_sc_hd__o211a_1
X_10656_ _11136_/A _10656_/B vssd1 vssd1 vccd1 vccd1 _10656_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16163_ _17499_/CLK _16163_/D vssd1 vssd1 vccd1 vccd1 _16163_/Q sky130_fd_sc_hd__dfxtp_1
X_10587_ hold3486/X _10530_/A _10586_/X vssd1 vssd1 vccd1 vccd1 _10587_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13375_ hold5341/X _13874_/B _13374_/X _13684_/C1 vssd1 vssd1 vccd1 vccd1 _13375_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15114_ hold2605/X hold340/X _15113_/Y _15054_/A vssd1 vssd1 vccd1 vccd1 _15114_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12326_ _17266_/Q _12356_/B _13481_/S vssd1 vssd1 vccd1 vccd1 _12326_/X sky130_fd_sc_hd__and3_1
XFILLER_0_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16094_ _18418_/CLK _16094_/D vssd1 vssd1 vccd1 vccd1 _16094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15045_ _15099_/A hold2579/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15046_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12257_ hold1740/X _17243_/Q _13409_/S vssd1 vssd1 vccd1 vccd1 _12258_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11208_ hold4399/X _11127_/A _11207_/X vssd1 vssd1 vccd1 vccd1 _11208_/Y sky130_fd_sc_hd__a21oi_1
X_12188_ hold2599/X _17220_/Q _12305_/C vssd1 vssd1 vccd1 vccd1 _12189_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_236_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_236_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11139_ _11637_/A _11139_/B vssd1 vssd1 vccd1 vccd1 _11139_/X sky130_fd_sc_hd__or2_1
XFILLER_0_207_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16996_ _17856_/CLK _16996_/D vssd1 vssd1 vccd1 vccd1 _16996_/Q sky130_fd_sc_hd__dfxtp_1
X_15947_ _17337_/CLK _15947_/D vssd1 vssd1 vccd1 vccd1 hold528/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15878_ _17735_/CLK _15878_/D vssd1 vssd1 vccd1 vccd1 _15878_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_346_wb_clk_i clkbuf_6_42_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17737_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_188_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_231_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14829_ hold1064/X _14828_/B _14828_/Y _14895_/C1 vssd1 vssd1 vccd1 vccd1 _14829_/X
+ sky130_fd_sc_hd__o211a_1
X_17617_ _17617_/CLK _17617_/D vssd1 vssd1 vccd1 vccd1 _17617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08350_ _15085_/A hold963/X hold115/X vssd1 vssd1 vccd1 vccd1 hold964/A sky130_fd_sc_hd__mux2_1
X_17548_ _18217_/CLK _17548_/D vssd1 vssd1 vccd1 vccd1 _17548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08281_ hold1471/X _08268_/B _08280_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _08281_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17479_ _17481_/CLK _17479_/D vssd1 vssd1 vccd1 vccd1 _17479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6105 _17524_/Q vssd1 vssd1 vccd1 vccd1 hold6105/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6116 _16542_/Q vssd1 vssd1 vccd1 vccd1 hold6116/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6127 _16530_/Q vssd1 vssd1 vccd1 vccd1 hold6127/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5404 _17024_/Q vssd1 vssd1 vccd1 vccd1 hold5404/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5415 _13759_/X vssd1 vssd1 vccd1 vccd1 _17706_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5426 _16992_/Q vssd1 vssd1 vccd1 vccd1 hold5426/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5437 _11686_/X vssd1 vssd1 vccd1 vccd1 _17052_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4703 _17632_/Q vssd1 vssd1 vccd1 vccd1 hold4703/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5448 _16799_/Q vssd1 vssd1 vccd1 vccd1 hold5448/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4714 _09700_/X vssd1 vssd1 vccd1 vccd1 _16390_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5459 _12220_/X vssd1 vssd1 vccd1 vccd1 _17230_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4725 _16456_/Q vssd1 vssd1 vccd1 vccd1 hold4725/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4736 _09910_/X vssd1 vssd1 vccd1 vccd1 _16460_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_62_wb_clk_i clkbuf_6_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18461_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4747 _17508_/Q vssd1 vssd1 vccd1 vccd1 hold4747/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4758 _17631_/Q vssd1 vssd1 vccd1 vccd1 hold4758/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4769 _09814_/X vssd1 vssd1 vccd1 vccd1 _16428_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout203 fanout210/X vssd1 vssd1 vccd1 vccd1 _11210_/B sky130_fd_sc_hd__buf_4
Xfanout214 _11201_/B vssd1 vssd1 vccd1 vccd1 _11171_/B sky130_fd_sc_hd__clkbuf_8
Xfanout225 _10634_/B vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__buf_4
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout236 _10067_/B vssd1 vssd1 vccd1 vccd1 _10571_/B sky130_fd_sc_hd__buf_2
Xfanout247 _09494_/X vssd1 vssd1 vccd1 vccd1 _10634_/B sky130_fd_sc_hd__clkbuf_8
X_09804_ _11061_/A _09804_/B vssd1 vssd1 vccd1 vccd1 _09804_/X sky130_fd_sc_hd__or2_1
Xfanout258 _12216_/A vssd1 vssd1 vccd1 vccd1 _13482_/A sky130_fd_sc_hd__buf_4
XFILLER_0_227_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout269 _11655_/A vssd1 vssd1 vccd1 vccd1 _11649_/A sky130_fd_sc_hd__buf_4
XFILLER_0_5_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07996_ hold1600/X _08029_/B _07995_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _07996_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_1337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09735_ _11010_/A _09735_/B vssd1 vssd1 vccd1 vccd1 _09735_/X sky130_fd_sc_hd__or2_1
XFILLER_0_236_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09666_ _09978_/A _09666_/B vssd1 vssd1 vccd1 vccd1 _09666_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08617_ hold673/X hold859/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold860/A sky130_fd_sc_hd__mux2_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09987_/A _09597_/B vssd1 vssd1 vccd1 vccd1 _09597_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ hold452/X hold454/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08549_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_194_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08479_ hold1760/X _08486_/B _08478_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08479_/X
+ sky130_fd_sc_hd__o211a_1
X_10510_ _10604_/A _10646_/B _10509_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _16660_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11490_ _12285_/A _11490_/B vssd1 vssd1 vccd1 vccd1 _11490_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10441_ hold3830/X _10631_/B _10440_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10441_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13160_ _13153_/X _13159_/X _13296_/B1 vssd1 vssd1 vccd1 vccd1 _17538_/D sky130_fd_sc_hd__o21a_1
X_10372_ hold3720/X _10625_/B _10371_/X _14769_/C1 vssd1 vssd1 vccd1 vccd1 _10372_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12111_ _12198_/A _12111_/B vssd1 vssd1 vccd1 vccd1 _12111_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13091_ _13090_/X _16904_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13091_/X sky130_fd_sc_hd__mux2_1
Xhold5960 hold6093/X vssd1 vssd1 vccd1 vccd1 hold5960/X sky130_fd_sc_hd__buf_2
Xhold5971 _07826_/X vssd1 vssd1 vccd1 vccd1 hold5971/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold5982 _18461_/Q vssd1 vssd1 vccd1 vccd1 _07784_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5993 _16313_/Q vssd1 vssd1 vccd1 vccd1 hold5993/X sky130_fd_sc_hd__dlygate4sd3_1
X_12042_ _12234_/A _12042_/B vssd1 vssd1 vccd1 vccd1 _12042_/X sky130_fd_sc_hd__or2_1
Xhold290 hold290/A vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_217_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16850_ _18021_/CLK _16850_/D vssd1 vssd1 vccd1 vccd1 _16850_/Q sky130_fd_sc_hd__dfxtp_1
X_15801_ _17732_/CLK _15801_/D vssd1 vssd1 vccd1 vccd1 _15801_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout770 _08131_/A vssd1 vssd1 vccd1 vccd1 _08151_/A sky130_fd_sc_hd__buf_4
Xfanout781 _14526_/C1 vssd1 vssd1 vccd1 vccd1 _14392_/A sky130_fd_sc_hd__buf_4
Xfanout792 _15056_/A vssd1 vssd1 vccd1 vccd1 _15060_/A sky130_fd_sc_hd__buf_4
X_16781_ _18016_/CLK _16781_/D vssd1 vssd1 vccd1 vccd1 _16781_/Q sky130_fd_sc_hd__dfxtp_1
X_13993_ hold2639/X _13995_/A2 _13992_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _13993_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15732_ _17187_/CLK _15732_/D vssd1 vssd1 vccd1 vccd1 _15732_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12944_ hold4554/X _12943_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12945_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_172_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _18451_/CLK _18451_/D vssd1 vssd1 vccd1 vccd1 _18451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15663_ _17281_/CLK _15663_/D vssd1 vssd1 vccd1 vccd1 _15663_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ hold3306/X _12874_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12875_/X sky130_fd_sc_hd__mux2_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17402_ _18453_/CLK _17402_/D vssd1 vssd1 vccd1 vccd1 _17402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _15169_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14614_/X sky130_fd_sc_hd__or2_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _18382_/CLK _18382_/D vssd1 vssd1 vccd1 vccd1 _18382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11826_ _12093_/A _11826_/B vssd1 vssd1 vccd1 vccd1 _11826_/X sky130_fd_sc_hd__or2_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _17242_/CLK _15594_/D vssd1 vssd1 vccd1 vccd1 _15594_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _17339_/CLK hold51/X vssd1 vssd1 vccd1 vccd1 _17333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14545_ _15225_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14545_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ hold4549/X _12243_/A _11756_/X vssd1 vssd1 vccd1 vccd1 _11757_/Y sky130_fd_sc_hd__a21oi_1
X_10708_ hold4909/X _11186_/B _10707_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _10708_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17264_ _17264_/CLK _17264_/D vssd1 vssd1 vccd1 vccd1 _17264_/Q sky130_fd_sc_hd__dfxtp_1
X_14476_ hold1901/X _14481_/B _14475_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _14476_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11688_ _12234_/A _11688_/B vssd1 vssd1 vccd1 vccd1 _11688_/X sky130_fd_sc_hd__or2_1
XFILLER_0_154_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16215_ _17723_/CLK _16215_/D vssd1 vssd1 vccd1 vccd1 _16215_/Q sky130_fd_sc_hd__dfxtp_1
X_13427_ hold1125/X hold4697/X _13811_/C vssd1 vssd1 vccd1 vccd1 _13428_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_102_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10639_ _10651_/A _10639_/B vssd1 vssd1 vccd1 vccd1 _16703_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17195_ _18430_/CLK _17195_/D vssd1 vssd1 vccd1 vccd1 _17195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16146_ _17341_/CLK _16146_/D vssd1 vssd1 vccd1 vccd1 hold545/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ hold2246/X hold4402/X _13865_/C vssd1 vssd1 vccd1 vccd1 _13359_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_11_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12309_ hold3470/X _13797_/A _12308_/X vssd1 vssd1 vccd1 vccd1 _12309_/Y sky130_fd_sc_hd__a21oi_1
X_16077_ _18401_/CLK _16077_/D vssd1 vssd1 vccd1 vccd1 hold675/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13289_ _13289_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13289_/X sky130_fd_sc_hd__and2_1
XFILLER_0_122_1415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3309 _10327_/X vssd1 vssd1 vccd1 vccd1 _16599_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15028_ _15028_/A _15028_/B vssd1 vssd1 vccd1 vccd1 _18299_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2608 _14127_/X vssd1 vssd1 vccd1 vccd1 _17867_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2619 _07977_/X vssd1 vssd1 vccd1 vccd1 _15631_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07850_ hold2410/X _07869_/B _07849_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _07850_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1907 _18265_/Q vssd1 vssd1 vccd1 vccd1 hold1907/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1918 _15025_/X vssd1 vssd1 vccd1 vccd1 _15026_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1929 _16223_/Q vssd1 vssd1 vccd1 vccd1 hold1929/X sky130_fd_sc_hd__dlygate4sd3_1
X_07781_ hold220/X vssd1 vssd1 vccd1 vccd1 _07781_/Y sky130_fd_sc_hd__inv_2
Xinput3 input3/A vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
X_16979_ _18065_/CLK _16979_/D vssd1 vssd1 vccd1 vccd1 _16979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09520_ hold4777/X _11201_/B _09519_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _09520_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_180_wb_clk_i clkbuf_6_51_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18327_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_91_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09451_ _09456_/C _09456_/D _09450_/Y vssd1 vssd1 vccd1 vccd1 _16310_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_149_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08402_ hold2979/X _08442_/A2 _08401_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _08402_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09382_ _16103_/Q _09392_/B _09362_/D hold644/X _09381_/X vssd1 vssd1 vccd1 vccd1
+ _09383_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_59_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08333_ _15557_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08333_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08264_ _15543_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08264_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08195_ _15529_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08195_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5201 _16827_/Q vssd1 vssd1 vccd1 vccd1 hold5201/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5212 _13483_/X vssd1 vssd1 vccd1 vccd1 _17614_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5223 _17238_/Q vssd1 vssd1 vccd1 vccd1 hold5223/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5234 _13657_/X vssd1 vssd1 vccd1 vccd1 _17672_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5245 _16884_/Q vssd1 vssd1 vccd1 vccd1 hold5245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4500 _13843_/Y vssd1 vssd1 vccd1 vccd1 _17734_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4511 _17350_/Q vssd1 vssd1 vccd1 vccd1 hold4511/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5256 _12187_/X vssd1 vssd1 vccd1 vccd1 _17219_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4522 _10126_/X vssd1 vssd1 vccd1 vccd1 _16532_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5267 _16789_/Q vssd1 vssd1 vccd1 vccd1 hold5267/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5278 _09598_/X vssd1 vssd1 vccd1 vccd1 _16356_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4533 _11194_/Y vssd1 vssd1 vccd1 vccd1 _16888_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4544 _10168_/X vssd1 vssd1 vccd1 vccd1 _16546_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5289 _17701_/Q vssd1 vssd1 vccd1 vccd1 hold5289/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3810 _16691_/Q vssd1 vssd1 vccd1 vccd1 hold3810/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4555 _16598_/Q vssd1 vssd1 vccd1 vccd1 hold4555/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4566 _11830_/X vssd1 vssd1 vccd1 vccd1 _17100_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3821 _10837_/X vssd1 vssd1 vccd1 vccd1 _16769_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3832 _16689_/Q vssd1 vssd1 vccd1 vccd1 hold3832/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4577 _16640_/Q vssd1 vssd1 vccd1 vccd1 hold4577/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3843 _10759_/X vssd1 vssd1 vccd1 vccd1 _16743_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4588 _12022_/X vssd1 vssd1 vccd1 vccd1 _17164_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4599 _12989_/X vssd1 vssd1 vccd1 vccd1 _12990_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3854 _17136_/Q vssd1 vssd1 vccd1 vccd1 hold3854/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3865 _09685_/X vssd1 vssd1 vccd1 vccd1 _16385_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3876 _16582_/Q vssd1 vssd1 vccd1 vccd1 hold3876/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3887 _09970_/X vssd1 vssd1 vccd1 vccd1 _16480_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_268_wb_clk_i clkbuf_6_56_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18226_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_226_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3898 _10378_/X vssd1 vssd1 vccd1 vccd1 _16616_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07979_ hold2476/X _07978_/B _07978_/Y _08167_/A vssd1 vssd1 vccd1 vccd1 _07979_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_236_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09718_ hold4509/X _10028_/B _09717_/X _15048_/A vssd1 vssd1 vccd1 vccd1 _09718_/X
+ sky130_fd_sc_hd__o211a_1
X_10990_ hold4925/X _11186_/B _10989_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10990_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09649_ hold4034/X _10031_/B _09648_/X _15146_/C1 vssd1 vssd1 vccd1 vccd1 _09649_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12660_/A _12660_/B vssd1 vssd1 vccd1 vccd1 _17396_/D sky130_fd_sc_hd__and2_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11611_ hold4093/X _12335_/B _11610_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _11611_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12591_ _12597_/A _12591_/B vssd1 vssd1 vccd1 vccd1 _17373_/D sky130_fd_sc_hd__and2_1
XFILLER_0_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14330_ _14330_/A _14334_/B vssd1 vssd1 vccd1 vccd1 _14330_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11542_ hold5444/X _11732_/B _11541_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _11542_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14261_ hold2094/X _14268_/B _14260_/X _14342_/A vssd1 vssd1 vccd1 vccd1 _14261_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11473_ hold4989/X _11765_/B _11472_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _11473_/X
+ sky130_fd_sc_hd__o211a_1
X_16000_ _17291_/CLK _16000_/D vssd1 vssd1 vccd1 vccd1 hold877/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13212_ hold4381/X _13211_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13212_/X sky130_fd_sc_hd__mux2_2
X_10424_ hold2664/X hold4054/X _11213_/C vssd1 vssd1 vccd1 vccd1 _10425_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14192_ _15537_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14192_/X sky130_fd_sc_hd__or2_1
Xclkbuf_6_40_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_40_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13143_ _13199_/A1 _13141_/X _13142_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13143_/X
+ sky130_fd_sc_hd__o211a_1
X_10355_ hold2236/X hold4573/X _10646_/C vssd1 vssd1 vccd1 vccd1 _10356_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5790 _12076_/X vssd1 vssd1 vccd1 vccd1 _17182_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10286_ hold2035/X hold4013/X _11186_/C vssd1 vssd1 vccd1 vccd1 _10287_/B sky130_fd_sc_hd__mux2_1
X_17951_ _17983_/CLK _17951_/D vssd1 vssd1 vccd1 vccd1 _17951_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _17560_/Q _17094_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13074_/X sky130_fd_sc_hd__mux2_1
X_12025_ hold5062/X _12217_/A2 _12024_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _12025_/X
+ sky130_fd_sc_hd__o211a_1
X_16902_ _18427_/CLK _16902_/D vssd1 vssd1 vccd1 vccd1 _16902_/Q sky130_fd_sc_hd__dfxtp_1
X_17882_ _17882_/CLK hold885/X vssd1 vssd1 vccd1 vccd1 hold884/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16833_ _18070_/CLK _16833_/D vssd1 vssd1 vccd1 vccd1 _16833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16764_ _17967_/CLK _16764_/D vssd1 vssd1 vccd1 vccd1 _16764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13976_ _14477_/A _13994_/B vssd1 vssd1 vccd1 vccd1 _13976_/X sky130_fd_sc_hd__or2_1
XFILLER_0_232_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15715_ _17735_/CLK _15715_/D vssd1 vssd1 vccd1 vccd1 _15715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12927_ _12948_/A _12927_/B vssd1 vssd1 vccd1 vccd1 _17485_/D sky130_fd_sc_hd__and2_1
X_16695_ _18125_/CLK _16695_/D vssd1 vssd1 vccd1 vccd1 _16695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15646_ _17190_/CLK _15646_/D vssd1 vssd1 vccd1 vccd1 _15646_/Q sky130_fd_sc_hd__dfxtp_1
X_18434_ _18437_/CLK _18434_/D vssd1 vssd1 vccd1 vccd1 _18434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12858_ _12864_/A _12858_/B vssd1 vssd1 vccd1 vccd1 _17462_/D sky130_fd_sc_hd__and2_1
XFILLER_0_158_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18365_ _18399_/CLK _18365_/D vssd1 vssd1 vccd1 vccd1 _18365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11809_ hold4670/X _12308_/B _11808_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _11809_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15577_ _17107_/CLK _15577_/D vssd1 vssd1 vccd1 vccd1 _15577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12789_ _12810_/A _12789_/B vssd1 vssd1 vccd1 vccd1 _17439_/D sky130_fd_sc_hd__and2_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _17523_/CLK hold27/X vssd1 vssd1 vccd1 vccd1 _17316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14528_ hold1616/X _14541_/B _14527_/X _14528_/C1 vssd1 vssd1 vccd1 vccd1 _14528_/X
+ sky130_fd_sc_hd__o211a_1
X_18296_ _18296_/CLK _18296_/D vssd1 vssd1 vccd1 vccd1 _18296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17247_ _17247_/CLK _17247_/D vssd1 vssd1 vccd1 vccd1 _17247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14459_ _15193_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14459_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17178_ _17576_/CLK _17178_/D vssd1 vssd1 vccd1 vccd1 _17178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16129_ _16129_/CLK _16129_/D vssd1 vssd1 vccd1 vccd1 hold256/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3106 _18136_/Q vssd1 vssd1 vccd1 vccd1 hold3106/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3117 _07848_/X vssd1 vssd1 vccd1 vccd1 _15569_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08951_ hold452/X hold853/X _08991_/S vssd1 vssd1 vccd1 vccd1 _08952_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_11_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3128 _12824_/X vssd1 vssd1 vccd1 vccd1 _12825_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3139 _17387_/Q vssd1 vssd1 vccd1 vccd1 hold3139/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2405 _13012_/X vssd1 vssd1 vccd1 vccd1 _17514_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2416 _18176_/Q vssd1 vssd1 vccd1 vccd1 hold2416/X sky130_fd_sc_hd__dlygate4sd3_1
X_07902_ _15525_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07902_/X sky130_fd_sc_hd__or2_1
Xhold2427 _07844_/X vssd1 vssd1 vccd1 vccd1 _15567_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08882_ hold29/X hold285/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08883_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_196_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_361_wb_clk_i clkbuf_6_35_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17268_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2438 _15548_/X vssd1 vssd1 vccd1 vccd1 _18452_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1704 _15842_/Q vssd1 vssd1 vccd1 vccd1 hold1704/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2449 _15643_/Q vssd1 vssd1 vccd1 vccd1 hold2449/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1715 _14873_/X vssd1 vssd1 vccd1 vccd1 _18225_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1726 _15691_/Q vssd1 vssd1 vccd1 vccd1 hold1726/X sky130_fd_sc_hd__dlygate4sd3_1
X_07833_ hold915/X _07881_/B vssd1 vssd1 vccd1 vccd1 _07833_/X sky130_fd_sc_hd__or2_1
XFILLER_0_208_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1737 _14213_/X vssd1 vssd1 vccd1 vccd1 _17909_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1748 _16169_/Q vssd1 vssd1 vccd1 vccd1 hold1748/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1759 _14975_/X vssd1 vssd1 vccd1 vccd1 _18273_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09503_ hold2085/X _16325_/Q _10004_/C vssd1 vssd1 vccd1 vccd1 _09504_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_196_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09434_ hold704/X _16303_/Q vssd1 vssd1 vccd1 vccd1 hold714/A sky130_fd_sc_hd__or2_1
XFILLER_0_133_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09365_ _09386_/A _09365_/B _09392_/C _09392_/D vssd1 vssd1 vccd1 vccd1 _09369_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_0_118_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08316_ hold2011/X _08323_/B _08315_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _08316_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_30 _13212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ hold2361/X _09325_/B _09295_/X _12612_/A vssd1 vssd1 vccd1 vccd1 _09296_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_41 _13260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_52 hold87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_63 hold384/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08247_ hold3078/X _08268_/B _08246_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08247_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_74 hold597/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_85 _15145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_96 hold5955/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08178_ hold1877/X _08209_/B _08177_/X _13729_/C1 vssd1 vssd1 vccd1 vccd1 _08178_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5020 _16856_/Q vssd1 vssd1 vccd1 vccd1 hold5020/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5031 _09502_/X vssd1 vssd1 vccd1 vccd1 _16324_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5042 _16612_/Q vssd1 vssd1 vccd1 vccd1 hold5042/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5053 _11296_/X vssd1 vssd1 vccd1 vccd1 _16922_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5064 _16832_/Q vssd1 vssd1 vccd1 vccd1 hold5064/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4330 _16522_/Q vssd1 vssd1 vccd1 vccd1 hold4330/X sky130_fd_sc_hd__buf_2
Xhold5075 _11026_/X vssd1 vssd1 vccd1 vccd1 _16832_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_449_wb_clk_i clkbuf_6_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17723_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10140_ _10524_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10140_/X sky130_fd_sc_hd__or2_1
Xhold4341 _16723_/Q vssd1 vssd1 vccd1 vccd1 hold4341/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5086 _16962_/Q vssd1 vssd1 vccd1 vccd1 hold5086/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4352 _11182_/Y vssd1 vssd1 vccd1 vccd1 _16884_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5097 _17270_/Q vssd1 vssd1 vccd1 vccd1 _12338_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4363 _12304_/Y vssd1 vssd1 vccd1 vccd1 _17258_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4374 _12294_/Y vssd1 vssd1 vccd1 vccd1 _12295_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3640 _16427_/Q vssd1 vssd1 vccd1 vccd1 hold3640/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4385 _11760_/Y vssd1 vssd1 vccd1 vccd1 _11761_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3651 _09667_/X vssd1 vssd1 vccd1 vccd1 _16379_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10071_ _13302_/A _10986_/A _10070_/X vssd1 vssd1 vccd1 vccd1 _10071_/Y sky130_fd_sc_hd__a21oi_1
Xhold4396 _17589_/Q vssd1 vssd1 vccd1 vccd1 hold4396/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3662 _16386_/Q vssd1 vssd1 vccd1 vccd1 hold3662/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3673 _10474_/X vssd1 vssd1 vccd1 vccd1 _16648_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3684 _16560_/Q vssd1 vssd1 vccd1 vccd1 hold3684/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3695 _09613_/X vssd1 vssd1 vccd1 vccd1 _16361_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2950 _18345_/Q vssd1 vssd1 vccd1 vccd1 hold2950/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2961 _14027_/X vssd1 vssd1 vccd1 vccd1 _17819_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2972 _08290_/X vssd1 vssd1 vccd1 vccd1 _15778_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2983 _15856_/Q vssd1 vssd1 vccd1 vccd1 hold2983/X sky130_fd_sc_hd__dlygate4sd3_1
X_13830_ hold4239/X _13734_/A _13829_/X vssd1 vssd1 vccd1 vccd1 _13830_/Y sky130_fd_sc_hd__a21oi_1
Xhold2994 _07838_/X vssd1 vssd1 vccd1 vccd1 _15564_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13761_ _13773_/A _13761_/B vssd1 vssd1 vccd1 vccd1 _13761_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_1382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10973_ hold2646/X hold5066/X _11654_/S vssd1 vssd1 vccd1 vccd1 _10974_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_230_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15500_ _15502_/A _15500_/B vssd1 vssd1 vccd1 vccd1 _18429_/D sky130_fd_sc_hd__and2_1
X_12712_ _16235_/Q _17415_/Q _12766_/S vssd1 vssd1 vccd1 vccd1 _12712_/X sky130_fd_sc_hd__mux2_1
X_16480_ _16480_/CLK _16480_/D vssd1 vssd1 vccd1 vccd1 _16480_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _13788_/A _13692_/B vssd1 vssd1 vccd1 vccd1 _13692_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15431_ hold518/X _15441_/A2 _09386_/D hold411/X _15426_/X vssd1 vssd1 vccd1 vccd1
+ _15432_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_210_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12643_ hold2904/X hold3343/X _12844_/S vssd1 vssd1 vccd1 vccd1 _12643_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_167_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18150_ _18150_/CLK _18150_/D vssd1 vssd1 vccd1 vccd1 _18150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15362_ _15480_/A _15362_/B _15362_/C _15362_/D vssd1 vssd1 vccd1 vccd1 _15362_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12574_ hold1996/X _17369_/Q _12970_/S vssd1 vssd1 vccd1 vccd1 _12574_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_142_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17101_ _17261_/CLK _17101_/D vssd1 vssd1 vccd1 vccd1 _17101_/Q sky130_fd_sc_hd__dfxtp_1
X_14313_ hold2701/X _14333_/A2 _14312_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _14313_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18081_ _18081_/CLK _18081_/D vssd1 vssd1 vccd1 vccd1 _18081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11525_ hold2189/X hold5669/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11526_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15293_ _15490_/A1 _15285_/X _15292_/X _15490_/B1 hold5935/A vssd1 vssd1 vccd1 vccd1
+ _15293_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_108_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17032_ _18448_/CLK _17032_/D vssd1 vssd1 vccd1 vccd1 _17032_/Q sky130_fd_sc_hd__dfxtp_1
X_14244_ hold423/X _14284_/B vssd1 vssd1 vccd1 vccd1 _14244_/X sky130_fd_sc_hd__or2_1
XFILLER_0_223_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11456_ hold2526/X _16976_/Q _12317_/C vssd1 vssd1 vccd1 vccd1 _11457_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10407_ _11103_/A _10407_/B vssd1 vssd1 vccd1 vccd1 _10407_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14175_ hold2487/X _14198_/B _14174_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _14175_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11387_ hold1676/X _16953_/Q _11783_/C vssd1 vssd1 vccd1 vccd1 _11388_/B sky130_fd_sc_hd__mux2_1
X_13126_ _13126_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13126_/X sky130_fd_sc_hd__or2_1
X_10338_ _10470_/A _10338_/B vssd1 vssd1 vccd1 vccd1 _10338_/X sky130_fd_sc_hd__or2_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_119_wb_clk_i clkbuf_6_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16120_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _13055_/C _13057_/B _17521_/Q vssd1 vssd1 vccd1 vccd1 _13057_/X sky130_fd_sc_hd__and3b_4
X_17934_ _18345_/CLK _17934_/D vssd1 vssd1 vccd1 vccd1 _17934_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10269_ _11091_/A _10269_/B vssd1 vssd1 vccd1 vccd1 _10269_/X sky130_fd_sc_hd__or2_1
X_12008_ hold1229/X hold4654/X _13811_/C vssd1 vssd1 vccd1 vccd1 _12009_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_84_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17865_ _17865_/CLK _17865_/D vssd1 vssd1 vccd1 vccd1 _17865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16816_ _18051_/CLK _16816_/D vssd1 vssd1 vccd1 vccd1 _16816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_1352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17796_ _17862_/CLK _17796_/D vssd1 vssd1 vccd1 vccd1 _17796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16747_ _18072_/CLK _16747_/D vssd1 vssd1 vccd1 vccd1 _16747_/Q sky130_fd_sc_hd__dfxtp_1
X_13959_ hold1656/X _13995_/A2 _13958_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _13959_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16678_ _18164_/CLK _16678_/D vssd1 vssd1 vccd1 vccd1 _16678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18417_ _18417_/CLK _18417_/D vssd1 vssd1 vccd1 vccd1 _18417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15629_ _18447_/CLK _15629_/D vssd1 vssd1 vccd1 vccd1 _15629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09150_ _15533_/A _09156_/B vssd1 vssd1 vccd1 vccd1 _09150_/X sky130_fd_sc_hd__or2_1
X_18348_ _18372_/CLK _18348_/D vssd1 vssd1 vccd1 vccd1 _18348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08101_ hold955/X _08088_/B _08100_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 hold956/A
+ sky130_fd_sc_hd__o211a_1
X_18279_ _18357_/CLK _18279_/D vssd1 vssd1 vccd1 vccd1 _18279_/Q sky130_fd_sc_hd__dfxtp_1
X_09081_ hold2914/X _09106_/B _09080_/X _12987_/A vssd1 vssd1 vccd1 vccd1 _09081_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08032_ hold2509/X _08033_/B _08031_/Y _13933_/A vssd1 vssd1 vccd1 vccd1 _08032_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput50 input50/A vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_6
XFILLER_0_31_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput61 input61/A vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__buf_6
Xhold801 hold801/A vssd1 vssd1 vccd1 vccd1 hold801/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold812 hold812/A vssd1 vssd1 vccd1 vccd1 hold812/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold823 hold823/A vssd1 vssd1 vccd1 vccd1 hold823/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold834 hold834/A vssd1 vssd1 vccd1 vccd1 hold834/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold845 hold845/A vssd1 vssd1 vccd1 vccd1 hold845/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold856 hold856/A vssd1 vssd1 vccd1 vccd1 hold856/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 hold867/A vssd1 vssd1 vccd1 vccd1 hold867/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold878 hold878/A vssd1 vssd1 vccd1 vccd1 hold878/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09983_ hold1722/X _16485_/Q _10004_/C vssd1 vssd1 vccd1 vccd1 _09984_/B sky130_fd_sc_hd__mux2_1
Xhold889 hold889/A vssd1 vssd1 vccd1 vccd1 hold889/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2202 _15540_/X vssd1 vssd1 vccd1 vccd1 _18448_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08934_ _08934_/A _12445_/B vssd1 vssd1 vccd1 vccd1 _08934_/X sky130_fd_sc_hd__or2_2
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2213 _18375_/Q vssd1 vssd1 vccd1 vccd1 hold2213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2224 _18311_/Q vssd1 vssd1 vccd1 vccd1 hold2224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2235 _08192_/X vssd1 vssd1 vccd1 vccd1 _15732_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2246 _15862_/Q vssd1 vssd1 vccd1 vccd1 hold2246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1501 _17957_/Q vssd1 vssd1 vccd1 vccd1 hold1501/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1512 _14071_/X vssd1 vssd1 vccd1 vccd1 _17840_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08865_ _15473_/A _08865_/B vssd1 vssd1 vccd1 vccd1 _16051_/D sky130_fd_sc_hd__and2_1
Xhold2257 _18330_/Q vssd1 vssd1 vccd1 vccd1 hold2257/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2268 next_key vssd1 vssd1 vccd1 vccd1 hold2268/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1523 _18033_/Q vssd1 vssd1 vccd1 vccd1 hold1523/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2279 _18077_/Q vssd1 vssd1 vccd1 vccd1 hold2279/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 _17896_/Q vssd1 vssd1 vccd1 vccd1 hold1534/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1545 _08081_/X vssd1 vssd1 vccd1 vccd1 _15680_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07816_ _15515_/A _14972_/A _14166_/A hold927/X vssd1 vssd1 vccd1 vccd1 _07817_/D
+ sky130_fd_sc_hd__or4_1
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1556 _15601_/Q vssd1 vssd1 vccd1 vccd1 hold1556/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1567 _08306_/X vssd1 vssd1 vccd1 vccd1 _15786_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08796_ _08868_/B _08934_/A _13046_/D vssd1 vssd1 vccd1 vccd1 _08801_/S sky130_fd_sc_hd__or3_2
XFILLER_0_74_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1578 hold1756/X vssd1 vssd1 vccd1 vccd1 hold1757/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1589 _14303_/X vssd1 vssd1 vccd1 vccd1 _17951_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09417_ _07804_/A _09456_/A _09440_/B _09416_/X vssd1 vssd1 vccd1 vccd1 _09417_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09348_ hold597/A _15541_/A _15182_/A _09352_/D vssd1 vssd1 vccd1 vccd1 _09364_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_47_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09279_ _15555_/A hold980/X _09283_/S vssd1 vssd1 vccd1 vccd1 hold981/A sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11310_ _11694_/A _11310_/B vssd1 vssd1 vccd1 vccd1 _11310_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12290_ hold1429/X _17254_/Q _13796_/S vssd1 vssd1 vccd1 vccd1 _12291_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11241_ _12210_/A _11241_/B vssd1 vssd1 vccd1 vccd1 _11241_/X sky130_fd_sc_hd__or2_1
XFILLER_0_142_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_283_wb_clk_i clkbuf_6_50_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18031_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11172_ hold4251/X _11010_/A _11171_/X vssd1 vssd1 vccd1 vccd1 _11172_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_212_wb_clk_i clkbuf_6_54_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18206_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4160 _11668_/X vssd1 vssd1 vccd1 vccd1 _17046_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10123_ hold3840/X _10601_/B _10122_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10123_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4171 _16406_/Q vssd1 vssd1 vccd1 vccd1 hold4171/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4182 _15263_/X vssd1 vssd1 vccd1 vccd1 _15264_/B sky130_fd_sc_hd__dlygate4sd3_1
X_15980_ _17295_/CLK _15980_/D vssd1 vssd1 vccd1 vccd1 hold869/A sky130_fd_sc_hd__dfxtp_1
XTAP_6355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4193 hold5911/X vssd1 vssd1 vccd1 vccd1 hold5912/A sky130_fd_sc_hd__buf_4
XTAP_6366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3470 _17100_/Q vssd1 vssd1 vccd1 vccd1 hold3470/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14931_ hold3100/X _14946_/B _14930_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _14931_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3481 hold3984/X vssd1 vssd1 vccd1 vccd1 _10589_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10054_ _11206_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _10054_/Y sky130_fd_sc_hd__nor2_1
XTAP_5654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3492 _11185_/Y vssd1 vssd1 vccd1 vccd1 _16885_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2780 _14035_/X vssd1 vssd1 vccd1 vccd1 _17823_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14862_ _15201_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14862_/X sky130_fd_sc_hd__or2_1
X_17650_ _17705_/CLK _17650_/D vssd1 vssd1 vccd1 vccd1 _17650_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2791 _08200_/X vssd1 vssd1 vccd1 vccd1 _15736_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16601_ _18191_/CLK _16601_/D vssd1 vssd1 vccd1 vccd1 _16601_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13813_ _13819_/A _13813_/B vssd1 vssd1 vccd1 vccd1 _13813_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_230_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17581_ _17741_/CLK _17581_/D vssd1 vssd1 vccd1 vccd1 _17581_/Q sky130_fd_sc_hd__dfxtp_1
X_14793_ hold1899/X _14828_/B _14792_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _14793_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16532_ _18220_/CLK _16532_/D vssd1 vssd1 vccd1 vccd1 _16532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13744_ hold5203/X _13856_/B _13743_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13744_/X
+ sky130_fd_sc_hd__o211a_1
X_10956_ _11136_/A _10956_/B vssd1 vssd1 vccd1 vccd1 _10956_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16463_ _18250_/CLK _16463_/D vssd1 vssd1 vccd1 vccd1 _16463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13675_ hold4048/X _13795_/A2 _13674_/X _13675_/C1 vssd1 vssd1 vccd1 vccd1 _13675_/X
+ sky130_fd_sc_hd__o211a_1
X_10887_ _11100_/A _10887_/B vssd1 vssd1 vccd1 vccd1 _10887_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15414_ _15414_/A _15414_/B vssd1 vssd1 vccd1 vccd1 _18417_/D sky130_fd_sc_hd__and2_1
XFILLER_0_155_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18202_ _18222_/CLK _18202_/D vssd1 vssd1 vccd1 vccd1 _18202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_241_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12626_ hold2277/X _12625_/X _12626_/S vssd1 vssd1 vccd1 vccd1 _12626_/X sky130_fd_sc_hd__mux2_1
XPHY_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16394_ _18371_/CLK _16394_/D vssd1 vssd1 vccd1 vccd1 _16394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_241_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18133_ _18215_/CLK _18133_/D vssd1 vssd1 vccd1 vccd1 _18133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15345_ hold478/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15345_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12557_ hold3599/X _12556_/X _12929_/S vssd1 vssd1 vccd1 vccd1 _12557_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11508_ _12174_/A _11508_/B vssd1 vssd1 vccd1 vccd1 _11508_/X sky130_fd_sc_hd__or2_1
X_18064_ _18064_/CLK _18064_/D vssd1 vssd1 vccd1 vccd1 _18064_/Q sky130_fd_sc_hd__dfxtp_1
X_15276_ _17331_/Q _15486_/B1 _15485_/B1 _16108_/Q vssd1 vssd1 vccd1 vccd1 _15276_/X
+ sky130_fd_sc_hd__a22o_1
X_12488_ _17337_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12488_/X sky130_fd_sc_hd__or2_1
Xhold108 hold108/A vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__buf_12
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17015_ _17895_/CLK _17015_/D vssd1 vssd1 vccd1 vccd1 _17015_/Q sky130_fd_sc_hd__dfxtp_1
Xhold119 hold119/A vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14227_ hold1117/X _14216_/Y _14226_/X _14354_/A vssd1 vssd1 vccd1 vccd1 _14227_/X
+ sky130_fd_sc_hd__o211a_1
X_11439_ _11631_/A _11439_/B vssd1 vssd1 vccd1 vccd1 _11439_/X sky130_fd_sc_hd__or2_1
XFILLER_0_112_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14158_ _15557_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14158_/X sky130_fd_sc_hd__or2_1
XFILLER_0_237_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13109_ _13108_/X hold4330/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13109_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14089_ hold3012/X _14094_/B _14088_/Y _12894_/A vssd1 vssd1 vccd1 vccd1 _14089_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_225_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_238_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17917_ _17949_/CLK _17917_/D vssd1 vssd1 vccd1 vccd1 _17917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_218_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_234_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08650_ _15344_/A _08650_/B vssd1 vssd1 vccd1 vccd1 _15947_/D sky130_fd_sc_hd__and2_1
X_17848_ _18429_/CLK _17848_/D vssd1 vssd1 vccd1 vccd1 _17848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08581_ _15414_/A _08581_/B vssd1 vssd1 vccd1 vccd1 _15914_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_87_wb_clk_i clkbuf_6_17_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17509_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17779_ _17779_/CLK _17779_/D vssd1 vssd1 vccd1 vccd1 _17779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_wb_clk_i clkbuf_6_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18438_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09202_ _15531_/A _09206_/B vssd1 vssd1 vccd1 vccd1 _09202_/X sky130_fd_sc_hd__or2_1
XFILLER_0_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09133_ hold2931/X _09177_/A2 _09132_/X _12864_/A vssd1 vssd1 vccd1 vccd1 _09133_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09064_ _18461_/Q hold353/A vssd1 vssd1 vccd1 vccd1 hold268/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08015_ _15529_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08015_/X sky130_fd_sc_hd__or2_1
XFILLER_0_128_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold620 hold620/A vssd1 vssd1 vccd1 vccd1 hold620/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold631 hold631/A vssd1 vssd1 vccd1 vccd1 hold631/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold642 hold642/A vssd1 vssd1 vccd1 vccd1 hold642/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold653 hold653/A vssd1 vssd1 vccd1 vccd1 hold653/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold664 hold664/A vssd1 vssd1 vccd1 vccd1 hold664/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold675 hold675/A vssd1 vssd1 vccd1 vccd1 hold675/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 hold686/A vssd1 vssd1 vccd1 vccd1 hold686/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold697 hold697/A vssd1 vssd1 vccd1 vccd1 hold697/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09966_ _10482_/A _09966_/B vssd1 vssd1 vccd1 vccd1 _09966_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2010 _15003_/X vssd1 vssd1 vccd1 vccd1 _18287_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2021 _18148_/Q vssd1 vssd1 vccd1 vccd1 hold2021/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08917_ _15244_/A hold467/X vssd1 vssd1 vccd1 vccd1 _16076_/D sky130_fd_sc_hd__and2_1
Xhold2032 _09115_/X vssd1 vssd1 vccd1 vccd1 _16172_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2043 _15828_/Q vssd1 vssd1 vccd1 vccd1 hold2043/X sky130_fd_sc_hd__dlygate4sd3_1
X_09897_ _09987_/A _09897_/B vssd1 vssd1 vccd1 vccd1 _09897_/X sky130_fd_sc_hd__or2_1
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2054 _14189_/X vssd1 vssd1 vccd1 vccd1 _17897_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2065 _14795_/X vssd1 vssd1 vccd1 vccd1 _18187_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1320 _09177_/X vssd1 vssd1 vccd1 vccd1 _16201_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1331 _08432_/X vssd1 vssd1 vccd1 vccd1 _15846_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2076 _14965_/X vssd1 vssd1 vccd1 vccd1 _18269_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ hold53/X hold656/X _08866_/S vssd1 vssd1 vccd1 vccd1 _08849_/B sky130_fd_sc_hd__mux2_1
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2087 _14534_/X vssd1 vssd1 vccd1 vccd1 _18063_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1342 _18020_/Q vssd1 vssd1 vccd1 vccd1 hold1342/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2098 _18017_/Q vssd1 vssd1 vccd1 vccd1 hold2098/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1353 _08042_/X vssd1 vssd1 vccd1 vccd1 _15662_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1364 hold6119/X vssd1 vssd1 vccd1 vccd1 hold909/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1375 _15152_/X vssd1 vssd1 vccd1 vccd1 _18359_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1386 _16158_/Q vssd1 vssd1 vccd1 vccd1 hold1386/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ hold143/X hold574/X _08779_/S vssd1 vssd1 vccd1 vccd1 _08780_/B sky130_fd_sc_hd__mux2_1
Xhold1397 _15738_/Q vssd1 vssd1 vccd1 vccd1 hold1397/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10810_ hold5535/X _11213_/B _10809_/X _14342_/A vssd1 vssd1 vccd1 vccd1 _10810_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ hold4390/X _11694_/A _11789_/X vssd1 vssd1 vccd1 vccd1 _11790_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_212_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10741_ hold3917/X _11222_/B _10740_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _10741_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13460_ hold2922/X hold4985/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13461_/B sky130_fd_sc_hd__mux2_1
X_10672_ hold5446/X _11723_/B _10671_/X _14364_/A vssd1 vssd1 vccd1 vccd1 _10672_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12411_ hold180/X hold770/X _12441_/S vssd1 vssd1 vccd1 vccd1 hold771/A sky130_fd_sc_hd__mux2_1
XFILLER_0_91_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13391_ hold2394/X hold4367/X _13865_/C vssd1 vssd1 vccd1 vccd1 _13392_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_106_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_464_wb_clk_i clkbuf_6_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17440_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_106_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15130_ hold1833/X _15165_/B _15129_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _15130_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12342_ hold4306/X _13407_/A _12341_/X vssd1 vssd1 vccd1 vccd1 _12342_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15061_ _15169_/A hold1179/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15062_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12273_ _12273_/A _12273_/B vssd1 vssd1 vccd1 vccd1 _12273_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14012_ _15519_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14012_/X sky130_fd_sc_hd__or2_1
X_11224_ _12331_/A _11224_/B vssd1 vssd1 vccd1 vccd1 _11224_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11155_ _11158_/A _11155_/B vssd1 vssd1 vccd1 vccd1 _11155_/Y sky130_fd_sc_hd__nor2_1
XTAP_6141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10106_ hold3163/X hold3486/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10107_/B sky130_fd_sc_hd__mux2_1
XTAP_6174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15963_ _16090_/CLK _15963_/D vssd1 vssd1 vccd1 vccd1 hold856/A sky130_fd_sc_hd__dfxtp_1
XTAP_5440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11086_ hold5245/X _11186_/B _11085_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _11086_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17702_ _17702_/CLK _17702_/D vssd1 vssd1 vccd1 vccd1 _17702_/Q sky130_fd_sc_hd__dfxtp_1
X_10037_ _16503_/Q _10577_/B _10385_/S vssd1 vssd1 vccd1 vccd1 _10037_/X sky130_fd_sc_hd__and3_1
X_14914_ _15183_/A hold407/X vssd1 vssd1 vccd1 vccd1 _14914_/X sky130_fd_sc_hd__or2_1
X_15894_ _17344_/CLK _15894_/D vssd1 vssd1 vccd1 vccd1 hold324/A sky130_fd_sc_hd__dfxtp_1
XTAP_5484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ _17729_/CLK _17633_/D vssd1 vssd1 vccd1 vccd1 _17633_/Q sky130_fd_sc_hd__dfxtp_1
X_14845_ hold2169/X _14880_/B _14844_/X _14853_/C1 vssd1 vssd1 vccd1 vccd1 _14845_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_231_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_231_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14776_ _15169_/A _14780_/B vssd1 vssd1 vccd1 vccd1 _14776_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17564_ _17628_/CLK _17564_/D vssd1 vssd1 vccd1 vccd1 _17564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11988_ _12273_/A _11988_/B vssd1 vssd1 vccd1 vccd1 _11988_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16515_ _18298_/CLK _16515_/D vssd1 vssd1 vccd1 vccd1 _16515_/Q sky130_fd_sc_hd__dfxtp_1
X_13727_ hold1877/X _17696_/Q _13766_/S vssd1 vssd1 vccd1 vccd1 _13728_/B sky130_fd_sc_hd__mux2_1
X_10939_ hold3927/X _11222_/B _10938_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _16803_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_188_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17495_ _17500_/CLK _17495_/D vssd1 vssd1 vccd1 vccd1 _17495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16446_ _18391_/CLK _16446_/D vssd1 vssd1 vccd1 vccd1 _16446_/Q sky130_fd_sc_hd__dfxtp_1
X_13658_ hold2400/X hold5557/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13659_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_45_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12609_ _12612_/A _12609_/B vssd1 vssd1 vccd1 vccd1 _17379_/D sky130_fd_sc_hd__and2_1
X_16377_ _18386_/CLK _16377_/D vssd1 vssd1 vccd1 vccd1 _16377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13589_ hold1037/X hold4125/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13590_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15328_ hold592/X _15484_/A2 _09392_/D hold810/X vssd1 vssd1 vccd1 vccd1 _15328_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18116_ _18154_/CLK _18116_/D vssd1 vssd1 vccd1 vccd1 _18116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_134_wb_clk_i clkbuf_6_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17345_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5608 _17705_/Q vssd1 vssd1 vccd1 vccd1 hold5608/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5619 _10912_/X vssd1 vssd1 vccd1 vccd1 _16794_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15259_ hold608/X _15485_/A2 _15488_/A2 hold830/X _15258_/X vssd1 vssd1 vccd1 vccd1
+ _15262_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_151_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18047_ _18047_/CLK hold637/X vssd1 vssd1 vccd1 vccd1 hold636/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4907 _16764_/Q vssd1 vssd1 vccd1 vccd1 hold4907/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4918 _11983_/X vssd1 vssd1 vccd1 vccd1 _17151_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4929 _16890_/Q vssd1 vssd1 vccd1 vccd1 hold4929/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09820_ hold5823/X _10022_/B _09819_/X _15202_/C1 vssd1 vssd1 vccd1 vccd1 _09820_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout407 _14286_/Y vssd1 vssd1 vccd1 vccd1 _14333_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_201_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout418 _14106_/B vssd1 vssd1 vccd1 vccd1 _14104_/B sky130_fd_sc_hd__buf_6
XFILLER_0_123_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout429 _13307_/S vssd1 vssd1 vccd1 vccd1 _13251_/S sky130_fd_sc_hd__buf_8
XFILLER_0_226_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_225_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09751_ hold3276/X _10577_/B _09750_/X _15146_/C1 vssd1 vssd1 vccd1 vccd1 _09751_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_197_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08702_ _15314_/A _08702_/B vssd1 vssd1 vccd1 vccd1 _15972_/D sky130_fd_sc_hd__and2_1
XFILLER_0_241_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09682_ hold3903/X _10046_/B _09681_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09682_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_234_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08633_ hold254/X hold472/X _08657_/S vssd1 vssd1 vccd1 vccd1 _08634_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ hold185/X hold745/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold746/A sky130_fd_sc_hd__mux2_1
XFILLER_0_77_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_234_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08495_ hold2575/X _08486_/B _08494_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _08495_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09116_ _15231_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09116_/X sky130_fd_sc_hd__or2_1
XFILLER_0_115_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09047_ _09047_/A hold139/X vssd1 vssd1 vccd1 vccd1 _16140_/D sky130_fd_sc_hd__and2_1
Xhold450 hold450/A vssd1 vssd1 vccd1 vccd1 input35/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 hold461/A vssd1 vssd1 vccd1 vccd1 hold461/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 hold472/A vssd1 vssd1 vccd1 vccd1 hold472/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold483 input49/X vssd1 vssd1 vccd1 vccd1 hold483/X sky130_fd_sc_hd__clkbuf_2
Xhold494 input26/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__buf_1
XFILLER_0_217_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout930 hold630/X vssd1 vssd1 vccd1 vccd1 _15537_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout941 hold1007/X vssd1 vssd1 vccd1 vccd1 _15205_/A sky130_fd_sc_hd__clkbuf_4
X_09949_ hold4707/X _10031_/B _09948_/X _15146_/C1 vssd1 vssd1 vccd1 vccd1 _09949_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ _14358_/A _12960_/B vssd1 vssd1 vccd1 vccd1 _17496_/D sky130_fd_sc_hd__and2_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 _09302_/X vssd1 vssd1 vccd1 vccd1 _16261_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1161 _15879_/Q vssd1 vssd1 vccd1 vccd1 hold1161/X sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ hold5028/X _13811_/B _11910_/X _08363_/A vssd1 vssd1 vccd1 vccd1 _11911_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_217_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1172 _15813_/Q vssd1 vssd1 vccd1 vccd1 hold1172/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1183 hold691/X vssd1 vssd1 vccd1 vccd1 hold1183/X sky130_fd_sc_hd__clkbuf_8
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _12894_/A _12891_/B vssd1 vssd1 vccd1 vccd1 _17473_/D sky130_fd_sc_hd__and2_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 _14164_/A vssd1 vssd1 vccd1 vccd1 _15509_/A sky130_fd_sc_hd__buf_4
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _15185_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14630_/X sky130_fd_sc_hd__or2_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ hold3854/X _12353_/B _11841_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _11842_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ hold915/X _14557_/Y _14560_/X _15019_/C1 vssd1 vssd1 vccd1 vccd1 hold916/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _12331_/A _11773_/B vssd1 vssd1 vccd1 vccd1 _11773_/Y sky130_fd_sc_hd__nor2_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _16319_/CLK hold734/X vssd1 vssd1 vccd1 vccd1 _16300_/Q sky130_fd_sc_hd__dfxtp_1
X_13512_ _13722_/A _13512_/B vssd1 vssd1 vccd1 vccd1 _13512_/X sky130_fd_sc_hd__or2_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10724_ hold2347/X hold4326/X _11204_/C vssd1 vssd1 vccd1 vccd1 _10725_/B sky130_fd_sc_hd__mux2_1
X_17280_ _17280_/CLK _17280_/D vssd1 vssd1 vccd1 vccd1 _17280_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ hold1956/X _14487_/B _14491_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _14492_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16231_ _17753_/CLK _16231_/D vssd1 vssd1 vccd1 vccd1 _16231_/Q sky130_fd_sc_hd__dfxtp_1
X_13443_ _13737_/A _13443_/B vssd1 vssd1 vccd1 vccd1 _13443_/X sky130_fd_sc_hd__or2_1
XFILLER_0_148_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10655_ hold2163/X hold4634/X _11732_/C vssd1 vssd1 vccd1 vccd1 _10656_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_64_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16162_ _18042_/CLK _16162_/D vssd1 vssd1 vccd1 vccd1 _16162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13374_ _13758_/A _13374_/B vssd1 vssd1 vccd1 vccd1 _13374_/X sky130_fd_sc_hd__or2_1
XFILLER_0_51_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10586_ _16686_/Q _10625_/B _10625_/C vssd1 vssd1 vccd1 vccd1 _10586_/X sky130_fd_sc_hd__and3_1
XFILLER_0_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15113_ _15547_/A hold340/X vssd1 vssd1 vccd1 vccd1 _15113_/Y sky130_fd_sc_hd__nand2_1
X_12325_ _13873_/A _12325_/B vssd1 vssd1 vccd1 vccd1 _12325_/Y sky130_fd_sc_hd__nor2_1
X_16093_ _16093_/CLK _16093_/D vssd1 vssd1 vccd1 vccd1 hold853/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15044_ _15044_/A _15044_/B vssd1 vssd1 vccd1 vccd1 _18307_/D sky130_fd_sc_hd__and2_1
XFILLER_0_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12256_ hold5793/X _12350_/B _12255_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _12256_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11207_ _11207_/A _11222_/B _11789_/C vssd1 vssd1 vccd1 vccd1 _11207_/X sky130_fd_sc_hd__and3_1
XFILLER_0_76_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12187_ hold5255/X _13886_/B _12186_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _12187_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11138_ _18073_/Q _16870_/Q _11723_/C vssd1 vssd1 vccd1 vccd1 _11139_/B sky130_fd_sc_hd__mux2_1
X_16995_ _17904_/CLK _16995_/D vssd1 vssd1 vccd1 vccd1 _16995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_235_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15946_ _17293_/CLK _15946_/D vssd1 vssd1 vccd1 vccd1 hold592/A sky130_fd_sc_hd__dfxtp_1
XTAP_5270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11069_ hold1855/X _16847_/Q _11168_/C vssd1 vssd1 vccd1 vccd1 _11070_/B sky130_fd_sc_hd__mux2_1
XTAP_5281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15877_ _17620_/CLK _15877_/D vssd1 vssd1 vccd1 vccd1 _15877_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17616_ _17648_/CLK _17616_/D vssd1 vssd1 vccd1 vccd1 _17616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14828_ _14952_/A _14828_/B vssd1 vssd1 vccd1 vccd1 _14828_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_188_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17547_ _18081_/CLK _17547_/D vssd1 vssd1 vccd1 vccd1 _17547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14759_ hold1919/X _14774_/B _14758_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14759_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_386_wb_clk_i clkbuf_6_35_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17277_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08280_ _15559_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08280_/X sky130_fd_sc_hd__or2_1
XFILLER_0_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17478_ _17481_/CLK _17478_/D vssd1 vssd1 vccd1 vccd1 _17478_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_315_wb_clk_i clkbuf_6_47_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18061_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16429_ _18374_/CLK _16429_/D vssd1 vssd1 vccd1 vccd1 _16429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6106 la_data_in[1] vssd1 vssd1 vccd1 vccd1 hold6106/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6117 _16519_/Q vssd1 vssd1 vccd1 vccd1 hold6117/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6128 _16317_/Q vssd1 vssd1 vccd1 vccd1 hold739/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5405 _11506_/X vssd1 vssd1 vccd1 vccd1 _16992_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5416 _17745_/Q vssd1 vssd1 vccd1 vccd1 hold5416/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5427 _11410_/X vssd1 vssd1 vccd1 vccd1 _16960_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5438 _17740_/Q vssd1 vssd1 vccd1 vccd1 hold5438/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5449 _10831_/X vssd1 vssd1 vccd1 vccd1 _16767_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4704 _13441_/X vssd1 vssd1 vccd1 vccd1 _17600_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4715 _17659_/Q vssd1 vssd1 vccd1 vccd1 hold4715/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4726 _09802_/X vssd1 vssd1 vccd1 vccd1 _16424_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4737 _17721_/Q vssd1 vssd1 vccd1 vccd1 hold4737/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4748 _12995_/X vssd1 vssd1 vccd1 vccd1 _12996_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4759 _13438_/X vssd1 vssd1 vccd1 vccd1 _17599_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout204 _11792_/B vssd1 vssd1 vccd1 vccd1 _12335_/B sky130_fd_sc_hd__buf_4
Xfanout215 _09992_/B vssd1 vssd1 vccd1 vccd1 _10022_/B sky130_fd_sc_hd__buf_4
Xfanout226 _10634_/B vssd1 vssd1 vccd1 vccd1 _10598_/B sky130_fd_sc_hd__buf_4
XFILLER_0_22_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout237 _10577_/B vssd1 vssd1 vccd1 vccd1 _10049_/B sky130_fd_sc_hd__clkbuf_8
X_09803_ hold2752/X hold3746/X _10028_/C vssd1 vssd1 vccd1 vccd1 _09804_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_226_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout248 _13722_/A vssd1 vssd1 vccd1 vccd1 _13719_/A sky130_fd_sc_hd__buf_4
Xfanout259 fanout299/X vssd1 vssd1 vccd1 vccd1 _12216_/A sky130_fd_sc_hd__clkbuf_4
X_07995_ _14395_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _07995_/X sky130_fd_sc_hd__or2_1
XFILLER_0_201_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09734_ _18315_/Q _16402_/Q _11171_/C vssd1 vssd1 vccd1 vccd1 _09735_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_96_1349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_31_wb_clk_i clkbuf_6_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17981_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_119_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09665_ hold2699/X hold3237/X _10067_/C vssd1 vssd1 vccd1 vccd1 _09666_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_210_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08616_ _15374_/A hold453/X vssd1 vssd1 vccd1 vccd1 _15930_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09596_ hold2075/X hold5030/X _09992_/C vssd1 vssd1 vccd1 vccd1 _09597_/B sky130_fd_sc_hd__mux2_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _12420_/A hold680/X vssd1 vssd1 vccd1 vccd1 _15897_/D sky130_fd_sc_hd__and2_1
XFILLER_0_221_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08478_ _14477_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08478_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10440_ _10536_/A _10440_/B vssd1 vssd1 vccd1 vccd1 _10440_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_30_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_30_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_116_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10371_ _10530_/A _10371_/B vssd1 vssd1 vccd1 vccd1 _10371_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12110_ hold2648/X _17194_/Q _12293_/C vssd1 vssd1 vccd1 vccd1 _12111_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5950 hold5950/A vssd1 vssd1 vccd1 vccd1 hold5950/X sky130_fd_sc_hd__clkbuf_4
X_13090_ _17562_/Q _17096_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13090_/X sky130_fd_sc_hd__mux2_1
Xhold5961 hold5961/A vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_12
XFILLER_0_130_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5972 hold6089/X vssd1 vssd1 vccd1 vccd1 hold5972/X sky130_fd_sc_hd__clkbuf_4
Xhold5983 hold6125/X vssd1 vssd1 vccd1 vccd1 _09463_/C sky130_fd_sc_hd__buf_1
Xhold5994 _16306_/Q vssd1 vssd1 vccd1 vccd1 hold5994/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12041_ hold2173/X _17171_/Q _12329_/C vssd1 vssd1 vccd1 vccd1 _12042_/B sky130_fd_sc_hd__mux2_1
Xhold280 hold280/A vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 hold291/A vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout760 _14131_/C1 vssd1 vssd1 vccd1 vccd1 _13923_/A sky130_fd_sc_hd__buf_4
XFILLER_0_205_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15800_ _17697_/CLK _15800_/D vssd1 vssd1 vccd1 vccd1 _15800_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout771 fanout791/X vssd1 vssd1 vccd1 vccd1 _08131_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_232_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout782 _14526_/C1 vssd1 vssd1 vccd1 vccd1 _14348_/A sky130_fd_sc_hd__buf_4
XFILLER_0_204_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16780_ _17983_/CLK _16780_/D vssd1 vssd1 vccd1 vccd1 _16780_/Q sky130_fd_sc_hd__dfxtp_1
X_13992_ _15553_/A _13994_/B vssd1 vssd1 vccd1 vccd1 _13992_/X sky130_fd_sc_hd__or2_1
Xfanout793 _15056_/A vssd1 vssd1 vccd1 vccd1 _15072_/A sky130_fd_sc_hd__buf_4
XFILLER_0_217_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12943_ hold2914/X hold4441/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12943_/X sky130_fd_sc_hd__mux2_1
X_15731_ _17734_/CLK _15731_/D vssd1 vssd1 vccd1 vccd1 _15731_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18450_ _18451_/CLK _18450_/D vssd1 vssd1 vccd1 vccd1 _18450_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 hold933/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15662_ _17906_/CLK _15662_/D vssd1 vssd1 vccd1 vccd1 _15662_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ hold1338/X _17469_/Q _12916_/S vssd1 vssd1 vccd1 vccd1 _12874_/X sky130_fd_sc_hd__mux2_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _18452_/CLK _17401_/D vssd1 vssd1 vccd1 vccd1 _17401_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ hold2380/X _14612_/B _14612_/Y _14697_/C1 vssd1 vssd1 vccd1 vccd1 _14613_/X
+ sky130_fd_sc_hd__o211a_1
X_11825_ hold1726/X hold4471/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11826_/B sky130_fd_sc_hd__mux2_1
X_18381_ _18381_/CLK _18381_/D vssd1 vssd1 vccd1 vccd1 _18381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15593_ _17209_/CLK _15593_/D vssd1 vssd1 vccd1 vccd1 _15593_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17332_ _17336_/CLK hold15/X vssd1 vssd1 vccd1 vccd1 _17332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ hold1127/X _14541_/B _14543_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _14544_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _17076_/Q _11771_/B _12242_/S vssd1 vssd1 vccd1 vccd1 _11756_/X sky130_fd_sc_hd__and3_1
XFILLER_0_154_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _11091_/A _10707_/B vssd1 vssd1 vccd1 vccd1 _10707_/X sky130_fd_sc_hd__or2_1
X_14475_ _14529_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14475_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17263_ _17899_/CLK _17263_/D vssd1 vssd1 vccd1 vccd1 _17263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11687_ hold3014/X hold5677/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11688_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_148_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13426_ hold5763/X _13814_/B _13425_/X _08361_/A vssd1 vssd1 vccd1 vccd1 _13426_/X
+ sky130_fd_sc_hd__o211a_1
X_16214_ _17723_/CLK _16214_/D vssd1 vssd1 vccd1 vccd1 _16214_/Q sky130_fd_sc_hd__dfxtp_1
X_10638_ hold3473/X _10542_/A _10637_/X vssd1 vssd1 vccd1 vccd1 _10638_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17194_ _17194_/CLK _17194_/D vssd1 vssd1 vccd1 vccd1 _17194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16145_ _17344_/CLK _16145_/D vssd1 vssd1 vccd1 vccd1 hold124/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13357_ hold5034/X _13856_/B _13356_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13357_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10569_ hold3428/X _10476_/A _10568_/X vssd1 vssd1 vccd1 vccd1 _10569_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12308_ _17260_/Q _12308_/B _13721_/S vssd1 vssd1 vccd1 vccd1 _12308_/X sky130_fd_sc_hd__and3_1
X_16076_ _17284_/CLK _16076_/D vssd1 vssd1 vccd1 vccd1 hold466/A sky130_fd_sc_hd__dfxtp_1
X_13288_ _13281_/X _13287_/X _13296_/B1 vssd1 vssd1 vccd1 vccd1 _17554_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_228_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15027_ _14850_/A hold2856/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15028_/B sky130_fd_sc_hd__mux2_1
X_12239_ hold3116/X _17237_/Q _12335_/C vssd1 vssd1 vccd1 vccd1 _12240_/B sky130_fd_sc_hd__mux2_1
Xhold2609 _17903_/Q vssd1 vssd1 vccd1 vccd1 hold2609/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1908 _14957_/X vssd1 vssd1 vccd1 vccd1 _18265_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1919 _18170_/Q vssd1 vssd1 vccd1 vccd1 hold1919/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07780_ hold235/X vssd1 vssd1 vccd1 vccd1 _07780_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_235_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16978_ _17858_/CLK _16978_/D vssd1 vssd1 vccd1 vccd1 _16978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput4 input4/A vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15929_ _16124_/CLK _15929_/D vssd1 vssd1 vccd1 vccd1 hold777/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09450_ _09456_/C _09456_/D _09478_/B vssd1 vssd1 vccd1 vccd1 _09450_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_204_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08401_ _15515_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08401_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09381_ hold513/X _09386_/A _09362_/C hold440/X vssd1 vssd1 vccd1 vccd1 _09381_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_203_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08332_ hold1515/X _08323_/B _08331_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _08332_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08263_ hold2893/X _08262_/B _08262_/Y _08385_/A vssd1 vssd1 vccd1 vccd1 _08263_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08194_ hold2758/X _08213_/B _08193_/X _13765_/C1 vssd1 vssd1 vccd1 vccd1 _08194_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5202 _10915_/X vssd1 vssd1 vccd1 vccd1 _16795_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5213 _16952_/Q vssd1 vssd1 vccd1 vccd1 hold5213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5224 _12148_/X vssd1 vssd1 vccd1 vccd1 _17206_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5235 _16976_/Q vssd1 vssd1 vccd1 vccd1 hold5235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4501 _16626_/Q vssd1 vssd1 vccd1 vccd1 hold4501/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5246 _11086_/X vssd1 vssd1 vccd1 vccd1 _16852_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4512 _16372_/Q vssd1 vssd1 vccd1 vccd1 hold4512/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5257 _17054_/Q vssd1 vssd1 vccd1 vccd1 hold5257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5268 _10801_/X vssd1 vssd1 vccd1 vccd1 _16757_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4523 _17355_/Q vssd1 vssd1 vccd1 vccd1 hold4523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4534 _17358_/Q vssd1 vssd1 vccd1 vccd1 hold4534/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5279 _16797_/Q vssd1 vssd1 vccd1 vccd1 hold5279/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3800 _10153_/X vssd1 vssd1 vccd1 vccd1 _16541_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4545 _16404_/Q vssd1 vssd1 vccd1 vccd1 hold4545/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3811 _16565_/Q vssd1 vssd1 vccd1 vccd1 hold3811/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4556 _10228_/X vssd1 vssd1 vccd1 vccd1 _16566_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4567 _16429_/Q vssd1 vssd1 vccd1 vccd1 hold4567/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3822 _16478_/Q vssd1 vssd1 vccd1 vccd1 hold3822/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3833 _10501_/X vssd1 vssd1 vccd1 vccd1 _16657_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4578 _10354_/X vssd1 vssd1 vccd1 vccd1 _16608_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3844 _16763_/Q vssd1 vssd1 vccd1 vccd1 hold3844/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4589 _17695_/Q vssd1 vssd1 vccd1 vccd1 hold4589/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3855 _11842_/X vssd1 vssd1 vccd1 vccd1 _17104_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3866 _17058_/Q vssd1 vssd1 vccd1 vccd1 hold3866/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3877 _10180_/X vssd1 vssd1 vccd1 vccd1 _16550_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3888 _17645_/Q vssd1 vssd1 vccd1 vccd1 hold3888/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3899 _16595_/Q vssd1 vssd1 vccd1 vccd1 hold3899/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07978_ _15547_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _07978_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09717_ _09933_/A _09717_/B vssd1 vssd1 vccd1 vccd1 _09717_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09648_ _09948_/A _09648_/B vssd1 vssd1 vccd1 vccd1 _09648_/X sky130_fd_sc_hd__or2_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_237_wb_clk_i clkbuf_6_62_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18213_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09579_ _10539_/A _09579_/B vssd1 vssd1 vccd1 vccd1 _09579_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _12240_/A _11610_/B vssd1 vssd1 vccd1 vccd1 _11610_/X sky130_fd_sc_hd__or2_1
XFILLER_0_194_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12590_ hold3295/X _12589_/X _12923_/S vssd1 vssd1 vccd1 vccd1 _12591_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_148_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11541_ _11637_/A _11541_/B vssd1 vssd1 vccd1 vccd1 _11541_/X sky130_fd_sc_hd__or2_1
XFILLER_0_147_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14260_ _14529_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14260_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ _11670_/A _11472_/B vssd1 vssd1 vccd1 vccd1 _11472_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13211_ _13210_/X _16919_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13211_/X sky130_fd_sc_hd__mux2_1
X_10423_ hold3298/X _10631_/B _10422_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10423_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14191_ hold1611/X _14202_/B _14190_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _14191_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13142_ _13142_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13142_/X sky130_fd_sc_hd__or2_1
X_10354_ hold4577/X _10646_/B _10353_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _10354_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13073_ _13073_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13073_/X sky130_fd_sc_hd__and2_1
X_17950_ _18072_/CLK _17950_/D vssd1 vssd1 vccd1 vccd1 _17950_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5780 _13714_/X vssd1 vssd1 vccd1 vccd1 _17691_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10285_ hold3608/X _10571_/B _10284_/X _14769_/C1 vssd1 vssd1 vccd1 vccd1 _10285_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5791 _17178_/Q vssd1 vssd1 vccd1 vccd1 hold5791/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12024_ _12216_/A _12024_/B vssd1 vssd1 vccd1 vccd1 _12024_/X sky130_fd_sc_hd__or2_1
X_16901_ _18427_/CLK _16901_/D vssd1 vssd1 vccd1 vccd1 _16901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17881_ _17881_/CLK _17881_/D vssd1 vssd1 vccd1 vccd1 _17881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16832_ _18067_/CLK _16832_/D vssd1 vssd1 vccd1 vccd1 _16832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_217_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_219_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout590 _13049_/Y vssd1 vssd1 vccd1 vccd1 _13311_/C1 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_205_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16763_ _18030_/CLK _16763_/D vssd1 vssd1 vccd1 vccd1 _16763_/Q sky130_fd_sc_hd__dfxtp_1
X_13975_ hold1440/X _13995_/A2 _13974_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _13975_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15714_ _17617_/CLK _15714_/D vssd1 vssd1 vccd1 vccd1 _15714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12926_ hold4530/X _12925_/X _12929_/S vssd1 vssd1 vccd1 vccd1 _12927_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_198_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16694_ _18156_/CLK _16694_/D vssd1 vssd1 vccd1 vccd1 _16694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18433_ _18437_/CLK _18433_/D vssd1 vssd1 vccd1 vccd1 _18433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15645_ _17157_/CLK _15645_/D vssd1 vssd1 vccd1 vccd1 _15645_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ hold3318/X _12856_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12857_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_200_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18364_ _18396_/CLK _18364_/D vssd1 vssd1 vccd1 vccd1 _18364_/Q sky130_fd_sc_hd__dfxtp_1
X_11808_ _13800_/A _11808_/B vssd1 vssd1 vccd1 vccd1 _11808_/X sky130_fd_sc_hd__or2_1
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12788_ hold3396/X _12787_/X _12812_/S vssd1 vssd1 vccd1 vccd1 _12788_/X sky130_fd_sc_hd__mux2_1
X_15576_ _17244_/CLK _15576_/D vssd1 vssd1 vccd1 vccd1 _15576_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _17335_/CLK _17315_/D vssd1 vssd1 vccd1 vccd1 _17315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11739_ hold4417/X _11649_/A _11738_/X vssd1 vssd1 vccd1 vccd1 _11739_/Y sky130_fd_sc_hd__a21oi_1
X_14527_ _15207_/A _14543_/B vssd1 vssd1 vccd1 vccd1 _14527_/X sky130_fd_sc_hd__or2_1
X_18295_ _18389_/CLK _18295_/D vssd1 vssd1 vccd1 vccd1 _18295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17246_ _17278_/CLK _17246_/D vssd1 vssd1 vccd1 vccd1 _17246_/Q sky130_fd_sc_hd__dfxtp_1
X_14458_ hold2328/X _14487_/B _14457_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _14458_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13409_ hold1161/X hold4681/X _13409_/S vssd1 vssd1 vccd1 vccd1 _13410_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_142_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14389_ _15231_/A hold1169/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14390_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17177_ _17743_/CLK _17177_/D vssd1 vssd1 vccd1 vccd1 _17177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16128_ _17321_/CLK _16128_/D vssd1 vssd1 vccd1 vccd1 hold433/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08950_ _09440_/B hold883/X vssd1 vssd1 vccd1 vccd1 _16092_/D sky130_fd_sc_hd__and2_1
Xhold3107 _14689_/X vssd1 vssd1 vccd1 vccd1 _18136_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16059_ _16082_/CLK _16059_/D vssd1 vssd1 vccd1 vccd1 hold285/A sky130_fd_sc_hd__dfxtp_1
Xhold3118 _17374_/Q vssd1 vssd1 vccd1 vccd1 hold3118/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3129 _17751_/Q vssd1 vssd1 vccd1 vccd1 hold3129/X sky130_fd_sc_hd__dlygate4sd3_1
X_07901_ hold1082/X _07918_/B _07900_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _07901_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2406 _15768_/Q vssd1 vssd1 vccd1 vccd1 hold2406/X sky130_fd_sc_hd__dlygate4sd3_1
X_08881_ _09047_/A _08881_/B vssd1 vssd1 vccd1 vccd1 _16058_/D sky130_fd_sc_hd__and2_1
Xhold2417 _14771_/X vssd1 vssd1 vccd1 vccd1 _18176_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2428 _15695_/Q vssd1 vssd1 vccd1 vccd1 hold2428/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2439 _15579_/Q vssd1 vssd1 vccd1 vccd1 hold2439/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1705 _08424_/X vssd1 vssd1 vccd1 vccd1 _15842_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1716 _15666_/Q vssd1 vssd1 vccd1 vccd1 hold1716/X sky130_fd_sc_hd__dlygate4sd3_1
X_07832_ hold1887/X _07865_/B _07831_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _07832_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1727 _08104_/X vssd1 vssd1 vccd1 vccd1 _08105_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1738 _18457_/Q vssd1 vssd1 vccd1 vccd1 hold1738/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1749 _09109_/X vssd1 vssd1 vccd1 vccd1 _16169_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09502_ hold5030/X _09992_/B _09501_/X _15404_/A vssd1 vssd1 vccd1 vccd1 _09502_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_330_wb_clk_i clkbuf_6_44_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17906_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09433_ _07785_/Y _09477_/A _09440_/B hold705/X vssd1 vssd1 vccd1 vccd1 hold706/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09364_ _09366_/A _09364_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09364_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_164_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08315_ _15539_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08315_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_20 _13164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ _15517_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09295_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_1347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_31 _13212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_42 _17524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 hold220/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ _15525_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08246_/X sky130_fd_sc_hd__or2_1
XANTENNA_64 hold597/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_75 hold679/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_86 _15145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_97 hold5941/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08177_ hold915/X _08225_/B vssd1 vssd1 vccd1 vccd1 _08177_/X sky130_fd_sc_hd__or2_1
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5010 _16812_/Q vssd1 vssd1 vccd1 vccd1 hold5010/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5021 _11002_/X vssd1 vssd1 vccd1 vccd1 _16824_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5032 _17186_/Q vssd1 vssd1 vccd1 vccd1 hold5032/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5043 _10270_/X vssd1 vssd1 vccd1 vccd1 _16580_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5054 _17083_/Q vssd1 vssd1 vccd1 vccd1 hold5054/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5065 _10930_/X vssd1 vssd1 vccd1 vccd1 _16800_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4320 _17123_/Q vssd1 vssd1 vccd1 vccd1 hold4320/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4331 _10575_/Y vssd1 vssd1 vccd1 vccd1 _10576_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5076 _17253_/Q vssd1 vssd1 vccd1 vccd1 hold5076/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4342 _11178_/Y vssd1 vssd1 vccd1 vccd1 _11179_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5087 _11320_/X vssd1 vssd1 vccd1 vccd1 _16930_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5098 _12244_/X vssd1 vssd1 vccd1 vccd1 _17238_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4353 _16920_/Q vssd1 vssd1 vccd1 vccd1 hold4353/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4364 _16923_/Q vssd1 vssd1 vccd1 vccd1 hold4364/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3630 _16509_/Q vssd1 vssd1 vccd1 vccd1 hold3630/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4375 _12295_/Y vssd1 vssd1 vccd1 vccd1 _17255_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3641 _09715_/X vssd1 vssd1 vccd1 vccd1 _16395_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10070_ _16514_/Q _10070_/B _10985_/S vssd1 vssd1 vccd1 vccd1 _10070_/X sky130_fd_sc_hd__and3_1
Xhold4386 _11761_/Y vssd1 vssd1 vccd1 vccd1 _17077_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3652 _16477_/Q vssd1 vssd1 vccd1 vccd1 hold3652/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4397 _13887_/Y vssd1 vssd1 vccd1 vccd1 _13888_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3663 _09592_/X vssd1 vssd1 vccd1 vccd1 _16354_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3674 _16699_/Q vssd1 vssd1 vccd1 vccd1 hold3674/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2940 _18221_/Q vssd1 vssd1 vccd1 vccd1 hold2940/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3685 _10114_/X vssd1 vssd1 vccd1 vccd1 _16528_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2951 _15122_/X vssd1 vssd1 vccd1 vccd1 _18345_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3696 _17709_/Q vssd1 vssd1 vccd1 vccd1 hold3696/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2962 _18031_/Q vssd1 vssd1 vccd1 vccd1 hold2962/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2973 _18005_/Q vssd1 vssd1 vccd1 vccd1 hold2973/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_418_wb_clk_i clkbuf_6_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17260_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2984 _08455_/X vssd1 vssd1 vccd1 vccd1 _15856_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2995 _17934_/Q vssd1 vssd1 vccd1 vccd1 hold2995/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13760_ hold2790/X _17707_/Q _13871_/C vssd1 vssd1 vccd1 vccd1 _13761_/B sky130_fd_sc_hd__mux2_1
X_10972_ hold4727/X _11162_/B _10971_/X _14372_/A vssd1 vssd1 vccd1 vccd1 _10972_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12711_ _12786_/A _12711_/B vssd1 vssd1 vccd1 vccd1 _17413_/D sky130_fd_sc_hd__and2_1
XFILLER_0_74_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13691_ hold1793/X _17684_/Q _13883_/C vssd1 vssd1 vccd1 vccd1 _13692_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15430_ hold389/X _09365_/B _09362_/D hold327/X _15428_/X vssd1 vssd1 vccd1 vccd1
+ _15432_/C sky130_fd_sc_hd__a221o_1
X_12642_ _12849_/A _12642_/B vssd1 vssd1 vccd1 vccd1 _17390_/D sky130_fd_sc_hd__and2_1
XFILLER_0_195_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15361_ _16300_/Q _15477_/A2 _15487_/B1 _16088_/Q _15360_/X vssd1 vssd1 vccd1 vccd1
+ _15362_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_182_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12573_ _14358_/A _12573_/B vssd1 vssd1 vccd1 vccd1 _17367_/D sky130_fd_sc_hd__and2_1
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17100_ _17260_/CLK _17100_/D vssd1 vssd1 vccd1 vccd1 _17100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14312_ _15099_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14312_/X sky130_fd_sc_hd__or2_1
X_11524_ hold4119/X _12305_/B _11523_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _11524_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15292_ _15489_/A _15292_/B _15292_/C _15292_/D vssd1 vssd1 vccd1 vccd1 _15292_/X
+ sky130_fd_sc_hd__or4_1
X_18080_ _18106_/CLK _18080_/D vssd1 vssd1 vccd1 vccd1 _18080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17031_ _17847_/CLK _17031_/D vssd1 vssd1 vccd1 vccd1 _17031_/Q sky130_fd_sc_hd__dfxtp_1
X_14243_ hold2635/X _14268_/B _14242_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _14243_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11455_ hold5307/X _11741_/B _11454_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _11455_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_1295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10406_ hold1692/X hold4501/X _11213_/C vssd1 vssd1 vccd1 vccd1 _10407_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14174_ _15193_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14174_/X sky130_fd_sc_hd__or2_1
X_11386_ hold4783/X _11798_/B _11385_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _11386_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13125_ _13124_/X hold3435/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13125_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10337_ hold2135/X _16603_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10338_/B sky130_fd_sc_hd__mux2_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _17523_/Q _17522_/Q _13056_/C _13056_/D vssd1 vssd1 vccd1 vccd1 _13267_/S
+ sky130_fd_sc_hd__and4b_4
XFILLER_0_178_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17933_ _17973_/CLK _17933_/D vssd1 vssd1 vccd1 vccd1 _17933_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10268_ hold2685/X hold3654/X _11186_/C vssd1 vssd1 vccd1 vccd1 _10269_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_218_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12007_ hold4793/X _13811_/B _12006_/X _08363_/A vssd1 vssd1 vccd1 vccd1 _12007_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_218_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17864_ _17936_/CLK _17864_/D vssd1 vssd1 vccd1 vccd1 _17864_/Q sky130_fd_sc_hd__dfxtp_1
X_10199_ hold3097/X hold3692/X _10595_/C vssd1 vssd1 vccd1 vccd1 _10200_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_178_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_159_wb_clk_i clkbuf_6_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17299_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16815_ _18050_/CLK _16815_/D vssd1 vssd1 vccd1 vccd1 _16815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17795_ _18065_/CLK _17795_/D vssd1 vssd1 vccd1 vccd1 _17795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16746_ _18045_/CLK _16746_/D vssd1 vssd1 vccd1 vccd1 _16746_/Q sky130_fd_sc_hd__dfxtp_1
X_13958_ _15519_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13958_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12909_ _12924_/A _12909_/B vssd1 vssd1 vccd1 vccd1 _17479_/D sky130_fd_sc_hd__and2_1
X_16677_ _18235_/CLK _16677_/D vssd1 vssd1 vccd1 vccd1 _16677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13889_ _07786_/Y _16286_/Q hold901/X _10964_/S vssd1 vssd1 vccd1 vccd1 _13889_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_201_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_235_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18416_ _18416_/CLK _18416_/D vssd1 vssd1 vccd1 vccd1 _18416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15628_ _17724_/CLK _15628_/D vssd1 vssd1 vccd1 vccd1 _15628_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18347_ _18347_/CLK _18347_/D vssd1 vssd1 vccd1 vccd1 _18347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15559_ _15559_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15559_/X sky130_fd_sc_hd__or2_1
X_08100_ _14732_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08100_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09080_ _14980_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09080_/X sky130_fd_sc_hd__or2_1
X_18278_ _18382_/CLK _18278_/D vssd1 vssd1 vccd1 vccd1 _18278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08031_ _15545_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _08031_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_163_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput40 input40/A vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_1
X_17229_ _17229_/CLK _17229_/D vssd1 vssd1 vccd1 vccd1 _17229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput51 input51/A vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_1
Xhold802 hold802/A vssd1 vssd1 vccd1 vccd1 hold802/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput62 input62/A vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_1
Xhold813 hold813/A vssd1 vssd1 vccd1 vccd1 hold813/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 hold824/A vssd1 vssd1 vccd1 vccd1 hold824/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 hold835/A vssd1 vssd1 vccd1 vccd1 hold835/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 hold846/A vssd1 vssd1 vccd1 vccd1 hold846/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold857 hold857/A vssd1 vssd1 vccd1 vccd1 hold857/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold868 hold868/A vssd1 vssd1 vccd1 vccd1 hold868/X sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ _13062_/A _10022_/B _09981_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _09982_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_204_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold879 hold879/A vssd1 vssd1 vccd1 vccd1 hold879/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08933_ _15284_/A hold650/X vssd1 vssd1 vccd1 vccd1 _16084_/D sky130_fd_sc_hd__and2_1
XFILLER_0_149_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2203 _15589_/Q vssd1 vssd1 vccd1 vccd1 hold2203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2214 _15186_/X vssd1 vssd1 vccd1 vccd1 _18375_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2225 la_data_in[8] vssd1 vssd1 vccd1 vccd1 hold2225/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2236 _18167_/Q vssd1 vssd1 vccd1 vccd1 hold2236/X sky130_fd_sc_hd__dlygate4sd3_1
X_08864_ hold320/X hold401/X _08866_/S vssd1 vssd1 vccd1 vccd1 _08865_/B sky130_fd_sc_hd__mux2_1
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2247 _08467_/X vssd1 vssd1 vccd1 vccd1 _15862_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1502 _14315_/X vssd1 vssd1 vccd1 vccd1 _17957_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2258 _15092_/X vssd1 vssd1 vccd1 vccd1 _18330_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1513 _15685_/Q vssd1 vssd1 vccd1 vccd1 hold1513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2269 hold2269/A vssd1 vssd1 vccd1 vccd1 input69/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1524 _14472_/X vssd1 vssd1 vccd1 vccd1 _18033_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1535 _14187_/X vssd1 vssd1 vccd1 vccd1 _17896_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07815_ hold933/A _14980_/A _15519_/A _15517_/A vssd1 vssd1 vccd1 vccd1 _07817_/C
+ sky130_fd_sc_hd__or4_1
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1546 _15653_/Q vssd1 vssd1 vccd1 vccd1 hold1546/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08795_ _13056_/C hold935/X vssd1 vssd1 vccd1 vccd1 _13046_/D sky130_fd_sc_hd__nand2_1
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1557 _07915_/X vssd1 vssd1 vccd1 vccd1 _15601_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1568 _15773_/Q vssd1 vssd1 vccd1 vccd1 hold1568/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1579 hold1758/X vssd1 vssd1 vccd1 vccd1 hold1579/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09416_ _09438_/B _16294_/Q vssd1 vssd1 vccd1 vccd1 _09416_/X sky130_fd_sc_hd__or2_1
XFILLER_0_220_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09347_ _09366_/A _09363_/B _09351_/B vssd1 vssd1 vccd1 vccd1 _09347_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_118_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09278_ _12798_/A _09278_/B vssd1 vssd1 vccd1 vccd1 _16250_/D sky130_fd_sc_hd__and2_1
XFILLER_0_62_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08229_ _08504_/A _15128_/A vssd1 vssd1 vccd1 vccd1 _08260_/B sky130_fd_sc_hd__or2_4
XFILLER_0_106_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11240_ hold2217/X hold4674/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11241_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11171_ _16881_/Q _11171_/B _11171_/C vssd1 vssd1 vccd1 vccd1 _11171_/X sky130_fd_sc_hd__and3_1
XTAP_6301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4150 _11485_/X vssd1 vssd1 vccd1 vccd1 _16985_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10122_ _10482_/A _10122_/B vssd1 vssd1 vccd1 vccd1 _10122_/X sky130_fd_sc_hd__or2_1
Xhold4161 _16995_/Q vssd1 vssd1 vccd1 vccd1 hold4161/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4172 _09652_/X vssd1 vssd1 vccd1 vccd1 _16374_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4183 hold5973/X vssd1 vssd1 vccd1 vccd1 hold5974/A sky130_fd_sc_hd__buf_6
XTAP_5600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4194 _15283_/X vssd1 vssd1 vccd1 vccd1 _15284_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3460 _10641_/Y vssd1 vssd1 vccd1 vccd1 _10642_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14930_ _15199_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14930_/X sky130_fd_sc_hd__or2_1
XTAP_5633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10053_ _13254_/A _09957_/A _10052_/X vssd1 vssd1 vccd1 vccd1 _10053_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3471 _12309_/Y vssd1 vssd1 vccd1 vccd1 _12310_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3482 _10590_/Y vssd1 vssd1 vccd1 vccd1 _10591_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3493 _17583_/Q vssd1 vssd1 vccd1 vccd1 hold3493/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_252_wb_clk_i clkbuf_6_59_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18232_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2770 _09089_/X vssd1 vssd1 vccd1 vccd1 _16159_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14861_ hold2261/X _14880_/B _14860_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _14861_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2781 _18058_/Q vssd1 vssd1 vccd1 vccd1 hold2781/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2792 _15603_/Q vssd1 vssd1 vccd1 vccd1 hold2792/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16600_ _18194_/CLK _16600_/D vssd1 vssd1 vccd1 vccd1 _16600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13812_ hold4270/X _13716_/A _13811_/X vssd1 vssd1 vccd1 vccd1 _13812_/Y sky130_fd_sc_hd__a21oi_1
X_17580_ _17740_/CLK _17580_/D vssd1 vssd1 vccd1 vccd1 _17580_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14792_ _15185_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14792_/X sky130_fd_sc_hd__or2_1
XFILLER_0_203_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16531_ _18177_/CLK _16531_/D vssd1 vssd1 vccd1 vccd1 _16531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10955_ hold3031/X hold4053/X _11153_/C vssd1 vssd1 vccd1 vccd1 _10956_/B sky130_fd_sc_hd__mux2_1
X_13743_ _13773_/A _13743_/B vssd1 vssd1 vccd1 vccd1 _13743_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16462_ _18375_/CLK _16462_/D vssd1 vssd1 vccd1 vccd1 _16462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13674_ _13794_/A _13674_/B vssd1 vssd1 vccd1 vccd1 _13674_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10886_ _17989_/Q hold4059/X _11753_/C vssd1 vssd1 vccd1 vccd1 _10887_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18201_ _18224_/CLK _18201_/D vssd1 vssd1 vccd1 vccd1 _18201_/Q sky130_fd_sc_hd__dfxtp_1
X_15413_ _15490_/A1 _15405_/X _15412_/X _15490_/B1 hold5967/A vssd1 vssd1 vccd1 vccd1
+ _15413_/X sky130_fd_sc_hd__a32o_1
XPHY_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12625_ _18437_/Q _17386_/Q _12850_/S vssd1 vssd1 vccd1 vccd1 _12625_/X sky130_fd_sc_hd__mux2_1
XPHY_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16393_ _18370_/CLK _16393_/D vssd1 vssd1 vccd1 vccd1 _16393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18132_ _18236_/CLK _18132_/D vssd1 vssd1 vccd1 vccd1 _18132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15344_ _15344_/A _15344_/B vssd1 vssd1 vccd1 vccd1 _18410_/D sky130_fd_sc_hd__and2_1
X_12556_ hold1149/X _17363_/Q _12985_/S vssd1 vssd1 vccd1 vccd1 _12556_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11507_ hold2244/X hold4089/X _12173_/S vssd1 vssd1 vccd1 vccd1 _11508_/B sky130_fd_sc_hd__mux2_1
X_18063_ _18063_/CLK _18063_/D vssd1 vssd1 vccd1 vccd1 _18063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12487_ hold5/X _12445_/A _12445_/B _12486_/X _09057_/A vssd1 vssd1 vccd1 vccd1 hold6/A
+ sky130_fd_sc_hd__o311a_1
X_15275_ hold479/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15275_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold109 hold109/A vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
X_17014_ _17862_/CLK _17014_/D vssd1 vssd1 vccd1 vccd1 _17014_/Q sky130_fd_sc_hd__dfxtp_1
X_14226_ hold945/X _14230_/B vssd1 vssd1 vccd1 vccd1 _14226_/X sky130_fd_sc_hd__or2_1
X_11438_ hold1911/X _16970_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _11439_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_227_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14157_ hold884/X _14148_/B _14156_/X _12660_/A vssd1 vssd1 vccd1 vccd1 hold885/A
+ sky130_fd_sc_hd__o211a_1
X_11369_ hold1783/X _16947_/Q _11753_/C vssd1 vssd1 vccd1 vccd1 _11370_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13108_ hold4469/X _13107_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13108_/X sky130_fd_sc_hd__mux2_2
X_14088_ _15541_/A _14094_/B vssd1 vssd1 vccd1 vccd1 _14088_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_237_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_237_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13039_ hold905/X _13039_/B vssd1 vssd1 vccd1 vccd1 hold906/A sky130_fd_sc_hd__and2_1
XFILLER_0_185_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17916_ _18046_/CLK _17916_/D vssd1 vssd1 vccd1 vccd1 _17916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17847_ _17847_/CLK _17847_/D vssd1 vssd1 vccd1 vccd1 _17847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_233_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08580_ hold143/X hold785/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08581_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17778_ _17905_/CLK _17778_/D vssd1 vssd1 vccd1 vccd1 _17778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16729_ _18060_/CLK _16729_/D vssd1 vssd1 vccd1 vccd1 _16729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09201_ hold2747/X _09214_/B _09200_/X _12804_/A vssd1 vssd1 vccd1 vccd1 _09201_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_56_wb_clk_i clkbuf_6_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18307_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_174_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09132_ _15515_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09132_/X sky130_fd_sc_hd__or2_1
XFILLER_0_174_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09063_ _12420_/A hold388/X vssd1 vssd1 vccd1 vccd1 _16148_/D sky130_fd_sc_hd__and2_1
XFILLER_0_163_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08014_ hold1229/X _08029_/B _08013_/X _08363_/A vssd1 vssd1 vccd1 vccd1 _08014_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold610 hold610/A vssd1 vssd1 vccd1 vccd1 hold610/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold621 hold621/A vssd1 vssd1 vccd1 vccd1 hold621/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold632 hold632/A vssd1 vssd1 vccd1 vccd1 hold632/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 hold643/A vssd1 vssd1 vccd1 vccd1 hold643/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold654 hold654/A vssd1 vssd1 vccd1 vccd1 hold654/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold665 hold665/A vssd1 vssd1 vccd1 vccd1 hold665/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold676 data_in[7] vssd1 vssd1 vccd1 vccd1 hold676/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold687 hold687/A vssd1 vssd1 vccd1 vccd1 hold687/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold698 hold698/A vssd1 vssd1 vccd1 vccd1 hold698/X sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ hold1165/X _16479_/Q _10601_/C vssd1 vssd1 vccd1 vccd1 _09966_/B sky130_fd_sc_hd__mux2_1
Xhold2000 _18453_/Q vssd1 vssd1 vccd1 vccd1 hold2000/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2011 _15791_/Q vssd1 vssd1 vccd1 vccd1 hold2011/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2022 _14713_/X vssd1 vssd1 vccd1 vccd1 _18148_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2033 _18159_/Q vssd1 vssd1 vccd1 vccd1 hold2033/X sky130_fd_sc_hd__dlygate4sd3_1
X_08916_ hold92/X hold466/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold467/A sky130_fd_sc_hd__mux2_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2044 _08396_/X vssd1 vssd1 vccd1 vccd1 _15828_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09896_ _18369_/Q hold4725/X _09992_/C vssd1 vssd1 vccd1 vccd1 _09897_/B sky130_fd_sc_hd__mux2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2055 _17756_/Q vssd1 vssd1 vccd1 vccd1 hold2055/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1310 _09336_/X vssd1 vssd1 vccd1 vccd1 _16278_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2066 _18023_/Q vssd1 vssd1 vccd1 vccd1 hold2066/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1321 _17892_/Q vssd1 vssd1 vccd1 vccd1 hold1321/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1332 _15797_/Q vssd1 vssd1 vccd1 vccd1 hold1332/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2077 _15665_/Q vssd1 vssd1 vccd1 vccd1 hold2077/X sky130_fd_sc_hd__dlygate4sd3_1
X_08847_ _12418_/A _08847_/B vssd1 vssd1 vccd1 vccd1 _16042_/D sky130_fd_sc_hd__and2_1
Xhold2088 _17933_/Q vssd1 vssd1 vccd1 vccd1 hold2088/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1343 _14444_/X vssd1 vssd1 vccd1 vccd1 _18020_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1354 _15637_/Q vssd1 vssd1 vccd1 vccd1 hold1354/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2099 _14438_/X vssd1 vssd1 vccd1 vccd1 _18017_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1365 hold909/X vssd1 vssd1 vccd1 vccd1 input59/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1376 _15885_/Q vssd1 vssd1 vccd1 vccd1 hold1376/X sky130_fd_sc_hd__dlygate4sd3_1
X_08778_ _15404_/A hold612/X vssd1 vssd1 vccd1 vccd1 _16009_/D sky130_fd_sc_hd__and2_1
Xhold1387 _09087_/X vssd1 vssd1 vccd1 vccd1 _16158_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1398 _08204_/X vssd1 vssd1 vccd1 vccd1 _15738_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10740_ _11124_/A _10740_/B vssd1 vssd1 vccd1 vccd1 _10740_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10671_ _11043_/A _10671_/B vssd1 vssd1 vccd1 vccd1 _10671_/X sky130_fd_sc_hd__or2_1
XFILLER_0_211_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ _12410_/A _12410_/B vssd1 vssd1 vccd1 vccd1 _17298_/D sky130_fd_sc_hd__and2_1
XFILLER_0_153_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13390_ hold5739/X _13847_/B _13389_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13390_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12341_ _12341_/A _13886_/B _13886_/C vssd1 vssd1 vccd1 vccd1 _12341_/X sky130_fd_sc_hd__and3_1
XFILLER_0_180_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15060_ _15060_/A hold236/X vssd1 vssd1 vccd1 vccd1 hold237/A sky130_fd_sc_hd__and2_1
XFILLER_0_133_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12272_ hold2402/X _17248_/Q _13886_/C vssd1 vssd1 vccd1 vccd1 _12273_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_105_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14011_ hold2597/X _14040_/B _14010_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _14011_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11223_ hold4414/X _11127_/A _11222_/X vssd1 vssd1 vccd1 vccd1 _11223_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_433_wb_clk_i clkbuf_6_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17630_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11154_ hold4259/X _11136_/A _11153_/X vssd1 vssd1 vccd1 vccd1 _11154_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10105_ hold3692/X _10625_/B _10104_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _10105_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15962_ _17324_/CLK _15962_/D vssd1 vssd1 vccd1 vccd1 hold865/A sky130_fd_sc_hd__dfxtp_1
XTAP_5430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11085_ _11109_/A _11085_/B vssd1 vssd1 vccd1 vccd1 _11085_/X sky130_fd_sc_hd__or2_1
XTAP_5441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17701_ _17707_/CLK _17701_/D vssd1 vssd1 vccd1 vccd1 _17701_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3290 _17375_/Q vssd1 vssd1 vccd1 vccd1 hold3290/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10036_ _11206_/A _10036_/B vssd1 vssd1 vccd1 vccd1 _16502_/D sky130_fd_sc_hd__nor2_1
X_14913_ hold406/X _15182_/B vssd1 vssd1 vccd1 vccd1 hold407/A sky130_fd_sc_hd__or2_1
XTAP_5474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15893_ _17339_/CLK _15893_/D vssd1 vssd1 vccd1 vccd1 hold815/A sky130_fd_sc_hd__dfxtp_1
XTAP_5485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17632_ _17728_/CLK _17632_/D vssd1 vssd1 vccd1 vccd1 _17632_/Q sky130_fd_sc_hd__dfxtp_1
X_14844_ _15183_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14844_/X sky130_fd_sc_hd__or2_1
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17563_ _17721_/CLK _17563_/D vssd1 vssd1 vccd1 vccd1 _17563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14775_ hold1033/X _14774_/B _14774_/Y _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14775_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11987_ hold1966/X hold4072/X _13748_/S vssd1 vssd1 vccd1 vccd1 _11988_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_105_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16514_ _18395_/CLK _16514_/D vssd1 vssd1 vccd1 vccd1 _16514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13726_ hold4612/X _13829_/B _13725_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13726_/X
+ sky130_fd_sc_hd__o211a_1
X_17494_ _17513_/CLK _17494_/D vssd1 vssd1 vccd1 vccd1 _17494_/Q sky130_fd_sc_hd__dfxtp_1
X_10938_ _11124_/A _10938_/B vssd1 vssd1 vccd1 vccd1 _10938_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16445_ _18388_/CLK _16445_/D vssd1 vssd1 vccd1 vccd1 _16445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10869_ _11136_/A _10869_/B vssd1 vssd1 vccd1 vccd1 _10869_/X sky130_fd_sc_hd__or2_1
X_13657_ hold5233/X _13868_/B _13656_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13657_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12608_ hold3263/X _12607_/X _12923_/S vssd1 vssd1 vccd1 vccd1 _12608_/X sky130_fd_sc_hd__mux2_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _18321_/CLK _16376_/D vssd1 vssd1 vccd1 vccd1 _16376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13588_ hold5460/X _13874_/B _13587_/X _13684_/C1 vssd1 vssd1 vccd1 vccd1 _13588_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18115_ _18115_/CLK _18115_/D vssd1 vssd1 vccd1 vccd1 _18115_/Q sky130_fd_sc_hd__dfxtp_1
X_15327_ _16141_/Q _15487_/A2 _15484_/B1 _15890_/Q _15326_/X vssd1 vssd1 vccd1 vccd1
+ _15332_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_14_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12539_ hold4536/X _12538_/X _12929_/S vssd1 vssd1 vccd1 vccd1 _12540_/B sky130_fd_sc_hd__mux2_1
Xhold5609 _13660_/X vssd1 vssd1 vccd1 vccd1 _17673_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18046_ _18046_/CLK _18046_/D vssd1 vssd1 vccd1 vccd1 _18046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15258_ hold472/X _15484_/A2 _09392_/D hold390/X vssd1 vssd1 vccd1 vccd1 _15258_/X
+ sky130_fd_sc_hd__a22o_1
Xhold4908 _10726_/X vssd1 vssd1 vccd1 vccd1 _16732_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4919 _16408_/Q vssd1 vssd1 vccd1 vccd1 hold4919/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14209_ hold3035/X _14202_/B _14208_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _14209_/X
+ sky130_fd_sc_hd__o211a_1
X_15189_ _15189_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15189_/X sky130_fd_sc_hd__or2_1
XFILLER_0_240_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_174_wb_clk_i clkbuf_6_48_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18385_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout408 _14286_/Y vssd1 vssd1 vccd1 vccd1 _14326_/B sky130_fd_sc_hd__clkbuf_8
Xfanout419 _14107_/A2 vssd1 vssd1 vccd1 vccd1 _14094_/B sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_103_wb_clk_i clkbuf_6_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17301_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_225_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09750_ _09954_/A _09750_/B vssd1 vssd1 vccd1 vccd1 _09750_/X sky130_fd_sc_hd__or2_1
XFILLER_0_225_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08701_ hold245/X hold846/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08702_/B sky130_fd_sc_hd__mux2_1
X_09681_ _09978_/A _09681_/B vssd1 vssd1 vccd1 vccd1 _09681_/X sky130_fd_sc_hd__or2_1
XFILLER_0_207_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08632_ _12438_/A hold186/X vssd1 vssd1 vccd1 vccd1 _15938_/D sky130_fd_sc_hd__and2_1
XFILLER_0_234_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08563_ _12426_/A hold543/X vssd1 vssd1 vccd1 vccd1 _15905_/D sky130_fd_sc_hd__and2_1
XFILLER_0_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_234_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08494_ _14726_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08494_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09115_ hold2031/X _09106_/B _09114_/X _15244_/A vssd1 vssd1 vccd1 vccd1 _09115_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_6_20_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_20_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09046_ hold92/X hold138/X _09056_/S vssd1 vssd1 vccd1 vccd1 hold139/A sky130_fd_sc_hd__mux2_1
XFILLER_0_142_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold440 hold440/A vssd1 vssd1 vccd1 vccd1 hold440/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 input35/X vssd1 vssd1 vccd1 vccd1 hold451/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 hold462/A vssd1 vssd1 vccd1 vccd1 hold462/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 hold473/A vssd1 vssd1 vccd1 vccd1 hold473/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 hold484/A vssd1 vssd1 vccd1 vccd1 hold484/X sky130_fd_sc_hd__buf_8
XFILLER_0_25_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold495 hold56/X vssd1 vssd1 vccd1 vccd1 hold495/X sky130_fd_sc_hd__buf_4
XFILLER_0_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout920 hold484/X vssd1 vssd1 vccd1 vccd1 _15549_/A sky130_fd_sc_hd__buf_12
Xfanout931 hold630/X vssd1 vssd1 vccd1 vccd1 _14477_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_217_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09948_ _09948_/A _09948_/B vssd1 vssd1 vccd1 vccd1 _09948_/X sky130_fd_sc_hd__or2_1
Xfanout942 _15203_/A vssd1 vssd1 vccd1 vccd1 _15529_/A sky130_fd_sc_hd__buf_12
XFILLER_0_102_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ _10986_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09879_/X sky130_fd_sc_hd__or2_1
Xhold1140 _15174_/X vssd1 vssd1 vccd1 vccd1 _18370_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1151 la_data_in[10] vssd1 vssd1 vccd1 vccd1 hold1151/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1162 _08501_/X vssd1 vssd1 vccd1 vccd1 _15879_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ _12198_/A _11910_/B vssd1 vssd1 vccd1 vccd1 _11910_/X sky130_fd_sc_hd__or2_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1173 _15660_/Q vssd1 vssd1 vccd1 vccd1 hold1173/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ hold3147/X _12889_/X _12905_/S vssd1 vssd1 vccd1 vccd1 _12890_/X sky130_fd_sc_hd__mux2_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 _15535_/A vssd1 vssd1 vccd1 vccd1 _09313_/A sky130_fd_sc_hd__buf_8
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1195 _09181_/X vssd1 vssd1 vccd1 vccd1 _16202_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11841_ _13314_/A _11841_/B vssd1 vssd1 vccd1 vccd1 _11841_/X sky130_fd_sc_hd__or2_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ _15492_/A _14573_/B _18075_/Q vssd1 vssd1 vccd1 vccd1 _14560_/X sky130_fd_sc_hd__a21o_1
X_11772_ hold4717/X _12243_/A _11771_/X vssd1 vssd1 vccd1 vccd1 _11772_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ hold3844/X _11171_/B _10722_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _10723_/X
+ sky130_fd_sc_hd__o211a_1
X_13511_ hold1098/X _17624_/Q _13817_/C vssd1 vssd1 vccd1 vccd1 _13512_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14491_ hold992/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14491_/X sky130_fd_sc_hd__or2_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16230_ _17434_/CLK _16230_/D vssd1 vssd1 vccd1 vccd1 _16230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10654_ hold3978/X _11723_/B _10653_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _10654_/X
+ sky130_fd_sc_hd__o211a_1
X_13442_ hold2591/X _17601_/Q _13862_/C vssd1 vssd1 vccd1 vccd1 _13443_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_222_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16161_ _17499_/CLK _16161_/D vssd1 vssd1 vccd1 vccd1 _16161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13373_ hold1819/X hold4421/X _13874_/C vssd1 vssd1 vccd1 vccd1 _13374_/B sky130_fd_sc_hd__mux2_1
X_10585_ _10651_/A _10585_/B vssd1 vssd1 vccd1 vccd1 _16685_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15112_ hold2534/X hold341/X _15111_/Y _15062_/A vssd1 vssd1 vccd1 vccd1 _15112_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12324_ hold4438/X _12219_/A _12323_/X vssd1 vssd1 vccd1 vccd1 _12324_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16092_ _18408_/CLK _16092_/D vssd1 vssd1 vccd1 vccd1 hold882/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_1_wb_clk_i clkbuf_6_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17437_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15043_ _14596_/A hold1423/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15043_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12255_ _12255_/A _12255_/B vssd1 vssd1 vccd1 vccd1 _12255_/X sky130_fd_sc_hd__or2_1
XFILLER_0_239_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11206_ _11206_/A _11206_/B vssd1 vssd1 vccd1 vccd1 _16892_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12186_ _13407_/A _12186_/B vssd1 vssd1 vccd1 vccd1 _12186_/X sky130_fd_sc_hd__or2_1
X_11137_ hold4634/X _11153_/B _11136_/X _14552_/C1 vssd1 vssd1 vccd1 vccd1 _11137_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16994_ _17874_/CLK _16994_/D vssd1 vssd1 vccd1 vccd1 _16994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_236_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15945_ _18417_/CLK _15945_/D vssd1 vssd1 vccd1 vccd1 hold487/A sky130_fd_sc_hd__dfxtp_1
X_11068_ hold4869/X _11162_/B _11067_/X _14372_/A vssd1 vssd1 vccd1 vccd1 _11068_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10019_ _10019_/A _10028_/B _10028_/C vssd1 vssd1 vccd1 vccd1 _10019_/X sky130_fd_sc_hd__and3_1
XTAP_5293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_222_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15876_ _17747_/CLK _15876_/D vssd1 vssd1 vccd1 vccd1 _15876_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17615_ _17672_/CLK _17615_/D vssd1 vssd1 vccd1 vccd1 _17615_/Q sky130_fd_sc_hd__dfxtp_1
X_14827_ hold2528/X _14826_/B _14826_/Y _14893_/C1 vssd1 vssd1 vccd1 vccd1 _14827_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_231_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17546_ _18296_/CLK _17546_/D vssd1 vssd1 vccd1 vccd1 _17546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14758_ _15205_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14758_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13709_ hold1327/X hold5781/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13710_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_86_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17477_ _17477_/CLK _17477_/D vssd1 vssd1 vccd1 vccd1 _17477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14689_ hold3106/X _14720_/B _14688_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14689_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16428_ _18242_/CLK _16428_/D vssd1 vssd1 vccd1 vccd1 _16428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6107 _16307_/Q vssd1 vssd1 vccd1 vccd1 hold6107/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16359_ _18421_/CLK _16359_/D vssd1 vssd1 vccd1 vccd1 _16359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6118 data_in[28] vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6129 _09468_/X vssd1 vssd1 vccd1 vccd1 _09470_/C sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_355_wb_clk_i clkbuf_6_40_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17738_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5406 _17065_/Q vssd1 vssd1 vccd1 vccd1 hold5406/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5417 _13780_/X vssd1 vssd1 vccd1 vccd1 _17713_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5428 _17046_/Q vssd1 vssd1 vccd1 vccd1 hold5428/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5439 _13765_/X vssd1 vssd1 vccd1 vccd1 _17708_/D sky130_fd_sc_hd__dlygate4sd3_1
X_18029_ _18066_/CLK _18029_/D vssd1 vssd1 vccd1 vccd1 _18029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4705 _16833_/Q vssd1 vssd1 vccd1 vccd1 hold4705/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4716 _13522_/X vssd1 vssd1 vccd1 vccd1 _17627_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4727 _16846_/Q vssd1 vssd1 vccd1 vccd1 hold4727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4738 _13708_/X vssd1 vssd1 vccd1 vccd1 _17689_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4749 _17212_/Q vssd1 vssd1 vccd1 vccd1 hold4749/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout205 _11792_/B vssd1 vssd1 vccd1 vccd1 _11798_/B sky130_fd_sc_hd__buf_4
Xfanout216 _11201_/B vssd1 vssd1 vccd1 vccd1 _09992_/B sky130_fd_sc_hd__clkbuf_8
Xfanout227 _10634_/B vssd1 vssd1 vccd1 vccd1 _10052_/B sky130_fd_sc_hd__buf_4
X_09802_ hold4725/X _09992_/B _09801_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _09802_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout238 _10577_/B vssd1 vssd1 vccd1 vccd1 _10601_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout249 _13800_/A vssd1 vssd1 vccd1 vccd1 _13722_/A sky130_fd_sc_hd__buf_4
X_07994_ _08504_/A _09498_/A vssd1 vssd1 vccd1 vccd1 _08043_/B sky130_fd_sc_hd__or2_4
XFILLER_0_226_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09733_ hold3536/X _10046_/B _09732_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _09733_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09664_ hold3708/X _10046_/B _09663_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09664_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08615_ hold452/X _15930_/Q _08657_/S vssd1 vssd1 vccd1 vccd1 hold453/A sky130_fd_sc_hd__mux2_1
XFILLER_0_96_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09595_ hold3698/X _10601_/B _09594_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09595_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_1253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_wb_clk_i clkbuf_6_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17499_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08546_ hold679/X _15897_/Q _08592_/S vssd1 vssd1 vccd1 vccd1 hold680/A sky130_fd_sc_hd__mux2_1
XFILLER_0_194_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08477_ hold1819/X _08486_/B _08476_/X _13684_/C1 vssd1 vssd1 vccd1 vccd1 _08477_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10370_ hold2111/X _16614_/Q _10625_/C vssd1 vssd1 vccd1 vccd1 _10371_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_33_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09029_ _12420_/A _09029_/B vssd1 vssd1 vccd1 vccd1 _16131_/D sky130_fd_sc_hd__and2_1
XFILLER_0_142_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5940 _16281_/Q vssd1 vssd1 vccd1 vccd1 hold5940/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5951 _18418_/Q vssd1 vssd1 vccd1 vccd1 hold5951/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5962 _16284_/Q vssd1 vssd1 vccd1 vccd1 hold5962/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5973 _18425_/Q vssd1 vssd1 vccd1 vccd1 hold5973/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12040_ hold5805/X _12362_/B _12039_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _12040_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5984 _09472_/D vssd1 vssd1 vccd1 vccd1 _09465_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold270 hold364/X vssd1 vssd1 vccd1 vccd1 hold270/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5995 _17519_/Q vssd1 vssd1 vccd1 vccd1 _09490_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold281 hold281/A vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold292 hold292/A vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_218_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout750 _08119_/A vssd1 vssd1 vccd1 vccd1 _12265_/C1 sky130_fd_sc_hd__buf_4
Xfanout761 _14528_/C1 vssd1 vssd1 vccd1 vccd1 _13911_/A sky130_fd_sc_hd__buf_4
XFILLER_0_233_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout772 _08385_/A vssd1 vssd1 vccd1 vccd1 _08389_/A sky130_fd_sc_hd__buf_4
XFILLER_0_205_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout783 fanout791/X vssd1 vssd1 vccd1 vccd1 _14526_/C1 sky130_fd_sc_hd__buf_4
X_13991_ hold1809/X _13986_/B _13990_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _13991_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_232_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout794 fanout816/X vssd1 vssd1 vccd1 vccd1 _15056_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_204_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15730_ _17707_/CLK _15730_/D vssd1 vssd1 vccd1 vccd1 _15730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _12987_/A _12942_/B vssd1 vssd1 vccd1 vccd1 _17490_/D sky130_fd_sc_hd__and2_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _17779_/CLK _15661_/D vssd1 vssd1 vccd1 vccd1 _15661_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 _15219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _12873_/A _12873_/B vssd1 vssd1 vccd1 vccd1 _17467_/D sky130_fd_sc_hd__and2_1
XFILLER_0_241_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_121 _15173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17400_ _18438_/CLK _17400_/D vssd1 vssd1 vccd1 vccd1 _17400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14612_ _15221_/A _14612_/B vssd1 vssd1 vccd1 vccd1 _14612_/Y sky130_fd_sc_hd__nand2_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18380_ _18380_/CLK _18380_/D vssd1 vssd1 vccd1 vccd1 _18380_/Q sky130_fd_sc_hd__dfxtp_1
X_11824_ hold4835/X _13811_/B _11823_/X _12103_/C1 vssd1 vssd1 vccd1 vccd1 _11824_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _17272_/CLK hold979/X vssd1 vssd1 vccd1 vccd1 hold978/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_233_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17331_ _17331_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 _17331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _14543_/A _14543_/B vssd1 vssd1 vccd1 vccd1 _14543_/X sky130_fd_sc_hd__or2_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _12331_/A _11755_/B vssd1 vssd1 vccd1 vccd1 _11755_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_200_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10706_ hold1670/X hold4318/X _11186_/C vssd1 vssd1 vccd1 vccd1 _10707_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17262_ _17262_/CLK _17262_/D vssd1 vssd1 vccd1 vccd1 _17262_/Q sky130_fd_sc_hd__dfxtp_1
X_14474_ hold2666/X _14481_/B _14473_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14474_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11686_ hold5436/X _12323_/B _11685_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _11686_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16213_ _17723_/CLK _16213_/D vssd1 vssd1 vccd1 vccd1 _16213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13425_ _13719_/A _13425_/B vssd1 vssd1 vccd1 vccd1 _13425_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10637_ _16703_/Q _10637_/B _10637_/C vssd1 vssd1 vccd1 vccd1 _10637_/X sky130_fd_sc_hd__and3_1
XFILLER_0_154_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17193_ _18447_/CLK _17193_/D vssd1 vssd1 vccd1 vccd1 _17193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16144_ _17339_/CLK _16144_/D vssd1 vssd1 vccd1 vccd1 hold396/A sky130_fd_sc_hd__dfxtp_1
X_10568_ _16680_/Q _10568_/B _10571_/C vssd1 vssd1 vccd1 vccd1 _10568_/X sky130_fd_sc_hd__and3_1
XFILLER_0_148_1288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13356_ _13773_/A _13356_/B vssd1 vssd1 vccd1 vccd1 _13356_/X sky130_fd_sc_hd__or2_1
XFILLER_0_11_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12307_ _13819_/A _12307_/B vssd1 vssd1 vccd1 vccd1 _12307_/Y sky130_fd_sc_hd__nor2_1
X_16075_ _17338_/CLK _16075_/D vssd1 vssd1 vccd1 vccd1 _16075_/Q sky130_fd_sc_hd__dfxtp_1
X_10499_ hold2483/X hold3676/X _10595_/C vssd1 vssd1 vccd1 vccd1 _10500_/B sky130_fd_sc_hd__mux2_1
X_13287_ _13311_/A1 _13285_/X _13286_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13287_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15026_ _15026_/A _15026_/B vssd1 vssd1 vccd1 vccd1 _18298_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12238_ hold4583/X _12350_/B _12237_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _12238_/X
+ sky130_fd_sc_hd__o211a_1
X_12169_ hold5751/X _12362_/B _12168_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _12169_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1909 _16187_/Q vssd1 vssd1 vccd1 vccd1 hold1909/X sky130_fd_sc_hd__dlygate4sd3_1
X_16977_ _17825_/CLK _16977_/D vssd1 vssd1 vccd1 vccd1 _16977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput5 input5/A vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
X_15928_ _17347_/CLK _15928_/D vssd1 vssd1 vccd1 vccd1 hold207/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15859_ _17630_/CLK hold999/X vssd1 vssd1 vccd1 vccd1 hold998/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08400_ hold2987/X _08442_/A2 _08399_/X _12738_/A vssd1 vssd1 vccd1 vccd1 _08400_/X
+ sky130_fd_sc_hd__o211a_1
X_09380_ hold544/X _09365_/B _15477_/A2 vssd1 vssd1 vccd1 vccd1 _09383_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_59_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08331_ _15555_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08331_/X sky130_fd_sc_hd__or2_1
X_17529_ _17533_/CLK _17529_/D vssd1 vssd1 vccd1 vccd1 _17529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08262_ _15215_/A _08262_/B vssd1 vssd1 vccd1 vccd1 _08262_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08193_ _14413_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08193_/X sky130_fd_sc_hd__or2_1
XFILLER_0_172_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5203 _17733_/Q vssd1 vssd1 vccd1 vccd1 hold5203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5214 _11290_/X vssd1 vssd1 vccd1 vccd1 _16920_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5225 _16900_/Q vssd1 vssd1 vccd1 vccd1 hold5225/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5236 _11362_/X vssd1 vssd1 vccd1 vccd1 _16944_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4502 _10312_/X vssd1 vssd1 vccd1 vccd1 _16594_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5247 _16894_/Q vssd1 vssd1 vccd1 vccd1 hold5247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4513 _09550_/X vssd1 vssd1 vccd1 vccd1 _16340_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5258 _11596_/X vssd1 vssd1 vccd1 vccd1 _17022_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4524 _12536_/X vssd1 vssd1 vccd1 vccd1 _12537_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5269 _17028_/Q vssd1 vssd1 vccd1 vccd1 hold5269/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4535 _17489_/Q vssd1 vssd1 vccd1 vccd1 hold4535/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4546 _09646_/X vssd1 vssd1 vccd1 vccd1 _16372_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3801 _17741_/Q vssd1 vssd1 vccd1 vccd1 _13862_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3812 _10129_/X vssd1 vssd1 vccd1 vccd1 _16533_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4557 _16431_/Q vssd1 vssd1 vccd1 vccd1 hold4557/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4568 _09721_/X vssd1 vssd1 vccd1 vccd1 _16397_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3823 _09868_/X vssd1 vssd1 vccd1 vccd1 _16446_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3834 _16559_/Q vssd1 vssd1 vccd1 vccd1 hold3834/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4579 _16704_/Q vssd1 vssd1 vccd1 vccd1 hold4579/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3845 _10723_/X vssd1 vssd1 vccd1 vccd1 _16731_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3856 _17261_/Q vssd1 vssd1 vccd1 vccd1 _12311_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3867 _11608_/X vssd1 vssd1 vccd1 vccd1 _17026_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3878 _16670_/Q vssd1 vssd1 vccd1 vccd1 hold3878/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3889 _13480_/X vssd1 vssd1 vccd1 vccd1 _17613_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07977_ hold2618/X _07978_/B _07976_/Y _14147_/C1 vssd1 vssd1 vccd1 vccd1 _07977_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09716_ hold1262/X hold4463/X _10028_/C vssd1 vssd1 vccd1 vccd1 _09717_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_230_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09647_ hold1861/X hold3946/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09648_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_201_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09578_ hold1000/X _13270_/A _10040_/C vssd1 vssd1 vccd1 vccd1 _09579_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _12410_/A hold476/X vssd1 vssd1 vccd1 vccd1 _15889_/D sky130_fd_sc_hd__and2_1
XFILLER_0_194_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_277_wb_clk_i clkbuf_6_51_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18395_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11540_ hold2555/X hold5376/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11541_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_203_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_206_wb_clk_i clkbuf_6_55_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18081_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_147_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11471_ hold2967/X _16981_/Q _11765_/C vssd1 vssd1 vccd1 vccd1 _11472_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10422_ _10536_/A _10422_/B vssd1 vssd1 vccd1 vccd1 _10422_/X sky130_fd_sc_hd__or2_1
X_13210_ _17577_/Q _17111_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13210_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_135_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14190_ _14529_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14190_/X sky130_fd_sc_hd__or2_1
X_13141_ _13140_/X hold3486/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13141_/X sky130_fd_sc_hd__mux2_1
X_10353_ _10551_/A _10353_/B vssd1 vssd1 vccd1 vccd1 _10353_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13072_ _13065_/X _13071_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17527_/D sky130_fd_sc_hd__o21a_1
Xhold5770 _11860_/X vssd1 vssd1 vccd1 vccd1 _17110_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10284_ _10476_/A _10284_/B vssd1 vssd1 vccd1 vccd1 _10284_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5781 _17690_/Q vssd1 vssd1 vccd1 vccd1 hold5781/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5792 _11968_/X vssd1 vssd1 vccd1 vccd1 _17146_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12023_ hold1546/X hold4026/X _13481_/S vssd1 vssd1 vccd1 vccd1 _12024_/B sky130_fd_sc_hd__mux2_1
X_16900_ _18428_/CLK _16900_/D vssd1 vssd1 vccd1 vccd1 _16900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17880_ _18448_/CLK _17880_/D vssd1 vssd1 vccd1 vccd1 _17880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16831_ _18126_/CLK _16831_/D vssd1 vssd1 vccd1 vccd1 _16831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout580 _14163_/B vssd1 vssd1 vccd1 vccd1 _14502_/B sky130_fd_sc_hd__buf_6
Xfanout591 _12811_/S vssd1 vssd1 vccd1 vccd1 _12766_/S sky130_fd_sc_hd__buf_6
XFILLER_0_73_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16762_ _17997_/CLK _16762_/D vssd1 vssd1 vccd1 vccd1 _16762_/Q sky130_fd_sc_hd__dfxtp_1
X_13974_ _14529_/A _13994_/B vssd1 vssd1 vccd1 vccd1 _13974_/X sky130_fd_sc_hd__or2_1
X_15713_ _17153_/CLK _15713_/D vssd1 vssd1 vccd1 vccd1 _15713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12925_ hold1618/X hold4445/X _12925_/S vssd1 vssd1 vccd1 vccd1 _12925_/X sky130_fd_sc_hd__mux2_1
X_16693_ _18099_/CLK _16693_/D vssd1 vssd1 vccd1 vccd1 _16693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_214_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18432_ _18432_/CLK _18432_/D vssd1 vssd1 vccd1 vccd1 _18432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15644_ _17910_/CLK _15644_/D vssd1 vssd1 vccd1 vccd1 _15644_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12856_ hold2931/X _17463_/Q _12916_/S vssd1 vssd1 vccd1 vccd1 _12856_/X sky130_fd_sc_hd__mux2_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18363_ _18363_/CLK _18363_/D vssd1 vssd1 vccd1 vccd1 _18363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11807_ hold1451/X _17093_/Q _13796_/S vssd1 vssd1 vccd1 vccd1 _11808_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _17590_/CLK _15575_/D vssd1 vssd1 vccd1 vccd1 _15575_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12787_ hold2462/X _17440_/Q _12838_/S vssd1 vssd1 vccd1 vccd1 _12787_/X sky130_fd_sc_hd__mux2_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17314_ _17314_/CLK _17314_/D vssd1 vssd1 vccd1 vccd1 hold866/A sky130_fd_sc_hd__dfxtp_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14526_ hold1536/X _14541_/B _14525_/X _14526_/C1 vssd1 vssd1 vccd1 vccd1 _14526_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18294_ _18388_/CLK hold201/X vssd1 vssd1 vccd1 vccd1 _18294_/Q sky130_fd_sc_hd__dfxtp_1
X_11738_ _17070_/Q _11744_/B _11738_/C vssd1 vssd1 vccd1 vccd1 _11738_/X sky130_fd_sc_hd__and3_1
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17245_ _17277_/CLK _17245_/D vssd1 vssd1 vccd1 vccd1 _17245_/Q sky130_fd_sc_hd__dfxtp_1
X_14457_ _14457_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14457_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11669_ hold1273/X _17047_/Q _11765_/C vssd1 vssd1 vccd1 vccd1 _11670_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13408_ hold4981/X _13877_/B _13407_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _13408_/X
+ sky130_fd_sc_hd__o211a_1
X_17176_ _17272_/CLK _17176_/D vssd1 vssd1 vccd1 vccd1 _17176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14388_ _14388_/A _14388_/B vssd1 vssd1 vccd1 vccd1 _17993_/D sky130_fd_sc_hd__and2_1
XFILLER_0_141_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16127_ _16147_/CLK _16127_/D vssd1 vssd1 vccd1 vccd1 hold326/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13339_ hold4608/X _13829_/B _13338_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13339_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3108 _18382_/Q vssd1 vssd1 vccd1 vccd1 hold3108/X sky130_fd_sc_hd__dlygate4sd3_1
X_16058_ _16058_/CLK _16058_/D vssd1 vssd1 vccd1 vccd1 hold790/A sky130_fd_sc_hd__dfxtp_1
Xhold3119 _12593_/X vssd1 vssd1 vccd1 vccd1 _12594_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15009_ hold6059/X _15004_/B hold511/X _15146_/C1 vssd1 vssd1 vccd1 vccd1 hold512/A
+ sky130_fd_sc_hd__o211a_1
X_07900_ _14517_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07900_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2407 _08267_/X vssd1 vssd1 vccd1 vccd1 _15768_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08880_ hold147/X hold790/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08881_/B sky130_fd_sc_hd__mux2_1
Xhold2418 _17825_/Q vssd1 vssd1 vccd1 vccd1 hold2418/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2429 _17962_/Q vssd1 vssd1 vccd1 vccd1 hold2429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1706 _16254_/Q vssd1 vssd1 vccd1 vccd1 hold1706/X sky130_fd_sc_hd__dlygate4sd3_1
X_07831_ _15509_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07831_/X sky130_fd_sc_hd__or2_1
XFILLER_0_23_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1717 _08053_/X vssd1 vssd1 vccd1 vccd1 _15666_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1728 _18083_/Q vssd1 vssd1 vccd1 vccd1 hold1728/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1739 _15558_/X vssd1 vssd1 vccd1 vccd1 _18457_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_237_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09501_ _09987_/A _09501_/B vssd1 vssd1 vccd1 vccd1 _09501_/X sky130_fd_sc_hd__or2_1
XFILLER_0_155_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09432_ hold704/X _16302_/Q vssd1 vssd1 vccd1 vccd1 hold705/A sky130_fd_sc_hd__or2_1
XFILLER_0_172_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09363_ _09366_/A _09363_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09363_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_370_wb_clk_i clkbuf_6_34_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17739_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08314_ hold1585/X _08323_/B _08313_/X _12738_/A vssd1 vssd1 vccd1 vccd1 _08314_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09294_ hold2926/X _09325_/B _09293_/X _12612_/A vssd1 vssd1 vccd1 vccd1 _09294_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_10 _13116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _13164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_32 _13260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 _18419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08245_ hold1115/X _08262_/B _08244_/X _13765_/C1 vssd1 vssd1 vccd1 vccd1 _08245_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_54 hold220/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_65 hold597/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_76 hold915/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_87 _15145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_98 hold5947/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ hold1532/X _08209_/B _08175_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _08176_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5000 _16888_/Q vssd1 vssd1 vccd1 vccd1 hold5000/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5011 _10870_/X vssd1 vssd1 vccd1 vccd1 _16780_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5022 _17133_/Q vssd1 vssd1 vccd1 vccd1 hold5022/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5033 _11992_/X vssd1 vssd1 vccd1 vccd1 _17154_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5044 _16860_/Q vssd1 vssd1 vccd1 vccd1 hold5044/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5055 _11683_/X vssd1 vssd1 vccd1 vccd1 _17051_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4310 _11166_/Y vssd1 vssd1 vccd1 vccd1 _11167_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4321 _12378_/Y vssd1 vssd1 vccd1 vccd1 _12379_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5066 _16815_/Q vssd1 vssd1 vccd1 vccd1 hold5066/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4332 _17120_/Q vssd1 vssd1 vccd1 vccd1 hold4332/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5077 _12193_/X vssd1 vssd1 vccd1 vccd1 _17221_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5088 _16841_/Q vssd1 vssd1 vccd1 vccd1 hold5088/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4343 _17101_/Q vssd1 vssd1 vccd1 vccd1 hold4343/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5099 _17127_/Q vssd1 vssd1 vccd1 vccd1 hold5099/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4354 _11769_/Y vssd1 vssd1 vccd1 vccd1 _11770_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3620 _16369_/Q vssd1 vssd1 vccd1 vccd1 hold3620/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4365 _11778_/Y vssd1 vssd1 vccd1 vccd1 _11779_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3631 _09961_/X vssd1 vssd1 vccd1 vccd1 _16477_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4376 hold5930/X vssd1 vssd1 vccd1 vccd1 hold5931/A sky130_fd_sc_hd__buf_6
XTAP_6549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3642 _16660_/Q vssd1 vssd1 vccd1 vccd1 hold3642/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4387 _17122_/Q vssd1 vssd1 vccd1 vccd1 hold4387/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3653 _09865_/X vssd1 vssd1 vccd1 vccd1 _16445_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4398 _13888_/Y vssd1 vssd1 vccd1 vccd1 _17749_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3664 _16583_/Q vssd1 vssd1 vccd1 vccd1 hold3664/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3675 _10531_/X vssd1 vssd1 vccd1 vccd1 _16667_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2930 _17764_/Q vssd1 vssd1 vccd1 vccd1 hold2930/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2941 _14865_/X vssd1 vssd1 vccd1 vccd1 _18221_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3686 _16514_/Q vssd1 vssd1 vccd1 vccd1 hold3686/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2952 _17927_/Q vssd1 vssd1 vccd1 vccd1 hold2952/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3697 _13672_/X vssd1 vssd1 vccd1 vccd1 _17677_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2963 _14468_/X vssd1 vssd1 vccd1 vccd1 _18031_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2974 _14414_/X vssd1 vssd1 vccd1 vccd1 _18005_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2985 _17839_/Q vssd1 vssd1 vccd1 vccd1 hold2985/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2996 _14267_/X vssd1 vssd1 vccd1 vccd1 _17934_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10971_ _11067_/A _10971_/B vssd1 vssd1 vccd1 vccd1 _10971_/X sky130_fd_sc_hd__or2_1
XFILLER_0_97_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_458_wb_clk_i clkbuf_6_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17429_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12710_ hold3892/X _12709_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12711_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13690_ hold5412/X _13880_/B _13689_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13690_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12641_ hold3375/X _12640_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12642_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15360_ hold490/X _15448_/A2 _15446_/B1 hold531/X vssd1 vssd1 vccd1 vccd1 _15360_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_182_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12572_ hold3220/X _12571_/X _12971_/S vssd1 vssd1 vccd1 vccd1 _12572_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_182_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14311_ hold1851/X _14333_/A2 _14310_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _14311_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11523_ _12093_/A _11523_/B vssd1 vssd1 vccd1 vccd1 _11523_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15291_ _16293_/Q _15477_/A2 _15487_/B1 hold516/X _15290_/X vssd1 vssd1 vccd1 vccd1
+ _15292_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17030_ _17910_/CLK _17030_/D vssd1 vssd1 vccd1 vccd1 _17030_/Q sky130_fd_sc_hd__dfxtp_1
X_14242_ _15517_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14242_/X sky130_fd_sc_hd__or2_1
X_11454_ _11553_/A _11454_/B vssd1 vssd1 vccd1 vccd1 _11454_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10405_ hold3676/X _10619_/B _10404_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10405_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_1382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14173_ hold2505/X _14198_/B _14172_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _14173_/X
+ sky130_fd_sc_hd__o211a_1
X_11385_ _12174_/A _11385_/B vssd1 vssd1 vccd1 vccd1 _11385_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13124_ hold3479/X _13123_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13124_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_239_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10336_ hold3948/X _10649_/B _10335_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10336_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _17523_/Q _13056_/C _13055_/C _17522_/Q vssd1 vssd1 vccd1 vccd1 _13055_/X
+ sky130_fd_sc_hd__or4b_4
X_10267_ hold3326/X _10589_/B _10266_/X _14691_/C1 vssd1 vssd1 vccd1 vccd1 _10267_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17932_ _17968_/CLK _17932_/D vssd1 vssd1 vccd1 vccd1 _17932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12006_ _13716_/A _12006_/B vssd1 vssd1 vccd1 vccd1 _12006_/X sky130_fd_sc_hd__or2_1
XFILLER_0_206_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17863_ _17895_/CLK _17863_/D vssd1 vssd1 vccd1 vccd1 _17863_/Q sky130_fd_sc_hd__dfxtp_1
X_10198_ hold3884/X _10625_/B _10197_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _10198_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16814_ _18048_/CLK _16814_/D vssd1 vssd1 vccd1 vccd1 _16814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17794_ _17859_/CLK _17794_/D vssd1 vssd1 vccd1 vccd1 _17794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16745_ _18014_/CLK _16745_/D vssd1 vssd1 vccd1 vccd1 _16745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13957_ hold2627/X _13995_/A2 _13956_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _13957_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_199_wb_clk_i clkbuf_6_53_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18386_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_158_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12908_ hold3332/X _12907_/X _12923_/S vssd1 vssd1 vccd1 vccd1 _12908_/X sky130_fd_sc_hd__mux2_1
X_16676_ _18234_/CLK _16676_/D vssd1 vssd1 vccd1 vccd1 _16676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13888_ _13888_/A _13888_/B vssd1 vssd1 vccd1 vccd1 _13888_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_158_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_128_wb_clk_i clkbuf_6_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16090_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18415_ _18416_/CLK _18415_/D vssd1 vssd1 vccd1 vccd1 _18415_/Q sky130_fd_sc_hd__dfxtp_1
X_15627_ _17194_/CLK _15627_/D vssd1 vssd1 vccd1 vccd1 _15627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12839_ hold4052/X _12838_/X _12839_/S vssd1 vssd1 vccd1 vccd1 _12840_/B sky130_fd_sc_hd__mux2_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18346_ _18346_/CLK hold342/X vssd1 vssd1 vccd1 vccd1 _18346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15558_ hold1738/X _15560_/A2 _15557_/X _12849_/A vssd1 vssd1 vccd1 vccd1 _15558_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14509_ _14974_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14509_/X sky130_fd_sc_hd__or2_1
X_18277_ _18349_/CLK _18277_/D vssd1 vssd1 vccd1 vccd1 _18277_/Q sky130_fd_sc_hd__dfxtp_1
X_15489_ _15489_/A _15489_/B _15489_/C _15489_/D vssd1 vssd1 vccd1 vccd1 _15489_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08030_ hold2298/X _08029_/B _08029_/Y _08115_/A vssd1 vssd1 vccd1 vccd1 _08030_/X
+ sky130_fd_sc_hd__o211a_1
X_17228_ _17260_/CLK _17228_/D vssd1 vssd1 vccd1 vccd1 _17228_/Q sky130_fd_sc_hd__dfxtp_1
Xinput30 input30/A vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput41 input41/A vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput52 input52/A vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__buf_6
Xinput63 input63/A vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold803 hold803/A vssd1 vssd1 vccd1 vccd1 hold803/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold814 hold814/A vssd1 vssd1 vccd1 vccd1 hold814/X sky130_fd_sc_hd__dlygate4sd3_1
X_17159_ _17194_/CLK _17159_/D vssd1 vssd1 vccd1 vccd1 _17159_/Q sky130_fd_sc_hd__dfxtp_1
Xhold825 hold825/A vssd1 vssd1 vccd1 vccd1 hold825/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold836 hold836/A vssd1 vssd1 vccd1 vccd1 hold836/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold847 hold847/A vssd1 vssd1 vccd1 vccd1 hold847/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 hold858/A vssd1 vssd1 vccd1 vccd1 hold858/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 hold869/A vssd1 vssd1 vccd1 vccd1 hold869/X sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ _09981_/A _09981_/B vssd1 vssd1 vccd1 vccd1 _09981_/X sky130_fd_sc_hd__or2_1
XFILLER_0_229_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08932_ hold278/X hold649/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold650/A sky130_fd_sc_hd__mux2_1
XFILLER_0_149_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2204 _07891_/X vssd1 vssd1 vccd1 vccd1 _15589_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2215 _17885_/Q vssd1 vssd1 vccd1 vccd1 hold2215/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2226 hold2226/A vssd1 vssd1 vccd1 vccd1 input67/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2237 _14753_/X vssd1 vssd1 vccd1 vccd1 _18167_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1503 _18364_/Q vssd1 vssd1 vccd1 vccd1 hold1503/X sky130_fd_sc_hd__dlygate4sd3_1
X_08863_ _12426_/A hold557/X vssd1 vssd1 vccd1 vccd1 _16050_/D sky130_fd_sc_hd__and2_1
Xhold2248 _17893_/Q vssd1 vssd1 vccd1 vccd1 hold2248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2259 _18356_/Q vssd1 vssd1 vccd1 vccd1 hold2259/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1514 _08091_/X vssd1 vssd1 vccd1 vccd1 _15685_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1525 _17910_/Q vssd1 vssd1 vccd1 vccd1 hold1525/X sky130_fd_sc_hd__dlygate4sd3_1
X_07814_ _15539_/A _15103_/A _15535_/A _15099_/A vssd1 vssd1 vccd1 vccd1 _07817_/B
+ sky130_fd_sc_hd__or4_1
Xhold1536 _18059_/Q vssd1 vssd1 vccd1 vccd1 hold1536/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1547 _08024_/X vssd1 vssd1 vccd1 vccd1 _15653_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08794_ _15482_/A hold603/X vssd1 vssd1 vccd1 vccd1 _16017_/D sky130_fd_sc_hd__and2_1
Xhold1558 _17871_/Q vssd1 vssd1 vccd1 vccd1 hold1558/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1569 _08277_/X vssd1 vssd1 vccd1 vccd1 _15773_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09415_ _07804_/A _09456_/B _15284_/A _09414_/X vssd1 vssd1 vccd1 vccd1 _09415_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09346_ hold97/X hold220/A _09359_/C vssd1 vssd1 vccd1 vccd1 _09351_/B sky130_fd_sc_hd__or3_2
XFILLER_0_75_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09277_ _15553_/A hold2330/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09278_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08228_ _08504_/A _15128_/A vssd1 vssd1 vccd1 vccd1 _08228_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_50_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_1255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08159_ _08171_/A _08159_/B vssd1 vssd1 vccd1 vccd1 _15717_/D sky130_fd_sc_hd__and2_1
XFILLER_0_222_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11170_ _12301_/A _11170_/B vssd1 vssd1 vccd1 vccd1 _16880_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_28_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4140 hold5928/X vssd1 vssd1 vccd1 vccd1 hold5929/A sky130_fd_sc_hd__buf_4
XFILLER_0_30_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10121_ hold2282/X _16531_/Q _10601_/C vssd1 vssd1 vccd1 vccd1 _10122_/B sky130_fd_sc_hd__mux2_1
Xhold4151 _17495_/Q vssd1 vssd1 vccd1 vccd1 hold4151/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4162 _11419_/X vssd1 vssd1 vccd1 vccd1 _16963_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4173 _17000_/Q vssd1 vssd1 vccd1 vccd1 hold4173/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4184 _15490_/X vssd1 vssd1 vccd1 vccd1 _15491_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4195 hold5936/X vssd1 vssd1 vccd1 vccd1 hold5937/A sky130_fd_sc_hd__buf_6
Xhold3450 _16731_/Q vssd1 vssd1 vccd1 vccd1 hold3450/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3461 hold3810/X vssd1 vssd1 vccd1 vccd1 _10601_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10052_ _16508_/Q _10052_/B _10538_/S vssd1 vssd1 vccd1 vccd1 _10052_/X sky130_fd_sc_hd__and3_1
XTAP_6379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3472 _12310_/Y vssd1 vssd1 vccd1 vccd1 _17260_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3483 _16722_/Q vssd1 vssd1 vccd1 vccd1 hold3483/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3494 _13869_/Y vssd1 vssd1 vccd1 vccd1 _13870_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2760 _15622_/Q vssd1 vssd1 vccd1 vccd1 hold2760/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14860_ _15145_/A _14892_/B vssd1 vssd1 vccd1 vccd1 _14860_/X sky130_fd_sc_hd__or2_1
XTAP_5678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2771 _17845_/Q vssd1 vssd1 vccd1 vccd1 hold2771/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2782 _14524_/X vssd1 vssd1 vccd1 vccd1 _18058_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2793 _07919_/X vssd1 vssd1 vccd1 vccd1 _15603_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ _17724_/Q _13811_/B _13811_/C vssd1 vssd1 vccd1 vccd1 _13811_/X sky130_fd_sc_hd__and3_1
XFILLER_0_203_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14791_ hold1998/X _14826_/B _14790_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14791_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_292_wb_clk_i clkbuf_6_39_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18065_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_225_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16530_ _18228_/CLK _16530_/D vssd1 vssd1 vccd1 vccd1 _16530_/Q sky130_fd_sc_hd__dfxtp_1
X_13742_ hold2942/X _17701_/Q _13871_/C vssd1 vssd1 vccd1 vccd1 _13743_/B sky130_fd_sc_hd__mux2_1
X_10954_ hold3771/X _11144_/B _10953_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _10954_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_221_wb_clk_i clkbuf_6_61_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18223_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16461_ _18374_/CLK _16461_/D vssd1 vssd1 vccd1 vccd1 _16461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13673_ hold2848/X hold4003/X _13766_/S vssd1 vssd1 vccd1 vccd1 _13674_/B sky130_fd_sc_hd__mux2_1
X_10885_ hold5060/X _11165_/B _10884_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _10885_/X
+ sky130_fd_sc_hd__o211a_1
X_18200_ _18200_/CLK _18200_/D vssd1 vssd1 vccd1 vccd1 _18200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15412_ _15489_/A _15412_/B _15412_/C _15412_/D vssd1 vssd1 vccd1 vccd1 _15412_/X
+ sky130_fd_sc_hd__or4_1
XPHY_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12624_ _12864_/A _12624_/B vssd1 vssd1 vccd1 vccd1 _17384_/D sky130_fd_sc_hd__and2_1
XPHY_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16392_ _18373_/CLK _16392_/D vssd1 vssd1 vccd1 vccd1 _16392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18131_ _18197_/CLK _18131_/D vssd1 vssd1 vccd1 vccd1 _18131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15343_ _15481_/A1 _15335_/X _15342_/X _15481_/B1 hold5929/A vssd1 vssd1 vccd1 vccd1
+ _15343_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12555_ _12948_/A _12555_/B vssd1 vssd1 vccd1 vccd1 _17361_/D sky130_fd_sc_hd__and2_1
XFILLER_0_93_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18062_ _18347_/CLK _18062_/D vssd1 vssd1 vccd1 vccd1 _18062_/Q sky130_fd_sc_hd__dfxtp_1
X_11506_ hold5404/X _12335_/B _11505_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _11506_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15274_ _15274_/A _15274_/B vssd1 vssd1 vccd1 vccd1 _18403_/D sky130_fd_sc_hd__and2_1
XFILLER_0_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12486_ _17336_/Q _12506_/B vssd1 vssd1 vccd1 vccd1 _12486_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17013_ _17861_/CLK _17013_/D vssd1 vssd1 vccd1 vccd1 _17013_/Q sky130_fd_sc_hd__dfxtp_1
X_14225_ hold2125/X _14216_/Y _14224_/X _14354_/A vssd1 vssd1 vccd1 vccd1 _14225_/X
+ sky130_fd_sc_hd__o211a_1
X_11437_ hold5368/X _11726_/B _11436_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _11437_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14156_ hold820/X _14160_/B vssd1 vssd1 vccd1 vccd1 _14156_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11368_ hold5140/X _11753_/B _11367_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _11368_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_237_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13107_ _13106_/X _16906_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13107_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10319_ hold2815/X _16597_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10320_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14087_ hold2218/X _14094_/B _14086_/X _12588_/A vssd1 vssd1 vccd1 vccd1 _14087_/X
+ sky130_fd_sc_hd__o211a_1
X_11299_ hold5138/X _12323_/B _11298_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _11299_/X
+ sky130_fd_sc_hd__o211a_1
X_13038_ _13048_/A _13034_/X _17523_/Q vssd1 vssd1 vccd1 vccd1 _13039_/B sky130_fd_sc_hd__a21o_1
X_17915_ _17976_/CLK _17915_/D vssd1 vssd1 vccd1 vccd1 _17915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17846_ _17846_/CLK _17846_/D vssd1 vssd1 vccd1 vccd1 _17846_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_309_wb_clk_i clkbuf_6_45_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18059_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14989_ hold2548/X _15004_/B _14988_/X _15048_/A vssd1 vssd1 vccd1 vccd1 _14989_/X
+ sky130_fd_sc_hd__o211a_1
X_17777_ _17843_/CLK _17777_/D vssd1 vssd1 vccd1 vccd1 _17777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16728_ _18057_/CLK _16728_/D vssd1 vssd1 vccd1 vccd1 _16728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_232_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16659_ _18217_/CLK _16659_/D vssd1 vssd1 vccd1 vccd1 _16659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09200_ _15529_/A _09206_/B vssd1 vssd1 vccd1 vccd1 _09200_/X sky130_fd_sc_hd__or2_1
XFILLER_0_53_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09131_ hold2924/X _09177_/A2 _09130_/X _12855_/A vssd1 vssd1 vccd1 vccd1 _09131_/X
+ sky130_fd_sc_hd__o211a_1
X_18329_ _18361_/CLK _18329_/D vssd1 vssd1 vccd1 vccd1 _18329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_10_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_10_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_09062_ hold278/X hold387/X _09062_/S vssd1 vssd1 vccd1 vccd1 hold388/A sky130_fd_sc_hd__mux2_1
XFILLER_0_127_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_96_wb_clk_i clkbuf_6_22_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18406_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_142_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08013_ hold951/X _08045_/B vssd1 vssd1 vccd1 vccd1 _08013_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold600 hold600/A vssd1 vssd1 vccd1 vccd1 hold600/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 hold611/A vssd1 vssd1 vccd1 vccd1 hold611/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_wb_clk_i clkbuf_6_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17360_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold622 hold622/A vssd1 vssd1 vccd1 vccd1 hold622/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 hold633/A vssd1 vssd1 vccd1 vccd1 hold633/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold644 hold644/A vssd1 vssd1 vccd1 vccd1 hold644/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold655 hold655/A vssd1 vssd1 vccd1 vccd1 hold655/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold666 hold666/A vssd1 vssd1 vccd1 vccd1 hold666/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 hold677/A vssd1 vssd1 vccd1 vccd1 input34/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 hold688/A vssd1 vssd1 vccd1 vccd1 hold688/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 hold699/A vssd1 vssd1 vccd1 vccd1 hold699/X sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ hold3944/X _10598_/B _09963_/X _15218_/C1 vssd1 vssd1 vccd1 vccd1 _09964_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2001 _15550_/X vssd1 vssd1 vccd1 vccd1 _18453_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2012 _08316_/X vssd1 vssd1 vccd1 vccd1 _15791_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08915_ _12426_/A hold430/X vssd1 vssd1 vccd1 vccd1 _16075_/D sky130_fd_sc_hd__and2_1
XFILLER_0_110_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2023 _17805_/Q vssd1 vssd1 vccd1 vccd1 hold2023/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2034 _14737_/X vssd1 vssd1 vccd1 vccd1 _18159_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09895_ hold3658/X _10004_/B _09894_/X _15042_/A vssd1 vssd1 vccd1 vccd1 _09895_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2045 _16316_/Q vssd1 vssd1 vccd1 vccd1 _09472_/C sky130_fd_sc_hd__clkbuf_2
Xhold1300 _14961_/X vssd1 vssd1 vccd1 vccd1 _18267_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1311 _18205_/Q vssd1 vssd1 vccd1 vccd1 hold1311/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2056 _17879_/Q vssd1 vssd1 vccd1 vccd1 hold2056/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1322 _14179_/X vssd1 vssd1 vccd1 vccd1 _17892_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08846_ hold373/X hold633/X _08866_/S vssd1 vssd1 vccd1 vccd1 _08847_/B sky130_fd_sc_hd__mux2_1
Xhold2067 _14452_/X vssd1 vssd1 vccd1 vccd1 _18023_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1333 _08328_/X vssd1 vssd1 vccd1 vccd1 _15797_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2078 _08051_/X vssd1 vssd1 vccd1 vccd1 _15665_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2089 _14265_/X vssd1 vssd1 vccd1 vccd1 _17933_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1344 _15634_/Q vssd1 vssd1 vccd1 vccd1 hold1344/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1355 _07989_/X vssd1 vssd1 vccd1 vccd1 _15637_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1366 input59/X vssd1 vssd1 vccd1 vccd1 hold910/A sky130_fd_sc_hd__buf_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1377 _08516_/X vssd1 vssd1 vccd1 vccd1 _15885_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08777_ hold92/X hold611/X _08793_/S vssd1 vssd1 vccd1 vccd1 hold612/A sky130_fd_sc_hd__mux2_1
XFILLER_0_169_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1388 _18321_/Q vssd1 vssd1 vccd1 vccd1 hold1388/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1399 _18305_/Q vssd1 vssd1 vccd1 vccd1 hold1399/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10670_ hold2514/X hold4469/X _11726_/C vssd1 vssd1 vccd1 vccd1 _10671_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_193_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09329_ hold992/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09329_/X sky130_fd_sc_hd__or2_1
XFILLER_0_192_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12340_ _13873_/A _12340_/B vssd1 vssd1 vccd1 vccd1 _12340_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_211_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12271_ hold4005/X _12365_/B _12270_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _12271_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14010_ _14457_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14010_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11222_ _16898_/Q _11222_/B _11789_/C vssd1 vssd1 vccd1 vccd1 _11222_/X sky130_fd_sc_hd__and3_1
XTAP_6110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11153_ _16875_/Q _11153_/B _11153_/C vssd1 vssd1 vccd1 vccd1 _11153_/X sky130_fd_sc_hd__and3_1
XFILLER_0_101_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10104_ _10530_/A _10104_/B vssd1 vssd1 vccd1 vccd1 _10104_/X sky130_fd_sc_hd__or2_1
XTAP_6154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15961_ _17321_/CLK _15961_/D vssd1 vssd1 vccd1 vccd1 hold851/A sky130_fd_sc_hd__dfxtp_1
X_11084_ hold1295/X hold4925/X _11204_/C vssd1 vssd1 vccd1 vccd1 _11085_/B sky130_fd_sc_hd__mux2_1
XTAP_6165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3280 _16635_/Q vssd1 vssd1 vccd1 vccd1 hold3280/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10035_ _13206_/A _09957_/A _10034_/X vssd1 vssd1 vccd1 vccd1 _10035_/Y sky130_fd_sc_hd__a21oi_1
X_14912_ hold406/X _15182_/B vssd1 vssd1 vccd1 vccd1 _14912_/Y sky130_fd_sc_hd__nor2_2
X_17700_ _17732_/CLK _17700_/D vssd1 vssd1 vccd1 vccd1 _17700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3291 _12596_/X vssd1 vssd1 vccd1 vccd1 _12597_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15892_ _16139_/CLK _15892_/D vssd1 vssd1 vccd1 vccd1 hold735/A sky130_fd_sc_hd__dfxtp_1
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2590 _08275_/X vssd1 vssd1 vccd1 vccd1 _15772_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_402_wb_clk_i clkbuf_6_37_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18050_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ hold330/X _14843_/B vssd1 vssd1 vccd1 vccd1 _14892_/B sky130_fd_sc_hd__or2_4
X_17631_ _17729_/CLK _17631_/D vssd1 vssd1 vccd1 vccd1 _17631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17562_ _17624_/CLK _17562_/D vssd1 vssd1 vccd1 vccd1 _17562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14774_ _14952_/A _14774_/B vssd1 vssd1 vccd1 vccd1 _14774_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_230_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11986_ hold4046/X _13886_/B _11985_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _11986_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16513_ _18298_/CLK _16513_/D vssd1 vssd1 vccd1 vccd1 _16513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13725_ _13734_/A _13725_/B vssd1 vssd1 vccd1 vccd1 _13725_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17493_ _17493_/CLK _17493_/D vssd1 vssd1 vccd1 vccd1 _17493_/Q sky130_fd_sc_hd__dfxtp_1
X_10937_ hold2805/X hold3824/X _11219_/C vssd1 vssd1 vccd1 vccd1 _10938_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16444_ _18357_/CLK _16444_/D vssd1 vssd1 vccd1 vccd1 _16444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13656_ _13752_/A _13656_/B vssd1 vssd1 vccd1 vccd1 _13656_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10868_ hold2015/X hold3324/X _11153_/C vssd1 vssd1 vccd1 vccd1 _10869_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12607_ hold1309/X _17380_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12607_/X sky130_fd_sc_hd__mux2_1
X_16375_ _18352_/CLK _16375_/D vssd1 vssd1 vccd1 vccd1 _16375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13587_ _13758_/A _13587_/B vssd1 vssd1 vccd1 vccd1 _13587_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ hold2850/X hold5181/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10800_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18114_ _18129_/CLK _18114_/D vssd1 vssd1 vccd1 vccd1 _18114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15326_ _17336_/Q _15486_/B1 _15485_/B1 hold100/X vssd1 vssd1 vccd1 vccd1 _15326_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12538_ hold1242/X hold4517/X _12925_/S vssd1 vssd1 vccd1 vccd1 _12538_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18045_ _18045_/CLK hold879/X vssd1 vssd1 vccd1 vccd1 hold878/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15257_ hold303/X _09357_/A _15484_/B1 hold460/X _15256_/X vssd1 vssd1 vccd1 vccd1
+ _15262_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_125_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12469_ hold163/X _12445_/A _12445_/B _12468_/X _12438_/A vssd1 vssd1 vccd1 vccd1
+ hold3/A sky130_fd_sc_hd__o311a_1
XFILLER_0_111_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4909 _16758_/Q vssd1 vssd1 vccd1 vccd1 hold4909/X sky130_fd_sc_hd__dlygate4sd3_1
X_14208_ _14726_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14208_/X sky130_fd_sc_hd__or2_1
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15188_ hold1847/X _15219_/B _15187_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _15188_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14139_ hold1570/X _14142_/B _14138_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _14139_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout409 _14282_/B vssd1 vssd1 vccd1 vccd1 _14284_/B sky130_fd_sc_hd__buf_6
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08700_ _15324_/A _08700_/B vssd1 vssd1 vccd1 vccd1 _15971_/D sky130_fd_sc_hd__and2_1
X_09680_ hold1527/X _16384_/Q _10067_/C vssd1 vssd1 vccd1 vccd1 _09681_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_143_wb_clk_i clkbuf_6_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18372_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08631_ hold185/X _15938_/Q _08657_/S vssd1 vssd1 vccd1 vccd1 hold186/A sky130_fd_sc_hd__mux2_1
X_17829_ _17840_/CLK _17829_/D vssd1 vssd1 vccd1 vccd1 _17829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08562_ hold180/X hold542/X _08592_/S vssd1 vssd1 vccd1 vccd1 hold543/A sky130_fd_sc_hd__mux2_1
XFILLER_0_194_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08493_ hold1442/X _08486_/B _08492_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _08493_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09114_ _15555_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09114_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09045_ _15314_/A _09045_/B vssd1 vssd1 vccd1 vccd1 _16139_/D sky130_fd_sc_hd__and2_1
XFILLER_0_27_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold430 hold430/A vssd1 vssd1 vccd1 vccd1 hold430/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 la_data_in[26] vssd1 vssd1 vccd1 vccd1 hold441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 hold452/A vssd1 vssd1 vccd1 vccd1 hold452/X sky130_fd_sc_hd__buf_4
Xhold463 hold463/A vssd1 vssd1 vccd1 vccd1 hold463/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold474 hold474/A vssd1 vssd1 vccd1 vccd1 hold474/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 hold485/A vssd1 vssd1 vccd1 vccd1 hold485/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 hold496/A vssd1 vssd1 vccd1 vccd1 hold496/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout910 hold820/X vssd1 vssd1 vccd1 vccd1 _15555_/A sky130_fd_sc_hd__buf_12
Xfanout921 hold484/X vssd1 vssd1 vccd1 vccd1 _14543_/A sky130_fd_sc_hd__clkbuf_8
X_09947_ hold1434/X hold4638/X _10031_/C vssd1 vssd1 vccd1 vccd1 _09948_/B sky130_fd_sc_hd__mux2_1
Xfanout932 hold630/X vssd1 vssd1 vccd1 vccd1 _15103_/A sky130_fd_sc_hd__clkbuf_16
Xfanout943 _15203_/A vssd1 vssd1 vccd1 vccd1 _14988_/A sky130_fd_sc_hd__buf_12
XFILLER_0_217_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ hold2211/X _16450_/Q _11204_/C vssd1 vssd1 vccd1 vccd1 _09879_/B sky130_fd_sc_hd__mux2_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 _16181_/Q vssd1 vssd1 vccd1 vccd1 hold1130/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 _15755_/Q vssd1 vssd1 vccd1 vccd1 hold1141/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08829_ _15374_/A _08829_/B vssd1 vssd1 vccd1 vccd1 _16033_/D sky130_fd_sc_hd__and2_1
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1152 hold1152/A vssd1 vssd1 vccd1 vccd1 input38/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1163 _16154_/Q vssd1 vssd1 vccd1 vccd1 hold1163/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1174 _08038_/X vssd1 vssd1 vccd1 vccd1 _15660_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1185 _09259_/X vssd1 vssd1 vccd1 vccd1 _09260_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1196 _17766_/Q vssd1 vssd1 vccd1 vccd1 hold1196/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11840_ hold1015/X _17104_/Q _12227_/S vssd1 vssd1 vccd1 vccd1 _11841_/B sky130_fd_sc_hd__mux2_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11771_ _17081_/Q _11771_/B _12242_/S vssd1 vssd1 vccd1 vccd1 _11771_/X sky130_fd_sc_hd__and3_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ hold5084/X _13814_/B _13509_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _13510_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10722_ _11106_/A _10722_/B vssd1 vssd1 vccd1 vccd1 _10722_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ hold1867/X _14487_/B _14489_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _14490_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13441_ hold4703/X _13795_/A2 _13440_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _13441_/X
+ sky130_fd_sc_hd__o211a_1
X_10653_ _11637_/A _10653_/B vssd1 vssd1 vccd1 vccd1 _10653_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16160_ _17500_/CLK _16160_/D vssd1 vssd1 vccd1 vccd1 _16160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13372_ hold5472/X _13880_/B _13371_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13372_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10584_ hold3501/X _10524_/A _10583_/X vssd1 vssd1 vccd1 vccd1 _10584_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15111_ _15165_/A hold341/X vssd1 vssd1 vccd1 vccd1 _15111_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_140_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12323_ _12323_/A _12323_/B _12323_/C vssd1 vssd1 vccd1 vccd1 _12323_/X sky130_fd_sc_hd__and3_1
X_16091_ _17300_/CLK _16091_/D vssd1 vssd1 vccd1 vccd1 hold667/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_1347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15042_ _15042_/A _15042_/B vssd1 vssd1 vccd1 vccd1 _18306_/D sky130_fd_sc_hd__and2_1
X_12254_ hold1762/X hold4739/X _13463_/S vssd1 vssd1 vccd1 vccd1 _12255_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11205_ hold4326/X _11109_/A _11204_/X vssd1 vssd1 vccd1 vccd1 _11205_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12185_ hold2792/X hold5156/X _13886_/C vssd1 vssd1 vccd1 vccd1 _12186_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_236_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_222_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11136_ _11136_/A _11136_/B vssd1 vssd1 vccd1 vccd1 _11136_/X sky130_fd_sc_hd__or2_1
X_16993_ _17873_/CLK _16993_/D vssd1 vssd1 vccd1 vccd1 _16993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15944_ _17314_/CLK _15944_/D vssd1 vssd1 vccd1 vccd1 hold793/A sky130_fd_sc_hd__dfxtp_1
X_11067_ _11067_/A _11067_/B vssd1 vssd1 vccd1 vccd1 _11067_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10018_ _11158_/A _10018_/B vssd1 vssd1 vccd1 vccd1 _16496_/D sky130_fd_sc_hd__nor2_1
XTAP_5294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15875_ _17653_/CLK _15875_/D vssd1 vssd1 vccd1 vccd1 _15875_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14826_ _15165_/A _14826_/B vssd1 vssd1 vccd1 vccd1 _14826_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_204_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17614_ _17614_/CLK _17614_/D vssd1 vssd1 vccd1 vccd1 _17614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17545_ _18392_/CLK _17545_/D vssd1 vssd1 vccd1 vccd1 _17545_/Q sky130_fd_sc_hd__dfxtp_1
X_14757_ hold2743/X _14772_/B _14756_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14757_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11969_ hold2503/X _17147_/Q _13409_/S vssd1 vssd1 vccd1 vccd1 _11970_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13708_ hold4737/X _13814_/B _13707_/X _08361_/A vssd1 vssd1 vccd1 vccd1 _13708_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17476_ _17476_/CLK _17476_/D vssd1 vssd1 vccd1 vccd1 _17476_/Q sky130_fd_sc_hd__dfxtp_1
X_14688_ _15189_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14688_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16427_ _18374_/CLK _16427_/D vssd1 vssd1 vccd1 vccd1 _16427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13639_ hold4569/X _13829_/B _13638_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13639_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16358_ _18411_/CLK _16358_/D vssd1 vssd1 vccd1 vccd1 _16358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6108 _09443_/Y vssd1 vssd1 vccd1 vccd1 _16307_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6119 la_data_in[2] vssd1 vssd1 vccd1 vccd1 hold6119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15309_ hold846/X _09365_/B _09392_/C hold890/X _15308_/X vssd1 vssd1 vccd1 vccd1
+ _15312_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16289_ _18404_/CLK _16289_/D vssd1 vssd1 vccd1 vccd1 _16289_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5407 _11629_/X vssd1 vssd1 vccd1 vccd1 _17033_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_129_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5418 _17619_/Q vssd1 vssd1 vccd1 vccd1 hold5418/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5429 _11572_/X vssd1 vssd1 vccd1 vccd1 _17014_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4706 _10933_/X vssd1 vssd1 vccd1 vccd1 _16801_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18028_ _18028_/CLK _18028_/D vssd1 vssd1 vccd1 vccd1 _18028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4717 _16921_/Q vssd1 vssd1 vccd1 vccd1 hold4717/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4728 _10972_/X vssd1 vssd1 vccd1 vccd1 _16814_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4739 _17242_/Q vssd1 vssd1 vccd1 vccd1 hold4739/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_395_wb_clk_i clkbuf_6_36_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17868_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_227_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout206 _11222_/B vssd1 vssd1 vccd1 vccd1 _11789_/B sky130_fd_sc_hd__buf_4
XFILLER_0_240_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout217 _10013_/B vssd1 vssd1 vccd1 vccd1 _11201_/B sky130_fd_sc_hd__buf_4
X_09801_ _09987_/A _09801_/B vssd1 vssd1 vccd1 vccd1 _09801_/X sky130_fd_sc_hd__or2_1
XFILLER_0_61_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_324_wb_clk_i clkbuf_6_46_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17269_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout228 _10616_/B vssd1 vssd1 vccd1 vccd1 _11213_/B sky130_fd_sc_hd__buf_4
Xfanout239 _10067_/B vssd1 vssd1 vccd1 vccd1 _10577_/B sky130_fd_sc_hd__buf_4
X_07993_ _08504_/A _09498_/A vssd1 vssd1 vccd1 vccd1 _07993_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_66_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09732_ _09978_/A _09732_/B vssd1 vssd1 vccd1 vccd1 _09732_/X sky130_fd_sc_hd__or2_1
XFILLER_0_198_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09663_ _09978_/A _09663_/B vssd1 vssd1 vccd1 vccd1 _09663_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08614_ _09061_/A hold778/X vssd1 vssd1 vccd1 vccd1 _15929_/D sky130_fd_sc_hd__and2_1
X_09594_ _10482_/A _09594_/B vssd1 vssd1 vccd1 vccd1 _09594_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08545_ _09061_/A hold197/X vssd1 vssd1 vccd1 vccd1 _15896_/D sky130_fd_sc_hd__and2_1
XFILLER_0_77_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08476_ _14529_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08476_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_40_wb_clk_i clkbuf_6_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17846_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_18_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09028_ hold172/X hold644/X _09060_/S vssd1 vssd1 vccd1 vccd1 _09029_/B sky130_fd_sc_hd__mux2_1
Xhold5930 _16280_/Q vssd1 vssd1 vccd1 vccd1 hold5930/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5941 hold5941/A vssd1 vssd1 vccd1 vccd1 hold5941/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5952 hold5952/A vssd1 vssd1 vccd1 vccd1 hold5952/X sky130_fd_sc_hd__clkbuf_4
Xhold5963 hold5963/A vssd1 vssd1 vccd1 vccd1 hold5963/X sky130_fd_sc_hd__clkbuf_4
Xhold5974 hold5974/A vssd1 vssd1 vccd1 vccd1 hold5974/X sky130_fd_sc_hd__buf_4
Xhold260 hold260/A vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5985 _09467_/Y vssd1 vssd1 vccd1 vccd1 _16316_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5996 _16527_/Q vssd1 vssd1 vccd1 vccd1 hold5996/X sky130_fd_sc_hd__buf_1
Xhold271 hold271/A vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__clkbuf_8
Xhold282 hold282/A vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 hold358/X vssd1 vssd1 vccd1 vccd1 hold359/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout740 _13675_/C1 vssd1 vssd1 vccd1 vccd1 _08377_/A sky130_fd_sc_hd__buf_4
XFILLER_0_102_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout751 _08119_/A vssd1 vssd1 vccd1 vccd1 _08133_/A sky130_fd_sc_hd__buf_4
Xfanout762 _14528_/C1 vssd1 vssd1 vccd1 vccd1 _14462_/C1 sky130_fd_sc_hd__buf_4
Xfanout773 _08385_/A vssd1 vssd1 vccd1 vccd1 _13792_/C1 sky130_fd_sc_hd__buf_4
X_13990_ _14330_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13990_/X sky130_fd_sc_hd__or2_1
XFILLER_0_219_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_233_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout784 _14143_/C1 vssd1 vssd1 vccd1 vccd1 _13943_/A sky130_fd_sc_hd__buf_4
Xfanout795 _15054_/A vssd1 vssd1 vccd1 vccd1 _15202_/C1 sky130_fd_sc_hd__buf_4
X_12941_ hold4467/X _12940_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12941_/X sky130_fd_sc_hd__mux2_1
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15660_ _17270_/CLK _15660_/D vssd1 vssd1 vccd1 vccd1 _15660_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ hold3120/X _12871_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12872_/X sky130_fd_sc_hd__mux2_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 _14479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_111 _14988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ hold2594/X _14610_/B _14610_/Y _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14611_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_122 _15173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11823_ _13716_/A _11823_/B vssd1 vssd1 vccd1 vccd1 _11823_/X sky130_fd_sc_hd__or2_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _17271_/CLK _15591_/D vssd1 vssd1 vccd1 vccd1 _15591_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17330_ _18410_/CLK hold173/X vssd1 vssd1 vccd1 vccd1 _17330_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14542_ hold2353/X _14541_/B _14541_/Y _14542_/C1 vssd1 vssd1 vccd1 vccd1 _14542_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11754_ hold4751/X _11658_/A _11753_/X vssd1 vssd1 vccd1 vccd1 _11754_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_166_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ hold5181/X _11225_/B _10704_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _10705_/X
+ sky130_fd_sc_hd__o211a_1
X_17261_ _17261_/CLK _17261_/D vssd1 vssd1 vccd1 vccd1 _17261_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14473_ _15099_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14473_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11685_ _12219_/A _11685_/B vssd1 vssd1 vccd1 vccd1 _11685_/X sky130_fd_sc_hd__or2_1
XFILLER_0_187_1250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16212_ _17725_/CLK _16212_/D vssd1 vssd1 vccd1 vccd1 _16212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13424_ hold2388/X _17595_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13425_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_180_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10636_ _11206_/A _10636_/B vssd1 vssd1 vccd1 vccd1 _16702_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17192_ _17724_/CLK _17192_/D vssd1 vssd1 vccd1 vccd1 _17192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16143_ _17299_/CLK _16143_/D vssd1 vssd1 vccd1 vccd1 hold864/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13355_ hold1043/X hold4378/X _13871_/C vssd1 vssd1 vccd1 vccd1 _13356_/B sky130_fd_sc_hd__mux2_1
X_10567_ _10603_/A _10567_/B vssd1 vssd1 vccd1 vccd1 _16679_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_183_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12306_ hold4471/X _12093_/A _12305_/X vssd1 vssd1 vccd1 vccd1 _12306_/Y sky130_fd_sc_hd__a21oi_1
X_16074_ _18405_/CLK _16074_/D vssd1 vssd1 vccd1 vccd1 hold399/A sky130_fd_sc_hd__dfxtp_1
X_13286_ _13286_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13286_/X sky130_fd_sc_hd__or2_1
X_10498_ hold3730/X _10598_/B _10497_/X _15019_/C1 vssd1 vssd1 vccd1 vccd1 _10498_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_220_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15025_ _15187_/A hold1917/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15025_/X sky130_fd_sc_hd__mux2_1
X_12237_ _12255_/A _12237_/B vssd1 vssd1 vccd1 vccd1 _12237_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12168_ _12267_/A _12168_/B vssd1 vssd1 vccd1 vccd1 _12168_/X sky130_fd_sc_hd__or2_1
XFILLER_0_194_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11119_ hold4881/X _11225_/B _11118_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _11119_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12099_ _13797_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12099_/X sky130_fd_sc_hd__or2_1
X_16976_ _17888_/CLK _16976_/D vssd1 vssd1 vccd1 vccd1 _16976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput6 input6/A vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
X_15927_ _17345_/CLK _15927_/D vssd1 vssd1 vccd1 vccd1 hold560/A sky130_fd_sc_hd__dfxtp_1
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ _17599_/CLK _15858_/D vssd1 vssd1 vccd1 vccd1 _15858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14809_ hold2928/X _14828_/B _14808_/X _14342_/A vssd1 vssd1 vccd1 vccd1 _14809_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15789_ _17426_/CLK _15789_/D vssd1 vssd1 vccd1 vccd1 _15789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08330_ hold2499/X _08336_/A2 _08329_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08330_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17528_ _17533_/CLK _17528_/D vssd1 vssd1 vccd1 vccd1 _17528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08261_ hold1793/X _08262_/B _08260_/X _08347_/A vssd1 vssd1 vccd1 vccd1 _08261_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17459_ _18455_/CLK _17459_/D vssd1 vssd1 vccd1 vccd1 _17459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08192_ hold2234/X _08213_/B _08191_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _08192_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5204 _13744_/X vssd1 vssd1 vccd1 vccd1 _17701_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5215 _16782_/Q vssd1 vssd1 vccd1 vccd1 hold5215/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5226 _11710_/X vssd1 vssd1 vccd1 vccd1 _17060_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5237 _17218_/Q vssd1 vssd1 vccd1 vccd1 hold5237/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4503 _17487_/Q vssd1 vssd1 vccd1 vccd1 hold4503/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5248 _11116_/X vssd1 vssd1 vccd1 vccd1 _16862_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4514 _17587_/Q vssd1 vssd1 vccd1 vccd1 hold4514/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5259 _17077_/Q vssd1 vssd1 vccd1 vccd1 hold5259/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4525 _16638_/Q vssd1 vssd1 vccd1 vccd1 hold4525/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4536 _17356_/Q vssd1 vssd1 vccd1 vccd1 hold4536/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4547 _16468_/Q vssd1 vssd1 vccd1 vccd1 hold4547/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3802 _13768_/X vssd1 vssd1 vccd1 vccd1 _17709_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4558 _09727_/X vssd1 vssd1 vccd1 vccd1 _16399_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3813 _17432_/Q vssd1 vssd1 vccd1 vccd1 hold3813/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3824 _16803_/Q vssd1 vssd1 vccd1 vccd1 hold3824/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4569 _17698_/Q vssd1 vssd1 vccd1 vccd1 hold4569/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3835 _10111_/X vssd1 vssd1 vccd1 vccd1 _16527_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3846 _16614_/Q vssd1 vssd1 vccd1 vccd1 hold3846/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3857 _12217_/X vssd1 vssd1 vccd1 vccd1 _17229_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3868 _16871_/Q vssd1 vssd1 vccd1 vccd1 hold3868/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3879 _10444_/X vssd1 vssd1 vccd1 vccd1 _16638_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07976_ _15545_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _07976_/Y sky130_fd_sc_hd__nand2_1
X_09715_ hold3640/X _10025_/B _09714_/X _15473_/A vssd1 vssd1 vccd1 vccd1 _09715_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09646_ hold4545/X _10028_/B _09645_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09646_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ hold3545/X _10601_/B _09576_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09577_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08528_ hold131/X hold475/X _08528_/S vssd1 vssd1 vccd1 vccd1 hold476/A sky130_fd_sc_hd__mux2_1
XFILLER_0_38_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08459_ hold2367/X _08488_/B _08458_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08459_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11470_ hold5362/X _11195_/B _11469_/X _14462_/C1 vssd1 vssd1 vccd1 vccd1 _11470_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10421_ hold2522/X _16631_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10422_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_246_wb_clk_i clkbuf_6_59_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18168_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13140_ hold4284/X _13139_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13140_/X sky130_fd_sc_hd__mux2_1
X_10352_ hold1113/X _16608_/Q _10646_/C vssd1 vssd1 vccd1 vccd1 _10353_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5760 _12253_/X vssd1 vssd1 vccd1 vccd1 _17241_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13071_ _13199_/A1 _13069_/X _13070_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13071_/X
+ sky130_fd_sc_hd__o211a_1
X_10283_ hold2659/X hold3292/X _10571_/C vssd1 vssd1 vccd1 vccd1 _10284_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5771 _17246_/Q vssd1 vssd1 vccd1 vccd1 hold5771/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5782 _13615_/X vssd1 vssd1 vccd1 vccd1 _17658_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5793 _17274_/Q vssd1 vssd1 vccd1 vccd1 hold5793/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12022_ hold4587/X _12308_/B _12021_/X _08167_/A vssd1 vssd1 vccd1 vccd1 _12022_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_1302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16830_ _18065_/CLK _16830_/D vssd1 vssd1 vccd1 vccd1 _16830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout570 _07916_/B vssd1 vssd1 vccd1 vccd1 _07936_/B sky130_fd_sc_hd__buf_8
Xfanout581 _13057_/X vssd1 vssd1 vccd1 vccd1 _13250_/S sky130_fd_sc_hd__buf_8
Xfanout592 _12811_/S vssd1 vssd1 vccd1 vccd1 _12838_/S sky130_fd_sc_hd__buf_6
X_13973_ hold1289/X _13995_/A2 _13972_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _13973_/X
+ sky130_fd_sc_hd__o211a_1
X_16761_ _17964_/CLK _16761_/D vssd1 vssd1 vccd1 vccd1 _16761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15712_ _17271_/CLK _15712_/D vssd1 vssd1 vccd1 vccd1 _15712_/Q sky130_fd_sc_hd__dfxtp_1
X_12924_ _12924_/A _12924_/B vssd1 vssd1 vccd1 vccd1 _17484_/D sky130_fd_sc_hd__and2_1
X_16692_ _18220_/CLK _16692_/D vssd1 vssd1 vccd1 vccd1 _16692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18431_ _18432_/CLK hold425/X vssd1 vssd1 vccd1 vccd1 _18431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15643_ _17153_/CLK _15643_/D vssd1 vssd1 vccd1 vccd1 _15643_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ _12855_/A _12855_/B vssd1 vssd1 vccd1 vccd1 _17461_/D sky130_fd_sc_hd__and2_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11806_ hold4022/X _13817_/B _11805_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _11806_/X
+ sky130_fd_sc_hd__o211a_1
X_18362_ _18394_/CLK hold632/X vssd1 vssd1 vccd1 vccd1 _18362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15574_ _17242_/CLK _15574_/D vssd1 vssd1 vccd1 vccd1 _15574_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _12786_/A _12786_/B vssd1 vssd1 vccd1 vccd1 _17438_/D sky130_fd_sc_hd__and2_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17313_ _17339_/CLK _17313_/D vssd1 vssd1 vccd1 vccd1 hold695/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14525_ _14596_/A _14543_/B vssd1 vssd1 vccd1 vccd1 _14525_/X sky130_fd_sc_hd__or2_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _12301_/A _11737_/B vssd1 vssd1 vccd1 vccd1 _17069_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_185_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18293_ _18325_/CLK _18293_/D vssd1 vssd1 vccd1 vccd1 _18293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14456_ hold3167/X _14481_/B _14455_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14456_/X
+ sky130_fd_sc_hd__o211a_1
X_17244_ _17244_/CLK _17244_/D vssd1 vssd1 vccd1 vccd1 _17244_/Q sky130_fd_sc_hd__dfxtp_1
X_11668_ _11762_/A _11771_/B _11667_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _11668_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13407_ _13407_/A _13407_/B vssd1 vssd1 vccd1 vccd1 _13407_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10619_ _16697_/Q _10619_/B _10619_/C vssd1 vssd1 vccd1 vccd1 _10619_/X sky130_fd_sc_hd__and3_1
X_17175_ _17281_/CLK _17175_/D vssd1 vssd1 vccd1 vccd1 _17175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14387_ _15229_/A hold2713/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14388_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11599_ hold5333/X _11789_/B _11598_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _11599_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16126_ _17321_/CLK _16126_/D vssd1 vssd1 vccd1 vccd1 hold775/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13338_ _13734_/A _13338_/B vssd1 vssd1 vccd1 vccd1 _13338_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16057_ _16093_/CLK _16057_/D vssd1 vssd1 vccd1 vccd1 hold772/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13269_ _13268_/X hold3441/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13269_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3109 _15200_/X vssd1 vssd1 vccd1 vccd1 _18382_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15008_ hold484/X hold510/A vssd1 vssd1 vccd1 vccd1 hold511/A sky130_fd_sc_hd__or2_1
XFILLER_0_196_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2408 _17961_/Q vssd1 vssd1 vccd1 vccd1 hold2408/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2419 _14039_/X vssd1 vssd1 vccd1 vccd1 _17825_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07830_ hold330/X hold355/X vssd1 vssd1 vccd1 vccd1 _07871_/B sky130_fd_sc_hd__or2_4
Xhold1707 _09288_/X vssd1 vssd1 vccd1 vccd1 _16254_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1718 _17874_/Q vssd1 vssd1 vccd1 vccd1 hold1718/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1729 _14579_/X vssd1 vssd1 vccd1 vccd1 _18083_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16959_ _17871_/CLK _16959_/D vssd1 vssd1 vccd1 vccd1 _16959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09500_ hold2177/X _16324_/Q _09992_/C vssd1 vssd1 vccd1 vccd1 _09501_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09431_ _07804_/A _09477_/B _09440_/B _09430_/X vssd1 vssd1 vccd1 vccd1 _09431_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09362_ _09362_/A _09392_/B _09362_/C _09362_/D vssd1 vssd1 vccd1 vccd1 _09369_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_59_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08313_ _15537_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08313_/X sky130_fd_sc_hd__or2_1
XFILLER_0_213_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09293_ _15515_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09293_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_11 _13116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _13180_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08244_ _14517_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08244_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_33 _13260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_44 _11774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_55 hold384/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_66 hold597/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_77 hold915/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08175_ _15509_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08175_/X sky130_fd_sc_hd__or2_1
XANTENNA_88 hold5963/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_99 _13148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5001 _11098_/X vssd1 vssd1 vccd1 vccd1 _16856_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5012 _16950_/Q vssd1 vssd1 vccd1 vccd1 hold5012/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5023 _11833_/X vssd1 vssd1 vccd1 vccd1 _17101_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5034 _17604_/Q vssd1 vssd1 vccd1 vccd1 hold5034/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4300 _17561_/Q vssd1 vssd1 vccd1 vccd1 hold4300/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5045 _11014_/X vssd1 vssd1 vccd1 vccd1 _16828_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5056 _17720_/Q vssd1 vssd1 vccd1 vccd1 hold5056/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4311 _11167_/Y vssd1 vssd1 vccd1 vccd1 _16879_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5067 _10879_/X vssd1 vssd1 vccd1 vccd1 _16783_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4322 _12379_/Y vssd1 vssd1 vccd1 vccd1 _17283_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput140 hold937/X vssd1 vssd1 vccd1 vccd1 load_status[0] sky130_fd_sc_hd__buf_12
Xhold5078 _17217_/Q vssd1 vssd1 vccd1 vccd1 hold5078/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4333 _12369_/Y vssd1 vssd1 vccd1 vccd1 _12370_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5089 _10957_/X vssd1 vssd1 vccd1 vccd1 _16809_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4344 _12312_/Y vssd1 vssd1 vccd1 vccd1 _12313_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3610 _16672_/Q vssd1 vssd1 vccd1 vccd1 hold3610/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4355 _11770_/Y vssd1 vssd1 vccd1 vccd1 _17080_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3621 _09541_/X vssd1 vssd1 vccd1 vccd1 _16337_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4366 _11779_/Y vssd1 vssd1 vccd1 vccd1 _17083_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3632 _16503_/Q vssd1 vssd1 vccd1 vccd1 hold3632/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4377 _09377_/X vssd1 vssd1 vccd1 vccd1 _16280_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3643 _10414_/X vssd1 vssd1 vccd1 vccd1 _16628_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4388 _12375_/Y vssd1 vssd1 vccd1 vccd1 _12376_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3654 _16580_/Q vssd1 vssd1 vccd1 vccd1 hold3654/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4399 _16733_/Q vssd1 vssd1 vccd1 vccd1 hold4399/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3665 _10183_/X vssd1 vssd1 vccd1 vccd1 _16551_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2920 _18188_/Q vssd1 vssd1 vccd1 vccd1 hold2920/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2931 _16179_/Q vssd1 vssd1 vccd1 vccd1 hold2931/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3676 _16657_/Q vssd1 vssd1 vccd1 vccd1 hold3676/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3687 _09976_/X vssd1 vssd1 vccd1 vccd1 _16482_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2942 _15730_/Q vssd1 vssd1 vccd1 vccd1 hold2942/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3698 _16387_/Q vssd1 vssd1 vccd1 vccd1 hold3698/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2953 _14253_/X vssd1 vssd1 vccd1 vccd1 _17927_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2964 _17817_/Q vssd1 vssd1 vccd1 vccd1 hold2964/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2975 _18013_/Q vssd1 vssd1 vccd1 vccd1 hold2975/X sky130_fd_sc_hd__dlygate4sd3_1
X_07959_ hold2760/X _07991_/A2 _07958_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _07959_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2986 _14069_/X vssd1 vssd1 vccd1 vccd1 _17839_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2997 _18002_/Q vssd1 vssd1 vccd1 vccd1 hold2997/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10970_ hold2098/X _16814_/Q _11162_/C vssd1 vssd1 vccd1 vccd1 _10971_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_214_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09629_ hold2548/X hold3218/X _10004_/C vssd1 vssd1 vccd1 vccd1 _09630_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12640_ hold1350/X hold3359/X _12844_/S vssd1 vssd1 vccd1 vccd1 _12640_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_214_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12571_ hold2846/X _17368_/Q _12970_/S vssd1 vssd1 vccd1 vccd1 _12571_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_109_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14310_ _14596_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14310_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_427_wb_clk_i clkbuf_6_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17686_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11522_ hold2079/X _16998_/Q _11717_/C vssd1 vssd1 vccd1 vccd1 _11523_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15290_ hold785/X _15448_/A2 _15446_/B1 hold790/X vssd1 vssd1 vccd1 vccd1 _15290_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14241_ hold3180/X _14268_/B _14240_/X _14372_/A vssd1 vssd1 vccd1 vccd1 _14241_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11453_ hold2779/X _16975_/Q _12323_/C vssd1 vssd1 vccd1 vccd1 _11454_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10404_ _10524_/A _10404_/B vssd1 vssd1 vccd1 vccd1 _10404_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14172_ _14457_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14172_/X sky130_fd_sc_hd__or2_1
X_11384_ hold2363/X _16952_/Q _12173_/S vssd1 vssd1 vccd1 vccd1 _11385_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_225_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13123_ _13122_/X hold5991/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13123_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_221_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10335_ _10554_/A _10335_/B vssd1 vssd1 vccd1 vccd1 _10335_/X sky130_fd_sc_hd__or2_1
XFILLER_0_221_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_237_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _17522_/Q _13056_/C _13056_/D _17523_/Q vssd1 vssd1 vccd1 vccd1 _13054_/X
+ sky130_fd_sc_hd__and4b_4
XFILLER_0_221_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17931_ _18057_/CLK _17931_/D vssd1 vssd1 vccd1 vccd1 _17931_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5590 _11698_/X vssd1 vssd1 vccd1 vccd1 _17056_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10266_ _10470_/A _10266_/B vssd1 vssd1 vccd1 vccd1 _10266_/X sky130_fd_sc_hd__or2_1
XFILLER_0_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12005_ hold2414/X _17159_/Q _13811_/C vssd1 vssd1 vccd1 vccd1 _12006_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17862_ _17862_/CLK _17862_/D vssd1 vssd1 vccd1 vccd1 _17862_/Q sky130_fd_sc_hd__dfxtp_1
X_10197_ _10530_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _10197_/X sky130_fd_sc_hd__or2_1
XFILLER_0_206_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16813_ _18016_/CLK _16813_/D vssd1 vssd1 vccd1 vccd1 _16813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17793_ _17858_/CLK _17793_/D vssd1 vssd1 vccd1 vccd1 _17793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_219_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16744_ _18045_/CLK _16744_/D vssd1 vssd1 vccd1 vccd1 _16744_/Q sky130_fd_sc_hd__dfxtp_1
X_13956_ _15517_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13956_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12907_ hold1641/X _17480_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12907_/X sky130_fd_sc_hd__mux2_1
X_16675_ _18233_/CLK _16675_/D vssd1 vssd1 vccd1 vccd1 _16675_/Q sky130_fd_sc_hd__dfxtp_1
X_13887_ hold4396/X _13407_/A _13886_/X vssd1 vssd1 vccd1 vccd1 _13887_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18414_ _18418_/CLK _18414_/D vssd1 vssd1 vccd1 vccd1 _18414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12838_ hold1921/X hold3366/X _12838_/S vssd1 vssd1 vccd1 vccd1 _12838_/X sky130_fd_sc_hd__mux2_1
X_15626_ _15886_/CLK _15626_/D vssd1 vssd1 vccd1 vccd1 _15626_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18345_ _18345_/CLK _18345_/D vssd1 vssd1 vccd1 vccd1 _18345_/Q sky130_fd_sc_hd__dfxtp_1
X_12769_ _16202_/Q hold3532/X _12838_/S vssd1 vssd1 vccd1 vccd1 _12769_/X sky130_fd_sc_hd__mux2_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15557_ _15557_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15557_/X sky130_fd_sc_hd__or2_1
XFILLER_0_189_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_168_wb_clk_i clkbuf_6_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18371_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14508_ hold1855/X _14537_/B _14507_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _14508_/X
+ sky130_fd_sc_hd__o211a_1
X_18276_ _18308_/CLK _18276_/D vssd1 vssd1 vccd1 vccd1 _18276_/Q sky130_fd_sc_hd__dfxtp_1
X_15488_ hold747/X _15488_/A2 _15485_/X vssd1 vssd1 vccd1 vccd1 _15489_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_126_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput20 hold90/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__buf_6
XFILLER_0_114_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17227_ _17259_/CLK _17227_/D vssd1 vssd1 vccd1 vccd1 _17227_/Q sky130_fd_sc_hd__dfxtp_1
Xinput31 input31/A vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14439_ _14726_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14439_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput42 input42/A vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__buf_6
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput53 input53/A vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__buf_6
Xinput64 input64/A vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_6
Xhold804 hold804/A vssd1 vssd1 vccd1 vccd1 hold804/X sky130_fd_sc_hd__dlygate4sd3_1
X_17158_ _17190_/CLK _17158_/D vssd1 vssd1 vccd1 vccd1 _17158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold815 hold815/A vssd1 vssd1 vccd1 vccd1 hold815/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold826 hold826/A vssd1 vssd1 vccd1 vccd1 hold826/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold837 hold837/A vssd1 vssd1 vccd1 vccd1 hold837/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16109_ _17336_/CLK _16109_/D vssd1 vssd1 vccd1 vccd1 hold145/A sky130_fd_sc_hd__dfxtp_1
Xhold848 hold848/A vssd1 vssd1 vccd1 vccd1 hold848/X sky130_fd_sc_hd__dlygate4sd3_1
X_09980_ hold2933/X _16484_/Q _10022_/C vssd1 vssd1 vccd1 vccd1 _09981_/B sky130_fd_sc_hd__mux2_1
X_17089_ _17843_/CLK _17089_/D vssd1 vssd1 vccd1 vccd1 _17089_/Q sky130_fd_sc_hd__dfxtp_1
Xhold859 hold859/A vssd1 vssd1 vccd1 vccd1 hold859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08931_ _15274_/A _08931_/B vssd1 vssd1 vccd1 vccd1 _16083_/D sky130_fd_sc_hd__and2_1
XFILLER_0_110_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2205 _17809_/Q vssd1 vssd1 vccd1 vccd1 hold2205/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2216 _14165_/X vssd1 vssd1 vccd1 vccd1 _17885_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08862_ hold495/X hold556/X _08866_/S vssd1 vssd1 vccd1 vccd1 hold557/A sky130_fd_sc_hd__mux2_1
Xhold2227 input67/X vssd1 vssd1 vccd1 vccd1 hold2227/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2238 _18080_/Q vssd1 vssd1 vccd1 vccd1 hold2238/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1504 _15162_/X vssd1 vssd1 vccd1 vccd1 _18364_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2249 _14181_/X vssd1 vssd1 vccd1 vccd1 _17893_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1515 _15799_/Q vssd1 vssd1 vccd1 vccd1 hold1515/X sky130_fd_sc_hd__dlygate4sd3_1
X_07813_ _14596_/A _14988_/A hold951/X _15199_/A vssd1 vssd1 vccd1 vccd1 _07813_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_58_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1526 _14215_/X vssd1 vssd1 vccd1 vccd1 _17910_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08793_ hold278/X hold602/X _08793_/S vssd1 vssd1 vccd1 vccd1 hold603/A sky130_fd_sc_hd__mux2_1
Xhold1537 _14526_/X vssd1 vssd1 vccd1 vccd1 _18059_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1548 _15841_/Q vssd1 vssd1 vccd1 vccd1 hold1548/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1559 _14135_/X vssd1 vssd1 vccd1 vccd1 _17871_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_233_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09414_ _09438_/B _16293_/Q vssd1 vssd1 vccd1 vccd1 _09414_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09345_ _15555_/A _15173_/A hold992/A _15169_/A vssd1 vssd1 vccd1 vccd1 _09359_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09276_ _12810_/A hold993/X vssd1 vssd1 vccd1 vccd1 _16249_/D sky130_fd_sc_hd__and2_1
XFILLER_0_8_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08227_ hold405/A hold337/A hold509/A hold444/A vssd1 vssd1 vccd1 vccd1 _15128_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_0_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08158_ _14164_/A hold1883/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08158_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_209_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_219_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08089_ hold2359/X _08088_/B _08088_/Y _08151_/A vssd1 vssd1 vccd1 vccd1 _08089_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4130 _13600_/X vssd1 vssd1 vccd1 vccd1 _17653_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4141 _15343_/X vssd1 vssd1 vccd1 vccd1 _15344_/B sky130_fd_sc_hd__dlygate4sd3_1
X_10120_ hold3901/X _10598_/B _10119_/X _14895_/C1 vssd1 vssd1 vccd1 vccd1 _10120_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4152 _16444_/Q vssd1 vssd1 vccd1 vccd1 hold4152/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4163 hold5956/X vssd1 vssd1 vccd1 vccd1 hold5957/A sky130_fd_sc_hd__buf_4
XFILLER_0_98_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4174 _11434_/X vssd1 vssd1 vccd1 vccd1 _16968_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3440 _10065_/Y vssd1 vssd1 vccd1 vccd1 _10066_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4185 hold5908/X vssd1 vssd1 vccd1 vccd1 hold4185/X sky130_fd_sc_hd__buf_4
XTAP_6358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10051_ _10603_/A _10051_/B vssd1 vssd1 vccd1 vccd1 _16507_/D sky130_fd_sc_hd__nor2_1
Xhold4196 _09388_/X vssd1 vssd1 vccd1 vccd1 _16282_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3451 _11202_/Y vssd1 vssd1 vccd1 vccd1 _11203_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3462 _10602_/Y vssd1 vssd1 vccd1 vccd1 _10603_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3473 _16543_/Q vssd1 vssd1 vccd1 vccd1 hold3473/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3484 _11175_/Y vssd1 vssd1 vccd1 vccd1 _11176_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2750 _08208_/X vssd1 vssd1 vccd1 vccd1 _15740_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3495 _13870_/Y vssd1 vssd1 vccd1 vccd1 _17743_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2761 _07959_/X vssd1 vssd1 vccd1 vccd1 _15622_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2772 _14081_/X vssd1 vssd1 vccd1 vccd1 _17845_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2783 _15677_/Q vssd1 vssd1 vccd1 vccd1 hold2783/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2794 _17928_/Q vssd1 vssd1 vccd1 vccd1 hold2794/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ _13819_/A _13810_/B vssd1 vssd1 vccd1 vccd1 _13810_/Y sky130_fd_sc_hd__nor2_1
X_14790_ _15183_/A _14830_/B vssd1 vssd1 vccd1 vccd1 _14790_/X sky130_fd_sc_hd__or2_1
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13741_ hold5265/X _13856_/B _13740_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13741_/X
+ sky130_fd_sc_hd__o211a_1
X_10953_ _11049_/A _10953_/B vssd1 vssd1 vccd1 vccd1 _10953_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16460_ _18242_/CLK _16460_/D vssd1 vssd1 vccd1 vccd1 _16460_/Q sky130_fd_sc_hd__dfxtp_1
X_13672_ hold3696/X _13795_/A2 _13671_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _13672_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10884_ _11655_/A _10884_/B vssd1 vssd1 vccd1 vccd1 _10884_/X sky130_fd_sc_hd__or2_1
XFILLER_0_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15411_ _16305_/Q _15477_/A2 _15487_/B1 hold853/X _15410_/X vssd1 vssd1 vccd1 vccd1
+ _15412_/D sky130_fd_sc_hd__a221o_1
X_12623_ hold3135/X _12622_/X _12851_/S vssd1 vssd1 vccd1 vccd1 _12624_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_109_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16391_ _18398_/CLK _16391_/D vssd1 vssd1 vccd1 vccd1 _16391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15342_ _15489_/A _15342_/B _15342_/C _15342_/D vssd1 vssd1 vccd1 vccd1 _15342_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_186_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18130_ _18162_/CLK _18130_/D vssd1 vssd1 vccd1 vccd1 _18130_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_261_wb_clk_i clkbuf_6_58_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18126_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12554_ hold4593/X _12553_/X _12929_/S vssd1 vssd1 vccd1 vccd1 _12555_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11505_ _12240_/A _11505_/B vssd1 vssd1 vccd1 vccd1 _11505_/X sky130_fd_sc_hd__or2_1
X_15273_ _15490_/A1 _15265_/X _15272_/X _15490_/B1 hold5927/A vssd1 vssd1 vccd1 vccd1
+ _15273_/X sky130_fd_sc_hd__a32o_1
X_18061_ _18061_/CLK _18061_/D vssd1 vssd1 vccd1 vccd1 _18061_/Q sky130_fd_sc_hd__dfxtp_1
X_12485_ hold32/X _12445_/A _12445_/B _12484_/X _15374_/A vssd1 vssd1 vccd1 vccd1
+ hold33/A sky130_fd_sc_hd__o311a_1
XFILLER_0_151_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14224_ _14974_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14224_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17012_ _17862_/CLK _17012_/D vssd1 vssd1 vccd1 vccd1 _17012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11436_ _11631_/A _11436_/B vssd1 vssd1 vccd1 vccd1 _11436_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14155_ hold2844/X _14148_/B _14154_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _14155_/X
+ sky130_fd_sc_hd__o211a_1
X_11367_ _11658_/A _11367_/B vssd1 vssd1 vccd1 vccd1 _11367_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_1332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13106_ _17564_/Q _17098_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13106_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_237_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10318_ hold3626/X _10604_/B _10317_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _10318_/X
+ sky130_fd_sc_hd__o211a_1
X_14086_ _15539_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14086_/X sky130_fd_sc_hd__or2_1
X_11298_ _12219_/A _11298_/B vssd1 vssd1 vccd1 vccd1 _11298_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13037_ _15374_/A hold908/X vssd1 vssd1 vccd1 vccd1 _17522_/D sky130_fd_sc_hd__and2_1
X_17914_ _18046_/CLK _17914_/D vssd1 vssd1 vccd1 vccd1 _17914_/Q sky130_fd_sc_hd__dfxtp_1
X_10249_ hold3814/X _10631_/B _10248_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10249_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17845_ _17883_/CLK _17845_/D vssd1 vssd1 vccd1 vccd1 _17845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17776_ _17840_/CLK _17776_/D vssd1 vssd1 vccd1 vccd1 _17776_/Q sky130_fd_sc_hd__dfxtp_1
X_14988_ _14988_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14988_/X sky130_fd_sc_hd__or2_1
XFILLER_0_135_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16727_ _18058_/CLK _16727_/D vssd1 vssd1 vccd1 vccd1 _16727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13939_ _13943_/A _13939_/B vssd1 vssd1 vccd1 vccd1 _17777_/D sky130_fd_sc_hd__and2_1
XFILLER_0_89_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_240_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_349_wb_clk_i clkbuf_6_40_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17745_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16658_ _18170_/CLK _16658_/D vssd1 vssd1 vccd1 vccd1 _16658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15609_ _18447_/CLK _15609_/D vssd1 vssd1 vccd1 vccd1 _15609_/Q sky130_fd_sc_hd__dfxtp_1
X_16589_ _18087_/CLK _16589_/D vssd1 vssd1 vccd1 vccd1 _16589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09130_ _15513_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09130_/X sky130_fd_sc_hd__or2_1
X_18328_ _18384_/CLK _18328_/D vssd1 vssd1 vccd1 vccd1 _18328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09061_ _09061_/A _09061_/B vssd1 vssd1 vccd1 vccd1 _16147_/D sky130_fd_sc_hd__and2_1
XFILLER_0_155_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18259_ _18361_/CLK _18259_/D vssd1 vssd1 vccd1 vccd1 _18259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08012_ hold2414/X _08029_/B _08011_/X _08363_/A vssd1 vssd1 vccd1 vccd1 _08012_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold601 hold601/A vssd1 vssd1 vccd1 vccd1 hold601/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold612 hold612/A vssd1 vssd1 vccd1 vccd1 hold612/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold623 hold623/A vssd1 vssd1 vccd1 vccd1 hold623/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold634 hold634/A vssd1 vssd1 vccd1 vccd1 hold634/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold645 hold645/A vssd1 vssd1 vccd1 vccd1 hold645/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold656 hold656/A vssd1 vssd1 vccd1 vccd1 hold656/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold667 hold667/A vssd1 vssd1 vccd1 vccd1 hold667/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold678 input34/X vssd1 vssd1 vccd1 vccd1 hold678/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09963_ _10563_/A _09963_/B vssd1 vssd1 vccd1 vccd1 _09963_/X sky130_fd_sc_hd__or2_1
XFILLER_0_228_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold689 hold689/A vssd1 vssd1 vccd1 vccd1 hold689/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_65_wb_clk_i clkbuf_6_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18462_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08914_ hold53/X _16075_/Q _08930_/S vssd1 vssd1 vccd1 vccd1 hold430/A sky130_fd_sc_hd__mux2_1
Xhold2002 _16162_/Q vssd1 vssd1 vccd1 vccd1 hold2002/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2013 _17998_/Q vssd1 vssd1 vccd1 vccd1 hold2013/X sky130_fd_sc_hd__dlygate4sd3_1
X_09894_ _09984_/A _09894_/B vssd1 vssd1 vccd1 vccd1 _09894_/X sky130_fd_sc_hd__or2_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2024 _13997_/X vssd1 vssd1 vccd1 vccd1 _17805_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2035 _18144_/Q vssd1 vssd1 vccd1 vccd1 hold2035/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2046 _09425_/X vssd1 vssd1 vccd1 vccd1 _16298_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1301 _16150_/Q vssd1 vssd1 vccd1 vccd1 hold1301/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _12438_/A _08845_/B vssd1 vssd1 vccd1 vccd1 _16041_/D sky130_fd_sc_hd__and2_1
XFILLER_0_209_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1312 _14831_/X vssd1 vssd1 vccd1 vccd1 _18205_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2057 _14151_/X vssd1 vssd1 vccd1 vccd1 _17879_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2068 _15626_/Q vssd1 vssd1 vccd1 vccd1 hold2068/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1323 _15598_/Q vssd1 vssd1 vccd1 vccd1 hold1323/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2079 _17846_/Q vssd1 vssd1 vccd1 vccd1 hold2079/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1334 _16200_/Q vssd1 vssd1 vccd1 vccd1 hold1334/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1345 _07983_/X vssd1 vssd1 vccd1 vccd1 _15634_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_1361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1356 _15584_/Q vssd1 vssd1 vccd1 vccd1 hold1356/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08776_ _15394_/A _08776_/B vssd1 vssd1 vccd1 vccd1 _16008_/D sky130_fd_sc_hd__and2_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1367 hold910/X vssd1 vssd1 vccd1 vccd1 hold1367/X sky130_fd_sc_hd__buf_8
Xhold1378 _15865_/Q vssd1 vssd1 vccd1 vccd1 hold1378/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1389 hold6049/X vssd1 vssd1 vccd1 vccd1 input2/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09328_ hold1552/X _09325_/B _09327_/X _12597_/A vssd1 vssd1 vccd1 vccd1 _09328_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09259_ _09313_/A _16241_/Q _09283_/S vssd1 vssd1 vccd1 vccd1 _09259_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _13749_/A _12270_/B vssd1 vssd1 vccd1 vccd1 _12270_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11221_ _12331_/A _11221_/B vssd1 vssd1 vccd1 vccd1 _11221_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_142_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11152_ _12301_/A _11152_/B vssd1 vssd1 vccd1 vccd1 _16874_/D sky130_fd_sc_hd__nor2_1
XTAP_6111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10103_ hold1728/X hold3501/X _10595_/C vssd1 vssd1 vccd1 vccd1 _10104_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_235_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15960_ _17322_/CLK _15960_/D vssd1 vssd1 vccd1 vccd1 hold323/A sky130_fd_sc_hd__dfxtp_1
XTAP_5410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11083_ hold5173/X _11204_/B _11082_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _11083_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3270 _16385_/Q vssd1 vssd1 vccd1 vccd1 hold3270/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3281 _10339_/X vssd1 vssd1 vccd1 vccd1 _16603_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10034_ _16502_/Q _10052_/B _10040_/C vssd1 vssd1 vccd1 vccd1 _10034_/X sky130_fd_sc_hd__and3_1
X_14911_ hold2497/X _14896_/Y _14910_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _14911_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3292 _16585_/Q vssd1 vssd1 vccd1 vccd1 hold3292/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15891_ _18412_/CLK _15891_/D vssd1 vssd1 vccd1 vccd1 hold741/A sky130_fd_sc_hd__dfxtp_1
XTAP_5465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2580 _16171_/Q vssd1 vssd1 vccd1 vccd1 hold2580/X sky130_fd_sc_hd__dlygate4sd3_1
X_17630_ _17630_/CLK _17630_/D vssd1 vssd1 vccd1 vccd1 _17630_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ hold330/X _14843_/B vssd1 vssd1 vccd1 vccd1 hold331/A sky130_fd_sc_hd__nor2_1
Xhold2591 _15838_/Q vssd1 vssd1 vccd1 vccd1 hold2591/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1890 _14657_/X vssd1 vssd1 vccd1 vccd1 _18121_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17561_ _17561_/CLK _17561_/D vssd1 vssd1 vccd1 vccd1 _17561_/Q sky130_fd_sc_hd__dfxtp_1
X_14773_ hold2544/X _14772_/B _14772_/Y _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14773_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11985_ _13407_/A _11985_/B vssd1 vssd1 vccd1 vccd1 _11985_/X sky130_fd_sc_hd__or2_1
XFILLER_0_203_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16512_ _18265_/CLK _16512_/D vssd1 vssd1 vccd1 vccd1 _16512_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_442_wb_clk_i clkbuf_6_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17719_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13724_ hold1532/X hold4589/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13725_/B sky130_fd_sc_hd__mux2_1
X_10936_ hold4817/X _11789_/B _10935_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _10936_/X
+ sky130_fd_sc_hd__o211a_1
X_17492_ _17492_/CLK _17492_/D vssd1 vssd1 vccd1 vccd1 _17492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16443_ _18388_/CLK _16443_/D vssd1 vssd1 vccd1 vccd1 _16443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10867_ hold4972/X _11153_/B _10866_/X _14552_/C1 vssd1 vssd1 vccd1 vccd1 _10867_/X
+ sky130_fd_sc_hd__o211a_1
X_13655_ hold2687/X _17672_/Q _13841_/C vssd1 vssd1 vccd1 vccd1 _13656_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12606_ _12612_/A _12606_/B vssd1 vssd1 vccd1 vccd1 _17378_/D sky130_fd_sc_hd__and2_1
XFILLER_0_184_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16374_ _18325_/CLK _16374_/D vssd1 vssd1 vccd1 vccd1 _16374_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ hold2956/X hold5394/X _13874_/C vssd1 vssd1 vccd1 vccd1 _13587_/B sky130_fd_sc_hd__mux2_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ hold5131/X _11186_/B _10797_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10798_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18113_ _18262_/CLK _18113_/D vssd1 vssd1 vccd1 vccd1 _18113_/Q sky130_fd_sc_hd__dfxtp_1
X_15325_ hold563/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15325_/X sky130_fd_sc_hd__or2_1
X_12537_ _12948_/A _12537_/B vssd1 vssd1 vccd1 vccd1 _17355_/D sky130_fd_sc_hd__and2_1
XFILLER_0_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18044_ _18047_/CLK _18044_/D vssd1 vssd1 vccd1 vccd1 _18044_/Q sky130_fd_sc_hd__dfxtp_1
X_12468_ _17327_/Q _12506_/B vssd1 vssd1 vccd1 vccd1 _12468_/X sky130_fd_sc_hd__or2_1
X_15256_ _17329_/Q _09362_/C _15485_/B1 hold398/X vssd1 vssd1 vccd1 vccd1 _15256_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_227_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14207_ hold1285/X _14202_/B _14206_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _14207_/X
+ sky130_fd_sc_hd__o211a_1
X_11419_ hold4161/X _11792_/B _11418_/X _14143_/C1 vssd1 vssd1 vccd1 vccd1 _11419_/X
+ sky130_fd_sc_hd__o211a_1
X_15187_ _15187_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15187_/X sky130_fd_sc_hd__or2_1
X_12399_ hold673/X hold810/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold811/A sky130_fd_sc_hd__mux2_1
XFILLER_0_240_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14138_ _14477_/A _14140_/B vssd1 vssd1 vccd1 vccd1 _14138_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14069_ hold2985/X _14107_/A2 _14068_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _14069_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08630_ _12390_/A hold526/X vssd1 vssd1 vccd1 vccd1 _15937_/D sky130_fd_sc_hd__and2_1
XFILLER_0_158_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17828_ _18060_/CLK _17828_/D vssd1 vssd1 vccd1 vccd1 _17828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08561_ _15434_/A _08561_/B vssd1 vssd1 vccd1 vccd1 _15904_/D sky130_fd_sc_hd__and2_1
XFILLER_0_222_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17759_ _17825_/CLK _17759_/D vssd1 vssd1 vccd1 vccd1 _17759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_183_wb_clk_i clkbuf_6_54_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18265_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08492_ _14330_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08492_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_112_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17523_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_147_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09113_ hold2580/X _09106_/B _09112_/X _12948_/A vssd1 vssd1 vccd1 vccd1 _09113_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09044_ hold53/X hold759/X _09060_/S vssd1 vssd1 vccd1 vccd1 _09045_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_115_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold420 hold420/A vssd1 vssd1 vccd1 vccd1 hold420/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 hold431/A vssd1 vssd1 vccd1 vccd1 hold431/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold442 hold442/A vssd1 vssd1 vccd1 vccd1 input55/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 hold453/A vssd1 vssd1 vccd1 vccd1 hold453/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold464 hold464/A vssd1 vssd1 vccd1 vccd1 hold464/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 hold475/A vssd1 vssd1 vccd1 vccd1 hold475/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 hold486/A vssd1 vssd1 vccd1 vccd1 hold486/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout900 _14972_/A vssd1 vssd1 vccd1 vccd1 _15513_/A sky130_fd_sc_hd__clkbuf_16
Xhold497 hold497/A vssd1 vssd1 vccd1 vccd1 hold497/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout911 _14960_/A vssd1 vssd1 vccd1 vccd1 _15229_/A sky130_fd_sc_hd__buf_8
XFILLER_0_217_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout922 hold484/X vssd1 vssd1 vccd1 vccd1 _15169_/A sky130_fd_sc_hd__clkbuf_16
X_09946_ hold5185/X _11204_/B _09945_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _09946_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout933 hold1183/X vssd1 vssd1 vccd1 vccd1 _15535_/A sky130_fd_sc_hd__buf_6
Xfanout944 hold1106/X vssd1 vssd1 vccd1 vccd1 hold1107/A sky130_fd_sc_hd__buf_6
XFILLER_0_216_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ hold3266/X _10067_/B _09876_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09877_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1120 _07795_/X vssd1 vssd1 vccd1 vccd1 _07796_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 _09137_/X vssd1 vssd1 vccd1 vccd1 _16181_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 _08241_/X vssd1 vssd1 vccd1 vccd1 _15755_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ hold77/X hold292/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08829_/B sky130_fd_sc_hd__mux2_1
Xhold1153 input38/X vssd1 vssd1 vccd1 vccd1 hold1153/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 _09079_/X vssd1 vssd1 vccd1 vccd1 _16154_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1175 _15749_/Q vssd1 vssd1 vccd1 vccd1 hold1175/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 _16183_/Q vssd1 vssd1 vccd1 vccd1 hold1186/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ hold172/X hold877/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08760_/B sky130_fd_sc_hd__mux2_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1197 _13916_/X vssd1 vssd1 vccd1 vccd1 _13917_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11770_ _12337_/A _11770_/B vssd1 vssd1 vccd1 vccd1 _11770_/Y sky130_fd_sc_hd__nor2_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10721_ hold2995/X hold3450/X _11201_/C vssd1 vssd1 vccd1 vccd1 _10722_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13440_ _13737_/A _13440_/B vssd1 vssd1 vccd1 vccd1 _13440_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10652_ hold2119/X _16708_/Q _11723_/C vssd1 vssd1 vccd1 vccd1 _10653_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_193_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13371_ _13791_/A _13371_/B vssd1 vssd1 vccd1 vccd1 _13371_/X sky130_fd_sc_hd__or2_1
X_10583_ _16685_/Q _10619_/B _10595_/C vssd1 vssd1 vccd1 vccd1 _10583_/X sky130_fd_sc_hd__and3_1
XFILLER_0_23_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15110_ hold2631/X hold340/X _15109_/Y _15176_/C1 vssd1 vssd1 vccd1 vccd1 _15110_/X
+ sky130_fd_sc_hd__o211a_1
X_12322_ _13819_/A _12322_/B vssd1 vssd1 vccd1 vccd1 _17264_/D sky130_fd_sc_hd__nor2_1
X_16090_ _16090_/CLK _16090_/D vssd1 vssd1 vccd1 vccd1 hold796/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15041_ _14988_/A hold2561/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15042_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12253_ hold5759/X _12362_/B _12252_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _12253_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11204_ _16892_/Q _11204_/B _11204_/C vssd1 vssd1 vccd1 vccd1 _11204_/X sky130_fd_sc_hd__and3_1
XFILLER_0_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12184_ hold5175/X _12374_/B _12183_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _12184_/X
+ sky130_fd_sc_hd__o211a_1
X_11135_ hold1893/X _16869_/Q _11153_/C vssd1 vssd1 vccd1 vccd1 _11136_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_101_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16992_ _17840_/CLK _16992_/D vssd1 vssd1 vccd1 vccd1 _16992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15943_ _17337_/CLK _15943_/D vssd1 vssd1 vccd1 vccd1 hold497/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11066_ hold2195/X hold4727/X _11162_/C vssd1 vssd1 vccd1 vccd1 _11067_/B sky130_fd_sc_hd__mux2_1
XTAP_5251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10017_ _13158_/A _09981_/A _10016_/X vssd1 vssd1 vccd1 vccd1 _10017_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ _17187_/CLK _15874_/D vssd1 vssd1 vccd1 vccd1 _15874_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17613_ _17709_/CLK _17613_/D vssd1 vssd1 vccd1 vccd1 _17613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ hold2376/X _14828_/B _14824_/Y _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14825_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_231_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ _18392_/CLK _17544_/D vssd1 vssd1 vccd1 vccd1 _17544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14756_ _14988_/A _14780_/B vssd1 vssd1 vccd1 vccd1 _14756_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11968_ hold5791/X _12350_/B _11967_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _11968_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13707_ _13722_/A _13707_/B vssd1 vssd1 vccd1 vccd1 _13707_/X sky130_fd_sc_hd__or2_1
X_17475_ _17476_/CLK _17475_/D vssd1 vssd1 vccd1 vccd1 _17475_/Q sky130_fd_sc_hd__dfxtp_1
X_10919_ hold2392/X _16797_/Q _11789_/C vssd1 vssd1 vccd1 vccd1 _10920_/B sky130_fd_sc_hd__mux2_1
X_14687_ hold1700/X _14720_/B _14686_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14687_/X
+ sky130_fd_sc_hd__o211a_1
X_11899_ hold4966/X _13886_/B _11898_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _11899_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16426_ _18371_/CLK _16426_/D vssd1 vssd1 vccd1 vccd1 _16426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13638_ _13734_/A _13638_/B vssd1 vssd1 vccd1 vccd1 _13638_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16357_ _18423_/CLK _16357_/D vssd1 vssd1 vccd1 vccd1 _16357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13569_ _13752_/A _13569_/B vssd1 vssd1 vccd1 vccd1 _13569_/X sky130_fd_sc_hd__or2_1
XFILLER_0_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6109 la_data_in[13] vssd1 vssd1 vccd1 vccd1 hold6109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15308_ hold793/X _09386_/A _15441_/A2 hold888/X vssd1 vssd1 vccd1 vccd1 _15308_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16288_ _16315_/CLK _16288_/D vssd1 vssd1 vccd1 vccd1 _16288_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5408 _17076_/Q vssd1 vssd1 vccd1 vccd1 hold5408/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_152_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5419 _13402_/X vssd1 vssd1 vccd1 vccd1 _17587_/D sky130_fd_sc_hd__dlygate4sd3_1
X_18027_ _18059_/CLK _18027_/D vssd1 vssd1 vccd1 vccd1 _18027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15239_ hold414/X _15485_/A2 _15488_/A2 hold837/X _15238_/X vssd1 vssd1 vccd1 vccd1
+ _15242_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_151_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4707 _16505_/Q vssd1 vssd1 vccd1 vccd1 hold4707/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4718 _11772_/Y vssd1 vssd1 vccd1 vccd1 _11773_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4729 _16877_/Q vssd1 vssd1 vccd1 vccd1 hold4729/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09800_ _18337_/Q _16424_/Q _09992_/C vssd1 vssd1 vccd1 vccd1 _09801_/B sky130_fd_sc_hd__mux2_1
Xfanout207 _11222_/B vssd1 vssd1 vccd1 vccd1 _11765_/B sky130_fd_sc_hd__buf_4
Xfanout218 _10004_/B vssd1 vssd1 vccd1 vccd1 _10028_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout229 _10616_/B vssd1 vssd1 vccd1 vccd1 _11225_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07992_ hold337/X hold509/X hold444/X hold405/X vssd1 vssd1 vccd1 vccd1 _09498_/A
+ sky130_fd_sc_hd__nand4b_4
XFILLER_0_238_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09731_ hold788/X _16401_/Q _10067_/C vssd1 vssd1 vccd1 vccd1 _09732_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09662_ hold2081/X hold3678/X _10067_/C vssd1 vssd1 vccd1 vccd1 _09663_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_364_wb_clk_i clkbuf_6_34_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17744_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_206_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08613_ hold679/X hold777/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold778/A sky130_fd_sc_hd__mux2_1
XFILLER_0_222_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09593_ _18268_/Q _13310_/A _10601_/C vssd1 vssd1 vccd1 vccd1 _09594_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08544_ hold29/X _15896_/Q _08544_/S vssd1 vssd1 vccd1 vccd1 hold197/A sky130_fd_sc_hd__mux2_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08475_ hold1380/X _08486_/B _08474_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _08475_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_6_9_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_9_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_80_wb_clk_i clkbuf_6_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17517_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09027_ _12420_/A hold345/X vssd1 vssd1 vccd1 vccd1 _16130_/D sky130_fd_sc_hd__and2_1
XFILLER_0_61_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5920 hold5920/A vssd1 vssd1 vccd1 vccd1 hold5920/X sky130_fd_sc_hd__buf_2
Xhold5931 hold5931/A vssd1 vssd1 vccd1 vccd1 hold5931/X sky130_fd_sc_hd__clkbuf_4
Xhold5942 hold6111/X vssd1 vssd1 vccd1 vccd1 hold907/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_103_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5953 hold6022/X vssd1 vssd1 vccd1 vccd1 _17754_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5964 _18420_/Q vssd1 vssd1 vccd1 vccd1 hold5964/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold250 hold250/A vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5975 hold6105/X vssd1 vssd1 vccd1 vccd1 _18463_/A sky130_fd_sc_hd__clkbuf_2
Xhold261 hold261/A vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5986 hold6133/X vssd1 vssd1 vccd1 vccd1 _09447_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold5997 _13149_/X vssd1 vssd1 vccd1 vccd1 hold5997/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 hold272/A vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 hold283/A vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 hold360/X vssd1 vssd1 vccd1 vccd1 hold361/A sky130_fd_sc_hd__buf_4
Xfanout730 _09003_/A vssd1 vssd1 vccd1 vccd1 _15434_/A sky130_fd_sc_hd__clkbuf_4
Xfanout741 _13675_/C1 vssd1 vssd1 vccd1 vccd1 _13729_/C1 sky130_fd_sc_hd__buf_2
XFILLER_0_217_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09929_ hold1857/X hold4606/X _10031_/C vssd1 vssd1 vccd1 vccd1 _09930_/B sky130_fd_sc_hd__mux2_1
Xfanout752 fanout843/X vssd1 vssd1 vccd1 vccd1 _08119_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout763 _14131_/C1 vssd1 vssd1 vccd1 vccd1 _14528_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout774 fanout791/X vssd1 vssd1 vccd1 vccd1 _08385_/A sky130_fd_sc_hd__buf_4
Xfanout785 _14143_/C1 vssd1 vssd1 vccd1 vccd1 _08125_/A sky130_fd_sc_hd__buf_4
XFILLER_0_226_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout796 _15054_/A vssd1 vssd1 vccd1 vccd1 _15068_/A sky130_fd_sc_hd__buf_4
XFILLER_0_198_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12940_ hold1163/X _17491_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12940_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_137_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12871_ hold3057/X _17468_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _12871_/X sky130_fd_sc_hd__mux2_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_101 _17571_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 _14988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _15165_/A _14610_/B vssd1 vssd1 vccd1 vccd1 _14610_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_123 hold1367/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11822_ hold2645/X hold4361/X _13811_/C vssd1 vssd1 vccd1 vccd1 _11823_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _17898_/CLK _15590_/D vssd1 vssd1 vccd1 vccd1 _15590_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14541_ _15221_/A _14541_/B vssd1 vssd1 vccd1 vccd1 _14541_/Y sky130_fd_sc_hd__nand2_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _17075_/Q _11753_/B _11753_/C vssd1 vssd1 vccd1 vccd1 _11753_/X sky130_fd_sc_hd__and3_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10704_ _11121_/A _10704_/B vssd1 vssd1 vccd1 vccd1 _10704_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _17260_/CLK _17260_/D vssd1 vssd1 vccd1 vccd1 _17260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14472_ hold1523/X _14481_/B _14471_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _14472_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ hold1484/X _17052_/Q _12323_/C vssd1 vssd1 vccd1 vccd1 _11685_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16211_ _17445_/CLK hold968/X vssd1 vssd1 vccd1 vccd1 _16211_/Q sky130_fd_sc_hd__dfxtp_1
X_10635_ hold3441/X _10563_/A _10634_/X vssd1 vssd1 vccd1 vccd1 _10636_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13423_ hold4066/X _13817_/B _13422_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _13423_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17191_ _17194_/CLK _17191_/D vssd1 vssd1 vccd1 vccd1 _17191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16142_ _18412_/CLK _16142_/D vssd1 vssd1 vccd1 vccd1 hold575/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13354_ hold3838/X _13862_/B _13353_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13354_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10566_ hold3417/X _10476_/A _10565_/X vssd1 vssd1 vccd1 vccd1 _10567_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12305_ _17259_/Q _12305_/B _12305_/C vssd1 vssd1 vccd1 vccd1 _12305_/X sky130_fd_sc_hd__and3_1
X_16073_ _17322_/CLK _16073_/D vssd1 vssd1 vccd1 vccd1 hold283/A sky130_fd_sc_hd__dfxtp_1
X_13285_ _13284_/X hold3459/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13285_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_133_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10497_ _10563_/A _10497_/B vssd1 vssd1 vccd1 vccd1 _10497_/X sky130_fd_sc_hd__or2_1
X_15024_ _15024_/A _15024_/B vssd1 vssd1 vccd1 vccd1 _18297_/D sky130_fd_sc_hd__and2_1
X_12236_ hold1039/X hold4563/X _12332_/C vssd1 vssd1 vccd1 vccd1 _12237_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_236_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12167_ hold2567/X hold4480/X _12362_/C vssd1 vssd1 vccd1 vccd1 _12168_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_209_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11118_ _11121_/A _11118_/B vssd1 vssd1 vccd1 vccd1 _11118_/X sky130_fd_sc_hd__or2_1
XFILLER_0_208_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12098_ hold2068/X _17190_/Q _13796_/S vssd1 vssd1 vccd1 vccd1 _12099_/B sky130_fd_sc_hd__mux2_1
X_16975_ _17823_/CLK _16975_/D vssd1 vssd1 vccd1 vccd1 _16975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15926_ _17288_/CLK _15926_/D vssd1 vssd1 vccd1 vccd1 hold829/A sky130_fd_sc_hd__dfxtp_1
X_11049_ _11049_/A _11049_/B vssd1 vssd1 vccd1 vccd1 _11049_/X sky130_fd_sc_hd__or2_1
Xinput7 input7/A vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_6
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ _17678_/CLK _15857_/D vssd1 vssd1 vccd1 vccd1 _15857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_231_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14808_ _15201_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14808_/X sky130_fd_sc_hd__or2_1
XFILLER_0_235_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15788_ _17720_/CLK _15788_/D vssd1 vssd1 vccd1 vccd1 _15788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17527_ _17533_/CLK _17527_/D vssd1 vssd1 vccd1 vccd1 _17527_/Q sky130_fd_sc_hd__dfxtp_1
X_14739_ hold1972/X _14772_/B _14738_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14739_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_188_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08260_ _14604_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08260_/X sky130_fd_sc_hd__or2_1
X_17458_ _18458_/CLK _17458_/D vssd1 vssd1 vccd1 vccd1 _17458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16409_ _18386_/CLK _16409_/D vssd1 vssd1 vccd1 vccd1 _16409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08191_ _15145_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08191_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17389_ _18455_/CLK _17389_/D vssd1 vssd1 vccd1 vccd1 _17389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5205 _16847_/Q vssd1 vssd1 vccd1 vccd1 hold5205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5216 _10780_/X vssd1 vssd1 vccd1 vccd1 _16750_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5227 _16768_/Q vssd1 vssd1 vccd1 vccd1 hold5227/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5238 _12088_/X vssd1 vssd1 vccd1 vccd1 _17186_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4504 _16596_/Q vssd1 vssd1 vccd1 vccd1 hold4504/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5249 _17614_/Q vssd1 vssd1 vccd1 vccd1 hold5249/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4515 _13881_/Y vssd1 vssd1 vccd1 vccd1 _13882_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4526 _10348_/X vssd1 vssd1 vccd1 vccd1 _16606_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4537 _16574_/Q vssd1 vssd1 vccd1 vccd1 hold4537/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3803 _16607_/Q vssd1 vssd1 vccd1 vccd1 hold3803/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4548 _09838_/X vssd1 vssd1 vccd1 vccd1 _16436_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3814 _16605_/Q vssd1 vssd1 vccd1 vccd1 hold3814/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4559 _17634_/Q vssd1 vssd1 vccd1 vccd1 hold4559/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3825 _10843_/X vssd1 vssd1 vccd1 vccd1 _16771_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3836 _16839_/Q vssd1 vssd1 vccd1 vccd1 hold3836/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3847 _10276_/X vssd1 vssd1 vccd1 vccd1 _16582_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3858 _16865_/Q vssd1 vssd1 vccd1 vccd1 hold3858/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3869 _11047_/X vssd1 vssd1 vccd1 vccd1 _16839_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07975_ hold2648/X _07978_/B _07974_/Y _12103_/C1 vssd1 vssd1 vccd1 vccd1 _07975_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09714_ _09912_/A _09714_/B vssd1 vssd1 vccd1 vccd1 _09714_/X sky130_fd_sc_hd__or2_1
XFILLER_0_208_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09645_ _09933_/A _09645_/B vssd1 vssd1 vccd1 vccd1 _09645_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09576_ _10482_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09576_/X sky130_fd_sc_hd__or2_1
XFILLER_0_139_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _12410_/A hold814/X vssd1 vssd1 vccd1 vccd1 _15888_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_9_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_212_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08458_ _15517_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08458_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_212_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08389_ _08389_/A _08389_/B vssd1 vssd1 vccd1 vccd1 _15826_/D sky130_fd_sc_hd__and2_1
XFILLER_0_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10420_ hold4452/X _10628_/B _10419_/X _14697_/C1 vssd1 vssd1 vccd1 vccd1 _10420_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10351_ hold3785/X _10631_/B _10350_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10351_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13070_ _13070_/A _13294_/B vssd1 vssd1 vccd1 vccd1 _13070_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5750 _11950_/X vssd1 vssd1 vccd1 vccd1 _17140_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10282_ hold3915/X _10568_/B _10281_/X _14769_/C1 vssd1 vssd1 vccd1 vccd1 _10282_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5761 _17278_/Q vssd1 vssd1 vccd1 vccd1 hold5761/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5772 _12172_/X vssd1 vssd1 vccd1 vccd1 _17214_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5783 _17722_/Q vssd1 vssd1 vccd1 vccd1 hold5783/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12021_ _13797_/A _12021_/B vssd1 vssd1 vccd1 vccd1 _12021_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_286_wb_clk_i clkbuf_6_48_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18054_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5794 _12256_/X vssd1 vssd1 vccd1 vccd1 _17242_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_215_wb_clk_i clkbuf_6_60_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18203_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_228_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout560 hold107/X vssd1 vssd1 vccd1 vccd1 _08152_/S sky130_fd_sc_hd__clkbuf_8
Xfanout571 _07884_/Y vssd1 vssd1 vccd1 vccd1 _07924_/B sky130_fd_sc_hd__buf_8
XFILLER_0_79_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16760_ _18057_/CLK _16760_/D vssd1 vssd1 vccd1 vccd1 _16760_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout582 _13057_/X vssd1 vssd1 vccd1 vccd1 _13306_/S sky130_fd_sc_hd__clkbuf_16
Xfanout593 _12871_/S vssd1 vssd1 vccd1 vccd1 _12811_/S sky130_fd_sc_hd__buf_6
X_13972_ _15207_/A _13994_/B vssd1 vssd1 vccd1 vccd1 _13972_/X sky130_fd_sc_hd__or2_1
X_15711_ _17281_/CLK _15711_/D vssd1 vssd1 vccd1 vccd1 _15711_/Q sky130_fd_sc_hd__dfxtp_1
X_12923_ hold3314/X _12922_/X _12923_/S vssd1 vssd1 vccd1 vccd1 _12923_/X sky130_fd_sc_hd__mux2_1
X_16691_ _18217_/CLK _16691_/D vssd1 vssd1 vccd1 vccd1 _16691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18430_ _18430_/CLK _18430_/D vssd1 vssd1 vccd1 vccd1 _18430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15642_ _17154_/CLK _15642_/D vssd1 vssd1 vccd1 vccd1 _15642_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ hold3349/X _12853_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12855_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_87_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18361_ _18361_/CLK _18361_/D vssd1 vssd1 vccd1 vccd1 _18361_/Q sky130_fd_sc_hd__dfxtp_1
X_11805_ _13800_/A _11805_/B vssd1 vssd1 vccd1 vccd1 _11805_/X sky130_fd_sc_hd__or2_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15573_ _17743_/CLK _15573_/D vssd1 vssd1 vccd1 vccd1 _15573_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12785_ hold3619/X _12784_/X _12839_/S vssd1 vssd1 vccd1 vccd1 _12786_/B sky130_fd_sc_hd__mux2_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17312_ _17336_/CLK _17312_/D vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__dfxtp_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14524_ hold2781/X _14537_/B _14523_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _14524_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18292_ _18346_/CLK _18292_/D vssd1 vssd1 vccd1 vccd1 _18292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11736_ hold4636/X _11649_/A _11735_/X vssd1 vssd1 vccd1 vccd1 _11736_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17243_ _17741_/CLK _17243_/D vssd1 vssd1 vccd1 vccd1 _17243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14455_ _15189_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14455_/X sky130_fd_sc_hd__or2_1
X_11667_ _11667_/A _11667_/B vssd1 vssd1 vccd1 vccd1 _11667_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13406_ hold1188/X hold4396/X _13886_/C vssd1 vssd1 vccd1 vccd1 _13407_/B sky130_fd_sc_hd__mux2_1
X_10618_ _11206_/A _10618_/B vssd1 vssd1 vccd1 vccd1 _16696_/D sky130_fd_sc_hd__nor2_1
X_17174_ _17898_/CLK _17174_/D vssd1 vssd1 vccd1 vccd1 _17174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14386_ _14390_/A _14386_/B vssd1 vssd1 vccd1 vccd1 _17992_/D sky130_fd_sc_hd__and2_1
X_11598_ _11694_/A _11598_/B vssd1 vssd1 vccd1 vccd1 _11598_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16125_ _16125_/CLK _16125_/D vssd1 vssd1 vccd1 vccd1 hold876/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10549_ hold4571/X _10646_/B _10548_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10549_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13337_ hold1395/X hold4335/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13338_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_40_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16056_ _17291_/CLK _16056_/D vssd1 vssd1 vccd1 vccd1 hold874/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13268_ hold3512/X _13267_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13268_/X sky130_fd_sc_hd__mux2_2
X_15007_ hold2424/X hold447/X _15006_/Y _15072_/A vssd1 vssd1 vccd1 vccd1 _15007_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_1324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12219_ _12219_/A _12219_/B vssd1 vssd1 vccd1 vccd1 _12219_/X sky130_fd_sc_hd__or2_1
X_13199_ _13199_/A1 _13197_/X _13198_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13199_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2409 _14323_/X vssd1 vssd1 vccd1 vccd1 _17961_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1708 _16226_/Q vssd1 vssd1 vccd1 vccd1 hold1708/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1719 _14141_/X vssd1 vssd1 vccd1 vccd1 _17874_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16958_ _17774_/CLK _16958_/D vssd1 vssd1 vccd1 vccd1 _16958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15909_ _17284_/CLK _15909_/D vssd1 vssd1 vccd1 vccd1 hold582/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16889_ _18060_/CLK _16889_/D vssd1 vssd1 vccd1 vccd1 _16889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09430_ _09438_/B _16301_/Q vssd1 vssd1 vccd1 vccd1 _09430_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09361_ _09366_/A _09364_/B _09361_/C vssd1 vssd1 vccd1 vccd1 _09361_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_19_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08312_ hold1841/X _08323_/B _08311_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _08312_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_19_wb_clk_i clkbuf_6_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17464_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_129_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09292_ hold1473/X _09325_/B _09291_/X _12948_/A vssd1 vssd1 vccd1 vccd1 _09292_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 _13116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_23 _13180_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ hold2946/X _08268_/B _08242_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08243_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_34 _13260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_45 _15056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_56 hold235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_67 hold597/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_78 hold951/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08174_ _08504_/A _15182_/A vssd1 vssd1 vccd1 vccd1 _08215_/B sky130_fd_sc_hd__or2_4
XFILLER_0_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_89 hold5957/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5002 _17035_/Q vssd1 vssd1 vccd1 vccd1 hold5002/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5013 _11284_/X vssd1 vssd1 vccd1 vccd1 _16918_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5024 _17694_/Q vssd1 vssd1 vccd1 vccd1 hold5024/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5035 _13357_/X vssd1 vssd1 vccd1 vccd1 _17572_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4301 _13803_/Y vssd1 vssd1 vccd1 vccd1 _13804_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5046 _17636_/Q vssd1 vssd1 vccd1 vccd1 hold5046/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5057 _13705_/X vssd1 vssd1 vccd1 vccd1 _17688_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4312 _16914_/Q vssd1 vssd1 vccd1 vccd1 hold4312/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4323 _17096_/Q vssd1 vssd1 vccd1 vccd1 hold4323/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput130 hold5963/X vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_12
Xhold5068 _17092_/Q vssd1 vssd1 vccd1 vccd1 hold5068/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput141 hold5909/X vssd1 vssd1 vccd1 vccd1 hold5910/A sky130_fd_sc_hd__buf_6
Xhold5079 _12085_/X vssd1 vssd1 vccd1 vccd1 _17185_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4334 _12370_/Y vssd1 vssd1 vccd1 vccd1 _17280_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3600 _12557_/X vssd1 vssd1 vccd1 vccd1 _12558_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4345 _16907_/Q vssd1 vssd1 vccd1 vccd1 hold4345/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3611 _10450_/X vssd1 vssd1 vccd1 vccd1 _16640_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4356 _16736_/Q vssd1 vssd1 vccd1 vccd1 hold4356/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3622 _16376_/Q vssd1 vssd1 vccd1 vccd1 hold3622/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4367 _17584_/Q vssd1 vssd1 vccd1 vccd1 hold4367/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3633 _09943_/X vssd1 vssd1 vccd1 vccd1 _16471_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4378 _17572_/Q vssd1 vssd1 vccd1 vccd1 hold4378/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3644 _16556_/Q vssd1 vssd1 vccd1 vccd1 hold3644/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4389 _12376_/Y vssd1 vssd1 vccd1 vccd1 _17282_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3655 _10174_/X vssd1 vssd1 vccd1 vccd1 _16548_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2910 _15619_/Q vssd1 vssd1 vccd1 vccd1 hold2910/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3666 _16652_/Q vssd1 vssd1 vccd1 vccd1 hold3666/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2921 _14797_/X vssd1 vssd1 vccd1 vccd1 _18188_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3677 _10405_/X vssd1 vssd1 vccd1 vccd1 _16625_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2932 _09133_/X vssd1 vssd1 vccd1 vccd1 _16179_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3688 _16584_/Q vssd1 vssd1 vccd1 vccd1 hold3688/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2943 _08188_/X vssd1 vssd1 vccd1 vccd1 _15730_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2954 _16218_/Q vssd1 vssd1 vccd1 vccd1 hold2954/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3699 _09595_/X vssd1 vssd1 vccd1 vccd1 _16355_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2965 _14023_/X vssd1 vssd1 vccd1 vccd1 _17817_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2976 _14430_/X vssd1 vssd1 vccd1 vccd1 _18013_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07958_ _14413_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07958_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2987 _15830_/Q vssd1 vssd1 vccd1 vccd1 hold2987/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2998 _14408_/X vssd1 vssd1 vccd1 vccd1 _18002_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07889_ hold1574/X _07924_/B _07888_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _07889_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09628_ hold4145/X _11201_/B _09627_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09628_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09559_ hold3224/X _10577_/B _09558_/X _15204_/C1 vssd1 vssd1 vccd1 vccd1 _09559_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12570_ _14358_/A _12570_/B vssd1 vssd1 vccd1 vccd1 _17366_/D sky130_fd_sc_hd__and2_1
XFILLER_0_66_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11521_ hold4083/X _12305_/B _11520_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _11521_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14240_ _15189_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14240_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11452_ hold5474/X _11165_/B _11451_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _11452_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10403_ hold1598/X _16625_/Q _10595_/C vssd1 vssd1 vccd1 vccd1 _10404_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_151_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14171_ hold6055/X _14198_/B hold1581/X _14352_/A vssd1 vssd1 vccd1 vccd1 _14171_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11383_ hold5183/X _11765_/B _11382_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _11383_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10334_ hold1972/X _16602_/Q _10640_/C vssd1 vssd1 vccd1 vccd1 _10335_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13122_ _17566_/Q _17100_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13122_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_225_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13053_ hold907/A _13056_/C _13055_/C _17523_/Q vssd1 vssd1 vccd1 vccd1 _13310_/B
+ sky130_fd_sc_hd__or4b_4
X_17930_ _18126_/CLK _17930_/D vssd1 vssd1 vccd1 vccd1 _17930_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5580 _13651_/X vssd1 vssd1 vccd1 vccd1 _17670_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10265_ hold2518/X _16579_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10266_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5591 _16965_/Q vssd1 vssd1 vccd1 vccd1 hold5591/X sky130_fd_sc_hd__dlygate4sd3_1
X_12004_ hold4903/X _12308_/B _12003_/X _08167_/A vssd1 vssd1 vccd1 vccd1 _12004_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4890 _11059_/X vssd1 vssd1 vccd1 vccd1 _16843_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17861_ _17861_/CLK _17861_/D vssd1 vssd1 vccd1 vccd1 _17861_/Q sky130_fd_sc_hd__dfxtp_1
X_10196_ hold1041/X hold3644/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10197_/B sky130_fd_sc_hd__mux2_1
X_16812_ _18047_/CLK _16812_/D vssd1 vssd1 vccd1 vccd1 _16812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17792_ _17867_/CLK _17792_/D vssd1 vssd1 vccd1 vccd1 _17792_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout390 _14680_/Y vssd1 vssd1 vccd1 vccd1 _14720_/B sky130_fd_sc_hd__buf_8
XFILLER_0_191_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16743_ _18010_/CLK _16743_/D vssd1 vssd1 vccd1 vccd1 _16743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13955_ hold3025/X _13995_/A2 _13954_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _13955_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_214_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12906_ _12906_/A _12906_/B vssd1 vssd1 vccd1 vccd1 _17478_/D sky130_fd_sc_hd__and2_1
X_16674_ _18200_/CLK _16674_/D vssd1 vssd1 vccd1 vccd1 _16674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13886_ _17749_/Q _13886_/B _13886_/C vssd1 vssd1 vccd1 vccd1 _13886_/X sky130_fd_sc_hd__and3_1
X_18413_ _18413_/CLK _18413_/D vssd1 vssd1 vccd1 vccd1 _18413_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_9_1262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15625_ _17221_/CLK _15625_/D vssd1 vssd1 vccd1 vccd1 _15625_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12837_ _12837_/A _12837_/B vssd1 vssd1 vccd1 vccd1 _17455_/D sky130_fd_sc_hd__and2_1
XFILLER_0_174_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _18376_/CLK _18344_/D vssd1 vssd1 vccd1 vccd1 _18344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15556_ hold1937/X _15560_/A2 _15555_/X _12843_/A vssd1 vssd1 vccd1 vccd1 _15556_/X
+ sky130_fd_sc_hd__o211a_1
X_12768_ _12777_/A _12768_/B vssd1 vssd1 vccd1 vccd1 _17432_/D sky130_fd_sc_hd__and2_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14507_ hold911/X _14553_/B vssd1 vssd1 vccd1 vccd1 _14507_/X sky130_fd_sc_hd__or2_1
XFILLER_0_154_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18275_ _18371_/CLK hold448/X vssd1 vssd1 vccd1 vccd1 _18275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11719_ _12301_/A _11719_/B vssd1 vssd1 vccd1 vccd1 _17063_/D sky130_fd_sc_hd__nor2_1
X_15487_ _17324_/Q _15487_/A2 _15487_/B1 hold737/X _15486_/X vssd1 vssd1 vccd1 vccd1
+ _15489_/C sky130_fd_sc_hd__a221o_1
X_12699_ _12777_/A _12699_/B vssd1 vssd1 vccd1 vccd1 _17409_/D sky130_fd_sc_hd__and2_1
XFILLER_0_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17226_ _18445_/CLK _17226_/D vssd1 vssd1 vccd1 vccd1 _17226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput10 input10/A vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_1
XFILLER_0_154_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14438_ hold2098/X _14433_/B _14437_/X _14372_/A vssd1 vssd1 vccd1 vccd1 _14438_/X
+ sky130_fd_sc_hd__o211a_1
Xinput21 input21/A vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_6
Xinput32 input32/A vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput43 input43/A vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_2
Xinput54 input54/A vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__buf_6
XFILLER_0_163_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17157_ _17157_/CLK _17157_/D vssd1 vssd1 vccd1 vccd1 _17157_/Q sky130_fd_sc_hd__dfxtp_1
Xhold805 hold805/A vssd1 vssd1 vccd1 vccd1 hold805/X sky130_fd_sc_hd__dlygate4sd3_1
X_14369_ _15103_/A hold1587/X _14381_/S vssd1 vssd1 vccd1 vccd1 _14370_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput65 input65/A vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_1
Xhold816 hold816/A vssd1 vssd1 vccd1 vccd1 hold816/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_137_wb_clk_i clkbuf_6_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16147_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16108_ _17331_/CLK _16108_/D vssd1 vssd1 vccd1 vccd1 _16108_/Q sky130_fd_sc_hd__dfxtp_1
Xhold827 hold827/A vssd1 vssd1 vccd1 vccd1 hold827/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold838 hold838/A vssd1 vssd1 vccd1 vccd1 hold838/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 hold849/A vssd1 vssd1 vccd1 vccd1 hold849/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17088_ _17904_/CLK _17088_/D vssd1 vssd1 vccd1 vccd1 _17088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16039_ _18416_/CLK _16039_/D vssd1 vssd1 vccd1 vccd1 hold500/A sky130_fd_sc_hd__dfxtp_1
X_08930_ hold320/X hold807/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08931_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2206 _14007_/X vssd1 vssd1 vccd1 vccd1 _17809_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2217 _18430_/Q vssd1 vssd1 vccd1 vccd1 hold2217/X sky130_fd_sc_hd__dlygate4sd3_1
X_08861_ _15374_/A hold88/X vssd1 vssd1 vccd1 vccd1 _16049_/D sky130_fd_sc_hd__and2_1
Xhold2228 _14807_/X vssd1 vssd1 vccd1 vccd1 _18193_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2239 _14570_/X vssd1 vssd1 vccd1 vccd1 hold2239/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1505 _17770_/Q vssd1 vssd1 vccd1 vccd1 hold1505/X sky130_fd_sc_hd__dlygate4sd3_1
X_07812_ _16286_/Q _07810_/Y hold2253/X _09339_/B vssd1 vssd1 vccd1 vccd1 _07812_/Y
+ sky130_fd_sc_hd__a31oi_1
Xhold1516 _08332_/X vssd1 vssd1 vccd1 vccd1 _15799_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08792_ _15473_/A hold321/X vssd1 vssd1 vccd1 vccd1 _16016_/D sky130_fd_sc_hd__and2_1
Xhold1527 _18297_/Q vssd1 vssd1 vccd1 vccd1 hold1527/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1538 _15764_/Q vssd1 vssd1 vccd1 vccd1 hold1538/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1549 _08422_/X vssd1 vssd1 vccd1 vccd1 _15841_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ _07804_/A hold5989/X _15284_/A _09412_/X vssd1 vssd1 vccd1 vccd1 _09413_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09344_ _15217_/A hold384/A _15182_/A _09352_/D vssd1 vssd1 vccd1 vccd1 _09363_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_168_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09275_ hold992/A _16249_/Q hold271/X vssd1 vssd1 vccd1 vccd1 hold993/A sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08226_ hold1175/X _08209_/B _08225_/X _13801_/C1 vssd1 vssd1 vccd1 vccd1 _08226_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ _08504_/A _15492_/A vssd1 vssd1 vccd1 vccd1 _08170_/S sky130_fd_sc_hd__nand2b_4
XFILLER_0_43_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08088_ _15221_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08088_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_101_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4120 _11524_/X vssd1 vssd1 vccd1 vccd1 _16998_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4131 _16958_/Q vssd1 vssd1 vccd1 vccd1 hold4131/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4142 _17366_/Q vssd1 vssd1 vccd1 vccd1 hold4142/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4153 _09766_/X vssd1 vssd1 vccd1 vccd1 _16412_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4164 _15463_/X vssd1 vssd1 vccd1 vccd1 _15464_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3430 _16347_/Q vssd1 vssd1 vccd1 vccd1 _13246_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4175 hold5958/X vssd1 vssd1 vccd1 vccd1 hold5959/A sky130_fd_sc_hd__buf_4
XTAP_6348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10050_ _13246_/A _09954_/A _10049_/X vssd1 vssd1 vccd1 vccd1 _10050_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3441 hold6116/X vssd1 vssd1 vccd1 vccd1 hold3441/X sky130_fd_sc_hd__buf_1
Xhold4186 _15353_/X vssd1 vssd1 vccd1 vccd1 _15354_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4197 hold5943/X vssd1 vssd1 vccd1 vccd1 hold5944/A sky130_fd_sc_hd__buf_4
XTAP_5614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3452 _11203_/Y vssd1 vssd1 vccd1 vccd1 _16891_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3463 _16541_/Q vssd1 vssd1 vccd1 vccd1 hold3463/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3474 _10638_/Y vssd1 vssd1 vccd1 vccd1 _10639_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2740 _14639_/X vssd1 vssd1 vccd1 vccd1 _18112_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3485 _11176_/Y vssd1 vssd1 vccd1 vccd1 _16882_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2751 _18319_/Q vssd1 vssd1 vccd1 vccd1 hold2751/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3496 _17119_/Q vssd1 vssd1 vccd1 vccd1 hold3496/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2762 _15760_/Q vssd1 vssd1 vccd1 vccd1 hold2762/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2773 _18139_/Q vssd1 vssd1 vccd1 vccd1 hold2773/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2784 _08075_/X vssd1 vssd1 vccd1 vccd1 _15677_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2795 _14255_/X vssd1 vssd1 vccd1 vccd1 _17928_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13740_ _13773_/A _13740_/B vssd1 vssd1 vccd1 vccd1 _13740_/X sky130_fd_sc_hd__or2_1
X_10952_ hold1933/X hold3724/X _11144_/C vssd1 vssd1 vccd1 vccd1 _10953_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_230_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13671_ _13794_/A _13671_/B vssd1 vssd1 vccd1 vccd1 _13671_/X sky130_fd_sc_hd__or2_1
XFILLER_0_210_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10883_ _17988_/Q _16785_/Q _11654_/S vssd1 vssd1 vccd1 vccd1 _10884_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15410_ hold829/X _15448_/A2 _15446_/B1 hold426/X vssd1 vssd1 vccd1 vccd1 _15410_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12622_ hold2881/X hold2277/X _12850_/S vssd1 vssd1 vccd1 vccd1 _12622_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16390_ _18411_/CLK _16390_/D vssd1 vssd1 vccd1 vccd1 _16390_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15341_ _16298_/Q _09362_/A _09392_/B hold716/X _15340_/X vssd1 vssd1 vccd1 vccd1
+ _15342_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_171_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12553_ hold2834/X hold3599/X _12925_/S vssd1 vssd1 vccd1 vccd1 _12553_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_164_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11504_ hold1511/X _16992_/Q _12335_/C vssd1 vssd1 vccd1 vccd1 _11505_/B sky130_fd_sc_hd__mux2_1
X_18060_ _18060_/CLK _18060_/D vssd1 vssd1 vccd1 vccd1 _18060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15272_ _15480_/A _15272_/B _15272_/C _15272_/D vssd1 vssd1 vccd1 vccd1 _15272_/X
+ sky130_fd_sc_hd__or4_1
X_12484_ _17335_/Q _12506_/B vssd1 vssd1 vccd1 vccd1 _12484_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17011_ _17859_/CLK _17011_/D vssd1 vssd1 vccd1 vccd1 _17011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14223_ hold2149/X _14216_/Y _14222_/X _13895_/A vssd1 vssd1 vccd1 vccd1 _14223_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11435_ hold2964/X hold5359/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11436_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_105_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_230_wb_clk_i clkbuf_6_63_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18149_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11366_ hold1440/X hold5103/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11367_/B sky130_fd_sc_hd__mux2_1
X_14154_ _15553_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14154_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13105_ _13105_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13105_/X sky130_fd_sc_hd__and2_1
X_10317_ _10551_/A _10317_/B vssd1 vssd1 vccd1 vccd1 _10317_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11297_ _17771_/Q hold4364/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11298_/B sky130_fd_sc_hd__mux2_1
X_14085_ hold2189/X _14094_/B _14084_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _14085_/X
+ sky130_fd_sc_hd__o211a_1
X_13036_ hold907/X _13035_/X hold904/A vssd1 vssd1 vccd1 vccd1 hold908/A sky130_fd_sc_hd__mux2_1
X_10248_ _10536_/A _10248_/B vssd1 vssd1 vccd1 vccd1 _10248_/X sky130_fd_sc_hd__or2_1
XFILLER_0_219_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17913_ _17913_/CLK _17913_/D vssd1 vssd1 vccd1 vccd1 _17913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17844_ _17856_/CLK _17844_/D vssd1 vssd1 vccd1 vccd1 _17844_/Q sky130_fd_sc_hd__dfxtp_1
X_10179_ _10563_/A _10179_/B vssd1 vssd1 vccd1 vccd1 _10179_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17775_ _17799_/CLK _17775_/D vssd1 vssd1 vccd1 vccd1 _17775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14987_ hold3072/X hold447/X _14986_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _14987_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_178_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16726_ _17929_/CLK _16726_/D vssd1 vssd1 vccd1 vccd1 _16726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13938_ _14726_/A hold2821/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13939_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_191_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16657_ _18215_/CLK _16657_/D vssd1 vssd1 vccd1 vccd1 _16657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13869_ hold3493/X _13581_/A _13868_/X vssd1 vssd1 vccd1 vccd1 _13869_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_201_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_233_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15608_ _17724_/CLK _15608_/D vssd1 vssd1 vccd1 vccd1 _15608_/Q sky130_fd_sc_hd__dfxtp_1
X_16588_ _18129_/CLK _16588_/D vssd1 vssd1 vccd1 vccd1 _16588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18327_ _18327_/CLK _18327_/D vssd1 vssd1 vccd1 vccd1 _18327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_389_wb_clk_i clkbuf_6_38_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17897_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15539_ _15539_/A _15549_/B vssd1 vssd1 vccd1 vccd1 _15539_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09060_ hold320/X hold459/X _09060_/S vssd1 vssd1 vccd1 vccd1 _09061_/B sky130_fd_sc_hd__mux2_1
X_18258_ _18356_/CLK hold646/X vssd1 vssd1 vccd1 vccd1 hold645/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_318_wb_clk_i clkbuf_6_47_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17895_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_142_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08011_ _15525_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08011_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17209_ _17209_/CLK _17209_/D vssd1 vssd1 vccd1 vccd1 _17209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18189_ _18221_/CLK _18189_/D vssd1 vssd1 vccd1 vccd1 _18189_/Q sky130_fd_sc_hd__dfxtp_1
Xhold602 hold602/A vssd1 vssd1 vccd1 vccd1 hold602/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold613 hold613/A vssd1 vssd1 vccd1 vccd1 hold613/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold624 hold624/A vssd1 vssd1 vccd1 vccd1 hold624/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 hold635/A vssd1 vssd1 vccd1 vccd1 hold635/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold646 hold646/A vssd1 vssd1 vccd1 vccd1 hold646/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold657 hold657/A vssd1 vssd1 vccd1 vccd1 hold657/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold668 hold668/A vssd1 vssd1 vccd1 vccd1 hold668/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold679 hold679/A vssd1 vssd1 vccd1 vccd1 hold679/X sky130_fd_sc_hd__buf_4
X_09962_ hold1177/X hold3822/X _10634_/C vssd1 vssd1 vccd1 vccd1 _09963_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_12_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08913_ _12394_/A _08913_/B vssd1 vssd1 vccd1 vccd1 _16074_/D sky130_fd_sc_hd__and2_1
Xhold2003 _09095_/X vssd1 vssd1 vccd1 vccd1 _16162_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09893_ hold1607/X _16455_/Q _10004_/C vssd1 vssd1 vccd1 vccd1 _09894_/B sky130_fd_sc_hd__mux2_1
Xhold2014 _14400_/X vssd1 vssd1 vccd1 vccd1 _17998_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2025 _18212_/Q vssd1 vssd1 vccd1 vccd1 hold2025/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2036 _14705_/X vssd1 vssd1 vccd1 vccd1 _18144_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2047 _18120_/Q vssd1 vssd1 vccd1 vccd1 hold2047/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1302 _09071_/X vssd1 vssd1 vccd1 vccd1 _16150_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08844_ hold5/X hold153/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08845_/B sky130_fd_sc_hd__mux2_1
Xhold1313 _18210_/Q vssd1 vssd1 vccd1 vccd1 hold1313/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2058 _18200_/Q vssd1 vssd1 vccd1 vccd1 hold2058/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2069 _07967_/X vssd1 vssd1 vccd1 vccd1 _15626_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1324 _07909_/X vssd1 vssd1 vccd1 vccd1 _15598_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1335 _09175_/X vssd1 vssd1 vccd1 vccd1 _16200_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1346 _15644_/Q vssd1 vssd1 vccd1 vccd1 hold1346/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1357 _07878_/X vssd1 vssd1 vccd1 vccd1 _15584_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_240_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08775_ hold53/X hold477/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08776_/B sky130_fd_sc_hd__mux2_1
Xhold1368 hold1368/A vssd1 vssd1 vccd1 vccd1 hold911/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_224_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1379 _08473_/X vssd1 vssd1 vccd1 vccd1 _15865_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_34_wb_clk_i clkbuf_6_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17850_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_135_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09327_ _15549_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09327_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09258_ _12753_/A _09258_/B vssd1 vssd1 vccd1 vccd1 _16240_/D sky130_fd_sc_hd__and2_1
XFILLER_0_211_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08209_ _15163_/A _08209_/B vssd1 vssd1 vccd1 vccd1 _08209_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09189_ hold2289/X _09218_/B _09188_/X _12786_/A vssd1 vssd1 vccd1 vccd1 _09189_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11220_ hold3476/X _11124_/A _11219_/X vssd1 vssd1 vccd1 vccd1 _11220_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_160_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11151_ hold4469/X _11043_/A _11150_/X vssd1 vssd1 vccd1 vccd1 _11151_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10102_ hold3644/X _10625_/B _10101_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _10102_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11082_ _11109_/A _11082_/B vssd1 vssd1 vccd1 vccd1 _11082_/X sky130_fd_sc_hd__or2_1
XTAP_6145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3260 _10279_/X vssd1 vssd1 vccd1 vccd1 _16583_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10033_ _11203_/A _10033_/B vssd1 vssd1 vccd1 vccd1 _10033_/Y sky130_fd_sc_hd__nor2_1
Xhold3271 _09589_/X vssd1 vssd1 vccd1 vccd1 _16353_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14910_ _14980_/A _14910_/B vssd1 vssd1 vccd1 vccd1 _14910_/X sky130_fd_sc_hd__or2_1
Xhold3282 _16651_/Q vssd1 vssd1 vccd1 vccd1 hold3282/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15890_ _17523_/CLK _15890_/D vssd1 vssd1 vccd1 vccd1 _15890_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3293 _10189_/X vssd1 vssd1 vccd1 vccd1 _16553_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2570 _15168_/X vssd1 vssd1 vccd1 vccd1 _18367_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ hold1313/X _14828_/B _14840_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14841_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2581 _09113_/X vssd1 vssd1 vccd1 vccd1 _16171_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2592 _08416_/X vssd1 vssd1 vccd1 vccd1 _15838_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1880 _09437_/X vssd1 vssd1 vccd1 vccd1 _16304_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ _17720_/CLK _17560_/D vssd1 vssd1 vccd1 vccd1 _17560_/Q sky130_fd_sc_hd__dfxtp_1
X_14772_ _15165_/A _14772_/B vssd1 vssd1 vccd1 vccd1 _14772_/Y sky130_fd_sc_hd__nand2_1
Xhold1891 _18285_/Q vssd1 vssd1 vccd1 vccd1 hold1891/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11984_ hold1837/X _17152_/Q _12371_/C vssd1 vssd1 vccd1 vccd1 _11985_/B sky130_fd_sc_hd__mux2_1
X_16511_ _18081_/CLK _16511_/D vssd1 vssd1 vccd1 vccd1 _16511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13723_ _13817_/A _13817_/B _13722_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _13723_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17491_ _17491_/CLK _17491_/D vssd1 vssd1 vccd1 vccd1 _17491_/Q sky130_fd_sc_hd__dfxtp_1
X_10935_ _11694_/A _10935_/B vssd1 vssd1 vccd1 vccd1 _10935_/X sky130_fd_sc_hd__or2_1
XFILLER_0_230_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16442_ _18323_/CLK _16442_/D vssd1 vssd1 vccd1 vccd1 _16442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ hold5490/X _13883_/B _13653_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13654_/X
+ sky130_fd_sc_hd__o211a_1
X_10866_ _11136_/A _10866_/B vssd1 vssd1 vccd1 vccd1 _10866_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ hold3265/X _12604_/X _12923_/S vssd1 vssd1 vccd1 vccd1 _12606_/B sky130_fd_sc_hd__mux2_1
X_16373_ _18324_/CLK _16373_/D vssd1 vssd1 vccd1 vccd1 _16373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ hold5285/X _13871_/B _13584_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13585_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10797_ _11091_/A _10797_/B vssd1 vssd1 vccd1 vccd1 _10797_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18112_ _18234_/CLK _18112_/D vssd1 vssd1 vccd1 vccd1 _18112_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15324_ _15324_/A _15324_/B vssd1 vssd1 vccd1 vccd1 _18408_/D sky130_fd_sc_hd__and2_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12536_ hold4523/X _12535_/X _12929_/S vssd1 vssd1 vccd1 vccd1 _12536_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_411_wb_clk_i clkbuf_6_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17899_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18043_ _18043_/CLK _18043_/D vssd1 vssd1 vccd1 vccd1 _18043_/Q sky130_fd_sc_hd__dfxtp_1
X_15255_ hold779/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15255_/X sky130_fd_sc_hd__or2_1
X_12467_ hold23/X _12445_/A _08868_/X _12466_/X _09003_/A vssd1 vssd1 vccd1 vccd1
+ hold24/A sky130_fd_sc_hd__o311a_1
X_14206_ _14330_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14206_/X sky130_fd_sc_hd__or2_1
X_11418_ _11697_/A _11418_/B vssd1 vssd1 vccd1 vccd1 _11418_/X sky130_fd_sc_hd__or2_1
XFILLER_0_201_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15186_ hold2213/X _15221_/B _15185_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _15186_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12398_ _12416_/A _12398_/B vssd1 vssd1 vccd1 vccd1 _17292_/D sky130_fd_sc_hd__and2_1
XFILLER_0_239_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14137_ hold2167/X _14142_/B _14136_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _14137_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_201_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11349_ _11637_/A _11349_/B vssd1 vssd1 vccd1 vccd1 _11349_/X sky130_fd_sc_hd__or2_1
XFILLER_0_240_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14068_ _14461_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14068_/X sky130_fd_sc_hd__or2_1
XFILLER_0_219_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13019_ _13019_/A hold899/X hold892/X hold920/X vssd1 vssd1 vccd1 vccd1 hold900/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_183_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17827_ _18065_/CLK _17827_/D vssd1 vssd1 vccd1 vccd1 _17827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08560_ hold172/X hold610/X _08592_/S vssd1 vssd1 vccd1 vccd1 _08561_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17758_ _17886_/CLK _17758_/D vssd1 vssd1 vccd1 vccd1 _17758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_234_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16709_ _18072_/CLK _16709_/D vssd1 vssd1 vccd1 vccd1 _16709_/Q sky130_fd_sc_hd__dfxtp_1
X_08491_ hold1340/X _08486_/B _08490_/X _08347_/A vssd1 vssd1 vccd1 vccd1 _08491_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17689_ _17689_/CLK _17689_/D vssd1 vssd1 vccd1 vccd1 _17689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09112_ _15553_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09112_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_152_wb_clk_i clkbuf_6_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18240_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_165_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09043_ _12440_/A _09043_/B vssd1 vssd1 vccd1 vccd1 _16138_/D sky130_fd_sc_hd__and2_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold410 hold410/A vssd1 vssd1 vccd1 vccd1 hold410/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold421 hold421/A vssd1 vssd1 vccd1 vccd1 input64/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 hold432/A vssd1 vssd1 vccd1 vccd1 hold432/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 input55/X vssd1 vssd1 vccd1 vccd1 hold443/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 hold454/A vssd1 vssd1 vccd1 vccd1 hold454/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold465 hold465/A vssd1 vssd1 vccd1 vccd1 hold465/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold476 hold476/A vssd1 vssd1 vccd1 vccd1 hold476/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 hold487/A vssd1 vssd1 vccd1 vccd1 hold487/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold498 hold498/A vssd1 vssd1 vccd1 vccd1 hold498/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 hold1367/X vssd1 vssd1 vccd1 vccd1 _14972_/A sky130_fd_sc_hd__buf_8
X_09945_ _11109_/A _09945_/B vssd1 vssd1 vccd1 vccd1 _09945_/X sky130_fd_sc_hd__or2_1
Xfanout912 hold820/X vssd1 vssd1 vccd1 vccd1 _14960_/A sky130_fd_sc_hd__buf_8
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout923 hold1022/X vssd1 vssd1 vccd1 vccd1 _14166_/A sky130_fd_sc_hd__buf_6
Xfanout934 hold1183/X vssd1 vssd1 vccd1 vccd1 _14529_/A sky130_fd_sc_hd__clkbuf_16
Xfanout945 hold1193/X vssd1 vssd1 vccd1 vccd1 _14164_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_216_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09876_ _10560_/A _09876_/B vssd1 vssd1 vccd1 vccd1 _09876_/X sky130_fd_sc_hd__or2_1
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 _18329_/Q vssd1 vssd1 vccd1 vccd1 hold1110/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 _16259_/Q vssd1 vssd1 vccd1 vccd1 hold1121/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1132 _16287_/Q vssd1 vssd1 vccd1 vccd1 _07786_/A sky130_fd_sc_hd__buf_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _12390_/A hold462/X vssd1 vssd1 vccd1 vccd1 _16032_/D sky130_fd_sc_hd__and2_1
XFILLER_0_99_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1143 _15853_/Q vssd1 vssd1 vccd1 vccd1 hold1143/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1154 _13914_/X vssd1 vssd1 vccd1 vccd1 _13915_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1165 _18392_/Q vssd1 vssd1 vccd1 vccd1 hold1165/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1176 _08226_/X vssd1 vssd1 vccd1 vccd1 _15749_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1187 _09141_/X vssd1 vssd1 vccd1 vccd1 _16183_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _15344_/A hold413/X vssd1 vssd1 vccd1 vccd1 _15999_/D sky130_fd_sc_hd__and2_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 _15815_/Q vssd1 vssd1 vccd1 vccd1 hold1198/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ hold77/X hold689/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08690_/B sky130_fd_sc_hd__mux2_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10720_ hold4056/X _11222_/B _10719_/X _14526_/C1 vssd1 vssd1 vccd1 vccd1 _10720_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10651_ _10651_/A _10651_/B vssd1 vssd1 vccd1 vccd1 _16707_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_82_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10582_ _10651_/A _10582_/B vssd1 vssd1 vccd1 vccd1 _10582_/Y sky130_fd_sc_hd__nor2_1
X_13370_ hold1380/X hold4495/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13371_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12321_ hold4298/X _13314_/A _12320_/X vssd1 vssd1 vccd1 vccd1 _12321_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15040_ _15394_/A _15040_/B vssd1 vssd1 vccd1 vccd1 _18305_/D sky130_fd_sc_hd__and2_1
XFILLER_0_107_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12252_ _12267_/A _12252_/B vssd1 vssd1 vccd1 vccd1 _12252_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11203_ _11203_/A _11203_/B vssd1 vssd1 vccd1 vccd1 _11203_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_121_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12183_ _13749_/A _12183_/B vssd1 vssd1 vccd1 vccd1 _12183_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11134_ hold5297/X _11732_/B _11133_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _11134_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16991_ _17871_/CLK _16991_/D vssd1 vssd1 vccd1 vccd1 _16991_/Q sky130_fd_sc_hd__dfxtp_1
X_15942_ _17335_/CLK _15942_/D vssd1 vssd1 vccd1 vccd1 hold165/A sky130_fd_sc_hd__dfxtp_1
X_11065_ hold4729/X _11162_/B _11064_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _11065_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3090 _15526_/X vssd1 vssd1 vccd1 vccd1 _18441_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10016_ _16496_/Q _10022_/B _10022_/C vssd1 vssd1 vccd1 vccd1 _10016_/X sky130_fd_sc_hd__and3_1
XFILLER_0_200_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ _17584_/CLK _15873_/D vssd1 vssd1 vccd1 vccd1 _15873_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14824_ _15163_/A _14828_/B vssd1 vssd1 vccd1 vccd1 _14824_/Y sky130_fd_sc_hd__nand2_1
X_17612_ _17734_/CLK _17612_/D vssd1 vssd1 vccd1 vccd1 _17612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17543_ _18392_/CLK _17543_/D vssd1 vssd1 vccd1 vccd1 _17543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ hold2836/X _14774_/B _14754_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _14755_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ _12255_/A _11967_/B vssd1 vssd1 vccd1 vccd1 _11967_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_230_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13706_ hold1370/X _17689_/Q _13817_/C vssd1 vssd1 vccd1 vccd1 _13707_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_86_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10918_ hold4955/X _11204_/B _10917_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _10918_/X
+ sky130_fd_sc_hd__o211a_1
X_17474_ _17881_/CLK _17474_/D vssd1 vssd1 vccd1 vccd1 _17474_/Q sky130_fd_sc_hd__dfxtp_1
X_14686_ hold911/X _14732_/B vssd1 vssd1 vccd1 vccd1 _14686_/X sky130_fd_sc_hd__or2_1
X_11898_ _13407_/A _11898_/B vssd1 vssd1 vccd1 vccd1 _11898_/X sky130_fd_sc_hd__or2_1
X_16425_ _18370_/CLK _16425_/D vssd1 vssd1 vccd1 vccd1 _16425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13637_ hold1515/X hold4541/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13638_/B sky130_fd_sc_hd__mux2_1
X_10849_ hold5187/X _11153_/B _10848_/X _14354_/A vssd1 vssd1 vccd1 vccd1 _10849_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16356_ _18369_/CLK _16356_/D vssd1 vssd1 vccd1 vccd1 _16356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13568_ hold1770/X _17643_/Q _13841_/C vssd1 vssd1 vccd1 vccd1 _13569_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_171_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15307_ hold759/X _09357_/A _09386_/D hold866/X _15306_/X vssd1 vssd1 vccd1 vccd1
+ _15312_/B sky130_fd_sc_hd__a221o_1
X_12519_ _12987_/A _12519_/B vssd1 vssd1 vccd1 vccd1 _17349_/D sky130_fd_sc_hd__and2_1
X_16287_ _18460_/CLK _16287_/D vssd1 vssd1 vccd1 vccd1 _16287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13499_ hold2718/X hold5507/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13500_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_180_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5409 _11662_/X vssd1 vssd1 vccd1 vccd1 _17044_/D sky130_fd_sc_hd__dlygate4sd3_1
X_18026_ _18056_/CLK _18026_/D vssd1 vssd1 vccd1 vccd1 _18026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15238_ hold525/X _15484_/A2 _09392_/D hold726/X vssd1 vssd1 vccd1 vccd1 _15238_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_160_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4708 _09949_/X vssd1 vssd1 vccd1 vccd1 _16473_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4719 _11773_/Y vssd1 vssd1 vccd1 vccd1 _17081_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15169_ _15169_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15169_/X sky130_fd_sc_hd__or2_1
XFILLER_0_238_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout208 _11792_/B vssd1 vssd1 vccd1 vccd1 _11222_/B sky130_fd_sc_hd__buf_4
Xfanout219 _10013_/B vssd1 vssd1 vccd1 vccd1 _10004_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07991_ hold1103/X _07991_/A2 _07990_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _07991_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_197_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09730_ hold4891/X _11171_/B _09729_/X _14372_/A vssd1 vssd1 vccd1 vccd1 _09730_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09661_ hold4687/X _10031_/B _09660_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09661_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08612_ _09061_/A _08612_/B vssd1 vssd1 vccd1 vccd1 _15928_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09592_ hold3662/X _10070_/B _09591_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _09592_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08543_ _09003_/A _08543_/B vssd1 vssd1 vccd1 vccd1 _15895_/D sky130_fd_sc_hd__and2_1
XFILLER_0_89_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_222_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_333_wb_clk_i clkbuf_6_41_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17279_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08474_ _15207_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08474_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5910 hold5910/A vssd1 vssd1 vccd1 vccd1 load_status[1] sky130_fd_sc_hd__buf_12
X_09026_ hold169/X hold344/X _09060_/S vssd1 vssd1 vccd1 vccd1 hold345/A sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5921 _17520_/Q vssd1 vssd1 vccd1 vccd1 hold935/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5932 _18414_/Q vssd1 vssd1 vccd1 vccd1 hold5932/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5943 _18412_/Q vssd1 vssd1 vccd1 vccd1 hold5943/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5954 _18421_/Q vssd1 vssd1 vccd1 vccd1 hold5954/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold240 hold240/A vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5965 hold5965/A vssd1 vssd1 vccd1 vccd1 hold5965/X sky130_fd_sc_hd__clkbuf_4
Xhold251 hold251/A vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5976 _17521_/Q vssd1 vssd1 vccd1 vccd1 hold5976/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold262 hold262/A vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5987 hold6123/X vssd1 vssd1 vccd1 vccd1 _09456_/C sky130_fd_sc_hd__buf_1
Xhold273 hold273/A vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5998 _16920_/Q vssd1 vssd1 vccd1 vccd1 hold5998/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 hold284/A vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 hold295/A vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__buf_2
Xfanout720 _15176_/C1 vssd1 vssd1 vccd1 vccd1 _15044_/A sky130_fd_sc_hd__buf_4
XFILLER_0_102_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout731 _09003_/A vssd1 vssd1 vccd1 vccd1 _09061_/A sky130_fd_sc_hd__buf_2
X_09928_ hold5807/X _10022_/B _09927_/X _15202_/C1 vssd1 vssd1 vccd1 vccd1 _09928_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout742 _13675_/C1 vssd1 vssd1 vccd1 vccd1 _08379_/A sky130_fd_sc_hd__buf_4
Xfanout753 _13929_/A vssd1 vssd1 vccd1 vccd1 _13927_/A sky130_fd_sc_hd__buf_4
Xfanout764 fanout843/X vssd1 vssd1 vccd1 vccd1 _14131_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_176_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout775 _08149_/A vssd1 vssd1 vccd1 vccd1 _08145_/A sky130_fd_sc_hd__buf_4
Xfanout786 fanout791/X vssd1 vssd1 vccd1 vccd1 _14143_/C1 sky130_fd_sc_hd__buf_4
X_09859_ hold3582/X _10049_/B _09858_/X _15146_/C1 vssd1 vssd1 vccd1 vccd1 _09859_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout797 fanout816/X vssd1 vssd1 vccd1 vccd1 _15054_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_232_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12870_ _12888_/A _12870_/B vssd1 vssd1 vccd1 vccd1 _17466_/D sky130_fd_sc_hd__and2_1
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 fanout299/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_113 _14988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11821_ hold5697/X _12299_/B _11820_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _11821_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 hold1367/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14540_ hold2443/X _14541_/B _14539_/Y _14344_/A vssd1 vssd1 vccd1 vccd1 _14540_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _12331_/A _11752_/B vssd1 vssd1 vccd1 vccd1 _11752_/Y sky130_fd_sc_hd__nor2_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ hold2794/X hold3490/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10704_/B sky130_fd_sc_hd__mux2_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14471_ _14596_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14471_/X sky130_fd_sc_hd__or2_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ hold5054/X _12317_/B _11682_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _11683_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16210_ _17445_/CLK _16210_/D vssd1 vssd1 vccd1 vccd1 _16210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13422_ _13722_/A _13422_/B vssd1 vssd1 vccd1 vccd1 _13422_/X sky130_fd_sc_hd__or2_1
X_10634_ _10634_/A _10634_/B _10634_/C vssd1 vssd1 vccd1 vccd1 _10634_/X sky130_fd_sc_hd__and3_1
X_17190_ _17190_/CLK _17190_/D vssd1 vssd1 vccd1 vccd1 _17190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16141_ _17336_/CLK _16141_/D vssd1 vssd1 vccd1 vccd1 _16141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13353_ _13794_/A _13353_/B vssd1 vssd1 vccd1 vccd1 _13353_/X sky130_fd_sc_hd__or2_1
X_10565_ _10565_/A _10568_/B _10571_/C vssd1 vssd1 vccd1 vccd1 _10565_/X sky130_fd_sc_hd__and3_1
XFILLER_0_183_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12304_ _13819_/A _12304_/B vssd1 vssd1 vccd1 vccd1 _12304_/Y sky130_fd_sc_hd__nor2_1
X_16072_ _17303_/CLK _16072_/D vssd1 vssd1 vccd1 vccd1 hold532/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13284_ hold4356/X _13283_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13284_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10496_ hold2727/X hold3257/X _10634_/C vssd1 vssd1 vccd1 vccd1 _10497_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15023_ _15185_/A hold1527/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15024_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12235_ hold5683/X _12329_/B _12234_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _12235_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12166_ hold5036/X _12356_/B _12165_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _12166_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11117_ hold2443/X hold3956/X _11216_/C vssd1 vssd1 vccd1 vccd1 _11118_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_236_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12097_ hold5090/X _12353_/B _12096_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _12097_/X
+ sky130_fd_sc_hd__o211a_1
X_16974_ _17886_/CLK _16974_/D vssd1 vssd1 vccd1 vccd1 _16974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15925_ _17300_/CLK _15925_/D vssd1 vssd1 vccd1 vccd1 hold886/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11048_ hold1956/X hold3771/X _11144_/C vssd1 vssd1 vccd1 vccd1 _11049_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_189_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 input8/A vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_1
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15856_ _15856_/CLK _15856_/D vssd1 vssd1 vccd1 vccd1 _15856_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14807_ hold6053/X _14828_/B _14806_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _14807_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_232_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15787_ _17686_/CLK _15787_/D vssd1 vssd1 vccd1 vccd1 _15787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12999_ _15244_/A _12999_/B vssd1 vssd1 vccd1 vccd1 _17509_/D sky130_fd_sc_hd__and2_1
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17526_ _17535_/CLK _17526_/D vssd1 vssd1 vccd1 vccd1 _17526_/Q sky130_fd_sc_hd__dfxtp_1
X_14738_ _15185_/A _14780_/B vssd1 vssd1 vccd1 vccd1 _14738_/X sky130_fd_sc_hd__or2_1
XFILLER_0_146_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17457_ _18458_/CLK _17457_/D vssd1 vssd1 vccd1 vccd1 _17457_/Q sky130_fd_sc_hd__dfxtp_1
X_14669_ hold1732/X _14664_/B _14668_/X _14853_/C1 vssd1 vssd1 vccd1 vccd1 _14669_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16408_ _18321_/CLK _16408_/D vssd1 vssd1 vccd1 vccd1 _16408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08190_ hold1099/X _08213_/B _08189_/X _13765_/C1 vssd1 vssd1 vccd1 vccd1 _08190_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17388_ _18455_/CLK _17388_/D vssd1 vssd1 vccd1 vccd1 _17388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16339_ _18342_/CLK _16339_/D vssd1 vssd1 vccd1 vccd1 _16339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5206 _10975_/X vssd1 vssd1 vccd1 vccd1 _16815_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5217 _17249_/Q vssd1 vssd1 vccd1 vccd1 hold5217/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5228 _10738_/X vssd1 vssd1 vccd1 vccd1 _16736_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5239 _17045_/Q vssd1 vssd1 vccd1 vccd1 hold5239/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4505 _10222_/X vssd1 vssd1 vccd1 vccd1 _16564_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18009_ _18041_/CLK _18009_/D vssd1 vssd1 vccd1 vccd1 _18009_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4516 _13882_/Y vssd1 vssd1 vccd1 vccd1 _17747_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4527 _16692_/Q vssd1 vssd1 vccd1 vccd1 hold4527/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4538 _10156_/X vssd1 vssd1 vccd1 vccd1 _16542_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3804 _10255_/X vssd1 vssd1 vccd1 vccd1 _16575_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4549 _16916_/Q vssd1 vssd1 vccd1 vccd1 hold4549/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3815 _10249_/X vssd1 vssd1 vccd1 vccd1 _16573_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3826 _17414_/Q vssd1 vssd1 vccd1 vccd1 hold3826/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3837 _10951_/X vssd1 vssd1 vccd1 vccd1 _16807_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3848 _16678_/Q vssd1 vssd1 vccd1 vccd1 hold3848/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3859 _11029_/X vssd1 vssd1 vccd1 vccd1 _16833_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07974_ _15543_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _07974_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09713_ hold2579/X hold3586/X _10025_/C vssd1 vssd1 vccd1 vccd1 _09714_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_214_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09644_ hold1891/X hold4512/X _10028_/C vssd1 vssd1 vccd1 vccd1 _09645_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_214_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09575_ hold2457/X _13262_/A _10601_/C vssd1 vssd1 vccd1 vccd1 _09576_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_210_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ hold618/X hold813/X _08528_/S vssd1 vssd1 vccd1 vccd1 hold814/A sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_212_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08457_ hold2826/X _08488_/B _08456_/X _13729_/C1 vssd1 vssd1 vccd1 vccd1 _08457_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_212_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08388_ _14443_/A hold1084/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08389_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10350_ _10536_/A _10350_/B vssd1 vssd1 vccd1 vccd1 _10350_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09009_ _09057_/A _09009_/B vssd1 vssd1 vccd1 vccd1 _16121_/D sky130_fd_sc_hd__and2_1
XFILLER_0_143_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5740 _13390_/X vssd1 vssd1 vccd1 vccd1 _17583_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10281_ _10476_/A _10281_/B vssd1 vssd1 vccd1 vccd1 _10281_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5751 _17245_/Q vssd1 vssd1 vccd1 vccd1 hold5751/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5762 _12268_/X vssd1 vssd1 vccd1 vccd1 _17246_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5773 _17150_/Q vssd1 vssd1 vccd1 vccd1 hold5773/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5784 _13711_/X vssd1 vssd1 vccd1 vccd1 _17690_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12020_ hold1953/X hold3935/X _13796_/S vssd1 vssd1 vccd1 vccd1 _12021_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_218_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5795 _17233_/Q vssd1 vssd1 vccd1 vccd1 hold5795/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_217_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout550 _08335_/B vssd1 vssd1 vccd1 vccd1 _08333_/B sky130_fd_sc_hd__buf_8
Xfanout561 _08100_/B vssd1 vssd1 vccd1 vccd1 _08094_/B sky130_fd_sc_hd__buf_6
XFILLER_0_233_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout572 _07884_/Y vssd1 vssd1 vccd1 vccd1 _07918_/B sky130_fd_sc_hd__buf_6
Xfanout583 _13055_/X vssd1 vssd1 vccd1 vccd1 _13244_/S sky130_fd_sc_hd__buf_8
X_13971_ hold1239/X _13995_/A2 _13970_/X _14211_/C1 vssd1 vssd1 vccd1 vccd1 _13971_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout594 _12871_/S vssd1 vssd1 vccd1 vccd1 _12844_/S sky130_fd_sc_hd__buf_6
X_15710_ _17278_/CLK hold110/X vssd1 vssd1 vccd1 vccd1 _15710_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_255_wb_clk_i clkbuf_6_58_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18024_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12922_ hold1319/X _17485_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12922_/X sky130_fd_sc_hd__mux2_1
X_16690_ _18170_/CLK _16690_/D vssd1 vssd1 vccd1 vccd1 _16690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15641_ _17187_/CLK _15641_/D vssd1 vssd1 vccd1 vccd1 _15641_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12853_ hold2924/X hold3318/X _12916_/S vssd1 vssd1 vccd1 vccd1 _12853_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_200_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18360_ _18384_/CLK _18360_/D vssd1 vssd1 vccd1 vccd1 _18360_/Q sky130_fd_sc_hd__dfxtp_1
X_11804_ hold1883/X _17092_/Q _12227_/S vssd1 vssd1 vccd1 vccd1 _11805_/B sky130_fd_sc_hd__mux2_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _17242_/CLK _15572_/D vssd1 vssd1 vccd1 vccd1 _15572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12784_ hold982/X hold3396/X _12838_/S vssd1 vssd1 vccd1 vccd1 _12784_/X sky130_fd_sc_hd__mux2_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _18413_/CLK _17311_/D vssd1 vssd1 vccd1 vccd1 hold118/A sky130_fd_sc_hd__dfxtp_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14988_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14523_/X sky130_fd_sc_hd__or2_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18291_ _18361_/CLK _18291_/D vssd1 vssd1 vccd1 vccd1 _18291_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11735_ _17069_/Q _11744_/B _11738_/C vssd1 vssd1 vccd1 vccd1 _11735_/X sky130_fd_sc_hd__and3_1
XFILLER_0_113_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17242_/CLK _17242_/D vssd1 vssd1 vccd1 vccd1 _17242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14454_ hold1688/X _14487_/B _14453_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _14454_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11666_ hold3006/X _17046_/Q _11783_/C vssd1 vssd1 vccd1 vccd1 _11667_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13405_ hold5507/X _13883_/B _13404_/X _08347_/A vssd1 vssd1 vccd1 vccd1 _13405_/X
+ sky130_fd_sc_hd__o211a_1
X_10617_ hold3515/X _11103_/A _10616_/X vssd1 vssd1 vccd1 vccd1 _10617_/Y sky130_fd_sc_hd__a21oi_1
X_17173_ _17779_/CLK _17173_/D vssd1 vssd1 vccd1 vccd1 _17173_/Q sky130_fd_sc_hd__dfxtp_1
X_14385_ _14726_/A hold2511/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14386_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11597_ hold1558/X hold5309/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11598_/B sky130_fd_sc_hd__mux2_1
X_16124_ _16124_/CLK _16124_/D vssd1 vssd1 vccd1 vccd1 hold755/A sky130_fd_sc_hd__dfxtp_1
X_13336_ hold4075/X _13808_/B _13335_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _13336_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10548_ _10551_/A _10548_/B vssd1 vssd1 vccd1 vccd1 _10548_/X sky130_fd_sc_hd__or2_1
XFILLER_0_45_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16055_ _17309_/CLK _16055_/D vssd1 vssd1 vccd1 vccd1 hold187/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13267_ _13266_/X _16926_/Q _13267_/S vssd1 vssd1 vccd1 vccd1 _13267_/X sky130_fd_sc_hd__mux2_1
X_10479_ _11091_/A _10479_/B vssd1 vssd1 vccd1 vccd1 _10479_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15006_ _15221_/A hold447/X vssd1 vssd1 vccd1 vccd1 _15006_/Y sky130_fd_sc_hd__nand2_1
X_12218_ hold1775/X hold5456/X _12323_/C vssd1 vssd1 vccd1 vccd1 _12219_/B sky130_fd_sc_hd__mux2_1
X_13198_ _13198_/A _13294_/B vssd1 vssd1 vccd1 vccd1 _13198_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12149_ hold2431/X hold4030/X _12371_/C vssd1 vssd1 vccd1 vccd1 _12150_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1709 _09229_/X vssd1 vssd1 vccd1 vccd1 _16226_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_236_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16957_ _17891_/CLK _16957_/D vssd1 vssd1 vccd1 vccd1 _16957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15908_ _16120_/CLK _15908_/D vssd1 vssd1 vccd1 vccd1 hold547/A sky130_fd_sc_hd__dfxtp_1
X_16888_ _18057_/CLK _16888_/D vssd1 vssd1 vccd1 vccd1 _16888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15839_ _17730_/CLK _15839_/D vssd1 vssd1 vccd1 vccd1 _15839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09360_ _09366_/A _09360_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09360_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08311_ _09313_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08311_/X sky130_fd_sc_hd__or2_1
X_17509_ _17509_/CLK _17509_/D vssd1 vssd1 vccd1 vccd1 _17509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09291_ _14972_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09291_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_13 _13116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _14461_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08242_/X sky130_fd_sc_hd__or2_1
XFILLER_0_144_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_24 _13180_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_35 _13260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 _15219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 hold484/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_wb_clk_i clkbuf_6_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17976_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08173_ _08504_/A _15182_/A vssd1 vssd1 vccd1 vccd1 _08173_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_68 hold597/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_79 _09313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5003 _11539_/X vssd1 vssd1 vccd1 vccd1 _17003_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5014 _16450_/Q vssd1 vssd1 vccd1 vccd1 hold5014/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5025 _13627_/X vssd1 vssd1 vccd1 vccd1 _17662_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5036 _17244_/Q vssd1 vssd1 vccd1 vccd1 hold5036/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4302 _13804_/Y vssd1 vssd1 vccd1 vccd1 _17721_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5047 _13453_/X vssd1 vssd1 vccd1 vccd1 _17604_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5058 _16854_/Q vssd1 vssd1 vccd1 vccd1 hold5058/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput120 hold5955/X vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_12
Xhold4313 _11751_/Y vssd1 vssd1 vccd1 vccd1 _11752_/B sky130_fd_sc_hd__dlygate4sd3_1
Xoutput131 hold5950/X vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_12
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4324 _12297_/Y vssd1 vssd1 vccd1 vccd1 _12298_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5069 _12286_/X vssd1 vssd1 vccd1 vccd1 _17252_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput142 hold935/X vssd1 vssd1 vccd1 vccd1 load_status[2] sky130_fd_sc_hd__buf_12
Xhold4335 _17566_/Q vssd1 vssd1 vccd1 vccd1 hold4335/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3601 _16421_/Q vssd1 vssd1 vccd1 vccd1 hold3601/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4346 _11730_/Y vssd1 vssd1 vccd1 vccd1 _11731_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3612 _16445_/Q vssd1 vssd1 vccd1 vccd1 hold3612/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4357 _11217_/Y vssd1 vssd1 vccd1 vccd1 _11218_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3623 _09562_/X vssd1 vssd1 vccd1 vccd1 _16344_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4368 _13872_/Y vssd1 vssd1 vccd1 vccd1 _13873_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3634 _16684_/Q vssd1 vssd1 vccd1 vccd1 hold3634/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4379 _13836_/Y vssd1 vssd1 vccd1 vccd1 _13837_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3645 _10102_/X vssd1 vssd1 vccd1 vccd1 _16524_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2900 _08463_/X vssd1 vssd1 vccd1 vccd1 _15860_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3656 _16342_/Q vssd1 vssd1 vccd1 vccd1 _13206_/A sky130_fd_sc_hd__buf_1
Xhold2911 _07953_/X vssd1 vssd1 vccd1 vccd1 _15619_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2922 _15844_/Q vssd1 vssd1 vccd1 vccd1 hold2922/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3667 _10390_/X vssd1 vssd1 vccd1 vccd1 _16620_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3678 _16378_/Q vssd1 vssd1 vccd1 vccd1 hold3678/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2933 _18397_/Q vssd1 vssd1 vccd1 vccd1 hold2933/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3689 _10186_/X vssd1 vssd1 vccd1 vccd1 _16552_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2944 _16271_/Q vssd1 vssd1 vccd1 vccd1 hold2944/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2955 _09213_/X vssd1 vssd1 vccd1 vccd1 _16218_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07957_ hold3095/X _07991_/A2 _07956_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _07957_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2966 _15693_/Q vssd1 vssd1 vccd1 vccd1 hold2966/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2977 _18249_/Q vssd1 vssd1 vccd1 vccd1 hold2977/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2988 _08400_/X vssd1 vssd1 vccd1 vccd1 _15830_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2999 _15719_/Q vssd1 vssd1 vccd1 vccd1 hold2999/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07888_ hold915/X _07936_/B vssd1 vssd1 vccd1 vccd1 _07888_/X sky130_fd_sc_hd__or2_1
XFILLER_0_214_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09627_ _11106_/A _09627_/B vssd1 vssd1 vccd1 vccd1 _09627_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09558_ _10386_/A _09558_/B vssd1 vssd1 vccd1 vccd1 _09558_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08509_ _15513_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08509_/X sky130_fd_sc_hd__or2_1
XFILLER_0_195_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09489_ _13048_/A _09489_/B vssd1 vssd1 vccd1 vccd1 _09494_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_210_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11520_ _11622_/A _11520_/B vssd1 vssd1 vccd1 vccd1 _11520_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11451_ _11655_/A _11451_/B vssd1 vssd1 vccd1 vccd1 _11451_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10402_ hold3257/X _10598_/B _10401_/X _15019_/C1 vssd1 vssd1 vccd1 vccd1 _10402_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14170_ _14974_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14170_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11382_ _11670_/A _11382_/B vssd1 vssd1 vccd1 vccd1 _11382_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13121_ _13121_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13121_/X sky130_fd_sc_hd__and2_1
X_10333_ hold3301/X _10637_/B _10332_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10333_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5570 _10960_/X vssd1 vssd1 vccd1 vccd1 _16810_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13052_ _17522_/Q _13056_/C _13056_/D _17523_/Q vssd1 vssd1 vccd1 vccd1 _13052_/X
+ sky130_fd_sc_hd__and4bb_4
X_10264_ hold4539/X _10628_/B _10263_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _10264_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5581 _17737_/Q vssd1 vssd1 vccd1 vccd1 hold5581/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5592 _11329_/X vssd1 vssd1 vccd1 vccd1 _16933_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12003_ _13797_/A _12003_/B vssd1 vssd1 vccd1 vccd1 _12003_/X sky130_fd_sc_hd__or2_1
Xhold4880 _13411_/X vssd1 vssd1 vccd1 vccd1 _17590_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10195_ hold3240/X _10577_/B _10194_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _10195_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4891 _16432_/Q vssd1 vssd1 vccd1 vccd1 hold4891/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_436_wb_clk_i clkbuf_6_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17425_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17860_ _17892_/CLK _17860_/D vssd1 vssd1 vccd1 vccd1 _17860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16811_ _18014_/CLK _16811_/D vssd1 vssd1 vccd1 vccd1 _16811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17791_ _17825_/CLK _17791_/D vssd1 vssd1 vccd1 vccd1 _17791_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout380 _14892_/B vssd1 vssd1 vccd1 vccd1 _14894_/B sky130_fd_sc_hd__buf_8
Xfanout391 _14680_/Y vssd1 vssd1 vccd1 vccd1 _14718_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13954_ _15515_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13954_/X sky130_fd_sc_hd__or2_1
X_16742_ _17949_/CLK _16742_/D vssd1 vssd1 vccd1 vccd1 _16742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_1259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12905_ hold3141/X _12904_/X _12905_/S vssd1 vssd1 vccd1 vccd1 _12905_/X sky130_fd_sc_hd__mux2_1
X_16673_ _18218_/CLK _16673_/D vssd1 vssd1 vccd1 vccd1 _16673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13885_ _13888_/A _13885_/B vssd1 vssd1 vccd1 vccd1 _13885_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_88_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18412_ _18412_/CLK _18412_/D vssd1 vssd1 vccd1 vccd1 _18412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12836_ hold4028/X _12835_/X _12839_/S vssd1 vssd1 vccd1 vccd1 _12836_/X sky130_fd_sc_hd__mux2_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15624_ _17878_/CLK _15624_/D vssd1 vssd1 vccd1 vccd1 _15624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18343_ _18375_/CLK _18343_/D vssd1 vssd1 vccd1 vccd1 _18343_/Q sky130_fd_sc_hd__dfxtp_1
X_15555_ _15555_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15555_/X sky130_fd_sc_hd__or2_1
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12767_ hold3813/X _12766_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12768_/B sky130_fd_sc_hd__mux2_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ hold2195/X _14537_/B _14505_/X _14372_/A vssd1 vssd1 vccd1 vccd1 _14506_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18274_ _18368_/CLK hold977/X vssd1 vssd1 vccd1 vccd1 _18274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11718_ hold3704/X _11622_/A _11717_/X vssd1 vssd1 vccd1 vccd1 _11718_/Y sky130_fd_sc_hd__a21oi_1
X_15486_ hold751/X _09367_/A _15486_/B1 hold845/X vssd1 vssd1 vccd1 vccd1 _15486_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12698_ hold3964/X _12697_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12699_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14437_ hold992/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14437_/X sky130_fd_sc_hd__or2_1
X_17225_ _18447_/CLK _17225_/D vssd1 vssd1 vccd1 vccd1 _17225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput11 input11/A vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_6
XFILLER_0_226_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11649_ _11649_/A _11649_/B vssd1 vssd1 vccd1 vccd1 _11649_/X sky130_fd_sc_hd__or2_1
Xinput22 input22/A vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_6
XFILLER_0_182_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput33 input33/A vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput44 input44/A vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_1
X_17156_ _17910_/CLK _17156_/D vssd1 vssd1 vccd1 vccd1 _17156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_226_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14368_ _14368_/A _14368_/B vssd1 vssd1 vccd1 vccd1 _17983_/D sky130_fd_sc_hd__and2_1
Xinput55 input55/A vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput66 input66/A vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__buf_6
XFILLER_0_3_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold806 hold806/A vssd1 vssd1 vccd1 vccd1 hold806/X sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ _16139_/CLK _16107_/D vssd1 vssd1 vccd1 vccd1 hold753/A sky130_fd_sc_hd__dfxtp_1
Xhold817 la_data_in[23] vssd1 vssd1 vccd1 vccd1 hold817/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 hold828/A vssd1 vssd1 vccd1 vccd1 hold828/X sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ hold2320/X _17560_/Q _13817_/C vssd1 vssd1 vccd1 vccd1 _13320_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_204_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold839 hold839/A vssd1 vssd1 vccd1 vccd1 hold839/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17087_ _18064_/CLK _17087_/D vssd1 vssd1 vccd1 vccd1 _17087_/Q sky130_fd_sc_hd__dfxtp_1
X_14299_ hold537/X _14333_/A2 _14298_/X _14364_/A vssd1 vssd1 vccd1 vccd1 hold538/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_228_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16038_ _16082_/CLK _16038_/D vssd1 vssd1 vccd1 vccd1 hold386/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08860_ hold87/X _16049_/Q _08860_/S vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_177_wb_clk_i clkbuf_6_49_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18375_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2207 _18226_/Q vssd1 vssd1 vccd1 vccd1 hold2207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2218 _17848_/Q vssd1 vssd1 vccd1 vccd1 hold2218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2229 _15784_/Q vssd1 vssd1 vccd1 vccd1 hold2229/X sky130_fd_sc_hd__dlygate4sd3_1
X_07811_ _13019_/A hold920/X hold892/X hold899/X vssd1 vssd1 vccd1 vccd1 _07811_/X
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_165_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1506 _15722_/Q vssd1 vssd1 vccd1 vccd1 hold1506/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_106_wb_clk_i clkbuf_6_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18401_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1517 _18044_/Q vssd1 vssd1 vccd1 vccd1 hold1517/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08791_ hold320/X _16016_/Q _08793_/S vssd1 vssd1 vccd1 vccd1 hold321/A sky130_fd_sc_hd__mux2_1
Xhold1528 _17511_/Q vssd1 vssd1 vccd1 vccd1 hold1528/X sky130_fd_sc_hd__dlygate4sd3_1
X_17989_ _18021_/CLK hold99/X vssd1 vssd1 vccd1 vccd1 _17989_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1539 _08259_/X vssd1 vssd1 vccd1 vccd1 _15764_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09412_ _09438_/B _09412_/B vssd1 vssd1 vccd1 vccd1 _09412_/X sky130_fd_sc_hd__or2_1
XFILLER_0_71_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09343_ _15559_/A _15231_/A hold353/A hold361/A vssd1 vssd1 vccd1 vccd1 _09352_/D
+ sky130_fd_sc_hd__or4_2
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09274_ _12753_/A _09274_/B vssd1 vssd1 vccd1 vccd1 _16248_/D sky130_fd_sc_hd__and2_1
XFILLER_0_63_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08225_ _15559_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08225_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08156_ hold444/X hold405/X hold337/X hold509/X vssd1 vssd1 vccd1 vccd1 _15492_/A
+ sky130_fd_sc_hd__and4b_4
XFILLER_0_31_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08087_ hold1287/X _08088_/B _08086_/Y _08145_/A vssd1 vssd1 vccd1 vccd1 _08087_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4110 _11302_/X vssd1 vssd1 vccd1 vccd1 _16924_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4121 _16690_/Q vssd1 vssd1 vccd1 vccd1 _10598_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4132 _11308_/X vssd1 vssd1 vccd1 vccd1 _16926_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4143 _16810_/Q vssd1 vssd1 vccd1 vccd1 hold4143/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4154 _17653_/Q vssd1 vssd1 vccd1 vccd1 hold4154/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3420 _16539_/Q vssd1 vssd1 vccd1 vccd1 hold3420/X sky130_fd_sc_hd__buf_1
Xhold4165 _16998_/Q vssd1 vssd1 vccd1 vccd1 hold4165/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3431 _10050_/Y vssd1 vssd1 vccd1 vccd1 _10051_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4176 _15481_/X vssd1 vssd1 vccd1 vccd1 _15482_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4187 hold5924/X vssd1 vssd1 vccd1 vccd1 hold5925/A sky130_fd_sc_hd__buf_4
Xhold3442 _16711_/Q vssd1 vssd1 vccd1 vccd1 hold3442/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4198 _15363_/X vssd1 vssd1 vccd1 vccd1 _15364_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3453 _17112_/Q vssd1 vssd1 vccd1 vccd1 hold3453/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3464 _10632_/Y vssd1 vssd1 vccd1 vccd1 _10633_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3475 hold6126/X vssd1 vssd1 vccd1 vccd1 hold3475/X sky130_fd_sc_hd__clkbuf_2
Xhold2730 _14279_/X vssd1 vssd1 vccd1 vccd1 _17940_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2741 _15837_/Q vssd1 vssd1 vccd1 vccd1 hold2741/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3486 _16526_/Q vssd1 vssd1 vccd1 vccd1 hold3486/X sky130_fd_sc_hd__buf_2
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08989_ hold82/X _16112_/Q _08991_/S vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__mux2_1
Xhold2752 _18338_/Q vssd1 vssd1 vccd1 vccd1 hold2752/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3497 _12366_/Y vssd1 vssd1 vccd1 vccd1 _12367_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2763 _08251_/X vssd1 vssd1 vccd1 vccd1 _15760_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2774 _14695_/X vssd1 vssd1 vccd1 vccd1 _18139_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2785 _17830_/Q vssd1 vssd1 vccd1 vccd1 hold2785/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2796 _18008_/Q vssd1 vssd1 vccd1 vccd1 hold2796/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10951_ hold3836/X _11144_/B _10950_/X _12978_/A vssd1 vssd1 vccd1 vccd1 _10951_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13670_ hold3078/X _17677_/Q _13766_/S vssd1 vssd1 vccd1 vccd1 _13671_/B sky130_fd_sc_hd__mux2_1
X_10882_ hold4167/X _11744_/B _10881_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _10882_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12621_ _12864_/A _12621_/B vssd1 vssd1 vccd1 vccd1 _12621_/X sky130_fd_sc_hd__and2_1
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15340_ hold599/X _09367_/A _09392_/A hold322/X vssd1 vssd1 vccd1 vccd1 _15340_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_241_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12552_ _12924_/A _12552_/B vssd1 vssd1 vccd1 vccd1 _17360_/D sky130_fd_sc_hd__and2_1
XPHY_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11503_ hold5309/X _11789_/B _11502_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _11503_/X
+ sky130_fd_sc_hd__o211a_1
X_15271_ _16291_/Q _09362_/A _15487_/B1 hold782/X _15270_/X vssd1 vssd1 vccd1 vccd1
+ _15272_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_191_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12483_ hold62/X _12509_/A2 _12501_/A3 _12482_/X _12410_/A vssd1 vssd1 vccd1 vccd1
+ hold63/A sky130_fd_sc_hd__o311a_1
XFILLER_0_108_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17010_ _17858_/CLK _17010_/D vssd1 vssd1 vccd1 vccd1 _17010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14222_ _14972_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14222_/X sky130_fd_sc_hd__or2_1
X_11434_ hold4173/X _11717_/B _11433_/X _12588_/A vssd1 vssd1 vccd1 vccd1 _11434_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14153_ hold2123/X _14148_/B _14152_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _14153_/X
+ sky130_fd_sc_hd__o211a_1
X_11365_ hold5370/X _11165_/B _11364_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _11365_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_4_wb_clk_i clkbuf_6_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18455_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13104_ _13097_/X _13103_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17531_/D sky130_fd_sc_hd__o21a_1
Xhold6090 la_data_in[14] vssd1 vssd1 vccd1 vccd1 hold627/A sky130_fd_sc_hd__dlygate4sd3_1
X_10316_ hold1766/X _16596_/Q _10604_/C vssd1 vssd1 vccd1 vccd1 _10317_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14084_ _15537_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14084_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11296_ hold5052/X _11771_/B _11295_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _11296_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_197_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13035_ _17523_/Q _13034_/X _13048_/A _13035_/D vssd1 vssd1 vccd1 vccd1 _13035_/X
+ sky130_fd_sc_hd__and4bb_1
X_17912_ _18073_/CLK _17912_/D vssd1 vssd1 vccd1 vccd1 _17912_/Q sky130_fd_sc_hd__dfxtp_1
X_10247_ hold1519/X hold3799/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10248_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_270_wb_clk_i clkbuf_6_57_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18124_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_238_1410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17843_ _17843_/CLK _17843_/D vssd1 vssd1 vccd1 vccd1 _17843_/Q sky130_fd_sc_hd__dfxtp_1
X_10178_ hold1652/X hold3740/X _10634_/C vssd1 vssd1 vccd1 vccd1 _10179_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_234_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17774_ _17774_/CLK hold299/X vssd1 vssd1 vccd1 vccd1 _17774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14986_ _15201_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14986_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16725_ _17960_/CLK _16725_/D vssd1 vssd1 vccd1 vccd1 _16725_/Q sky130_fd_sc_hd__dfxtp_1
X_13937_ _13943_/A _13937_/B vssd1 vssd1 vccd1 vccd1 _17776_/D sky130_fd_sc_hd__and2_1
XFILLER_0_88_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16656_ _18214_/CLK _16656_/D vssd1 vssd1 vccd1 vccd1 _16656_/Q sky130_fd_sc_hd__dfxtp_1
X_13868_ _17743_/Q _13868_/B _13868_/C vssd1 vssd1 vccd1 vccd1 _13868_/X sky130_fd_sc_hd__and3_1
XFILLER_0_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12819_ _12822_/A _12819_/B vssd1 vssd1 vccd1 vccd1 _17449_/D sky130_fd_sc_hd__and2_1
X_15607_ _18443_/CLK _15607_/D vssd1 vssd1 vccd1 vccd1 _15607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16587_ _18177_/CLK _16587_/D vssd1 vssd1 vccd1 vccd1 _16587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13799_ hold1175/X _17720_/Q _13817_/C vssd1 vssd1 vccd1 vccd1 _13800_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_226_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18326_ _18388_/CLK _18326_/D vssd1 vssd1 vccd1 vccd1 _18326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15538_ hold2179/X _15547_/B _15537_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _15538_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15469_ _17322_/Q _15487_/A2 _09392_/B hold688/X _15468_/X vssd1 vssd1 vccd1 vccd1
+ _15471_/C sky130_fd_sc_hd__a221o_1
X_18257_ _18327_/CLK _18257_/D vssd1 vssd1 vccd1 vccd1 _18257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08010_ hold1427/X _08029_/B _08009_/X _08167_/A vssd1 vssd1 vccd1 vccd1 _08010_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17208_ _17272_/CLK _17208_/D vssd1 vssd1 vccd1 vccd1 _17208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18188_ _18188_/CLK _18188_/D vssd1 vssd1 vccd1 vccd1 _18188_/Q sky130_fd_sc_hd__dfxtp_1
Xhold603 hold603/A vssd1 vssd1 vccd1 vccd1 hold603/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold614 hold614/A vssd1 vssd1 vccd1 vccd1 hold614/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_358_wb_clk_i clkbuf_6_41_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17576_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17139_ _17897_/CLK _17139_/D vssd1 vssd1 vccd1 vccd1 _17139_/Q sky130_fd_sc_hd__dfxtp_1
Xhold625 hold625/A vssd1 vssd1 vccd1 vccd1 hold625/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold636 hold636/A vssd1 vssd1 vccd1 vccd1 hold636/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 hold647/A vssd1 vssd1 vccd1 vccd1 hold647/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 hold658/A vssd1 vssd1 vccd1 vccd1 hold658/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09961_ hold3630/X _10601_/B _09960_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09961_/X
+ sky130_fd_sc_hd__o211a_1
Xhold669 hold669/A vssd1 vssd1 vccd1 vccd1 hold669/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08912_ hold373/X hold399/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08913_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_110_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09892_ hold5008/X _09992_/B _09891_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _09892_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2004 _17932_/Q vssd1 vssd1 vccd1 vccd1 hold2004/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2015 _17983_/Q vssd1 vssd1 vccd1 vccd1 hold2015/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2026 _14847_/X vssd1 vssd1 vccd1 vccd1 _18212_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08843_ _15364_/A _08843_/B vssd1 vssd1 vccd1 vccd1 _16040_/D sky130_fd_sc_hd__and2_1
Xhold2037 _18350_/Q vssd1 vssd1 vccd1 vccd1 hold2037/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2048 _14655_/X vssd1 vssd1 vccd1 vccd1 _18120_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1303 _15650_/Q vssd1 vssd1 vccd1 vccd1 hold1303/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1314 _14841_/X vssd1 vssd1 vccd1 vccd1 _18210_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2059 _14821_/X vssd1 vssd1 vccd1 vccd1 _18200_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1325 _15582_/Q vssd1 vssd1 vccd1 vccd1 hold1325/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1336 _15613_/Q vssd1 vssd1 vccd1 vccd1 hold1336/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08774_ _15482_/A _08774_/B vssd1 vssd1 vccd1 vccd1 _16007_/D sky130_fd_sc_hd__and2_1
XFILLER_0_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1347 _08006_/X vssd1 vssd1 vccd1 vccd1 _15644_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1358 _15663_/Q vssd1 vssd1 vccd1 vccd1 hold1358/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1369 _14345_/X vssd1 vssd1 vccd1 vccd1 _14346_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_74_wb_clk_i clkbuf_6_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18043_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_192_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09326_ hold961/X _09325_/B _09325_/Y _12906_/A vssd1 vssd1 vccd1 vccd1 hold962/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09257_ _15533_/A hold2459/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09258_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_211_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08208_ hold2749/X _08209_/B _08207_/Y _08381_/A vssd1 vssd1 vccd1 vccd1 _08208_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09188_ _15517_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09188_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_1307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08139_ _08139_/A hold623/X vssd1 vssd1 vccd1 vccd1 _15708_/D sky130_fd_sc_hd__and2_1
XFILLER_0_209_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11150_ _16874_/Q _11723_/B _11726_/C vssd1 vssd1 vccd1 vccd1 _11150_/X sky130_fd_sc_hd__and3_1
XTAP_6102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10101_ _10530_/A _10101_/B vssd1 vssd1 vccd1 vccd1 _10101_/X sky130_fd_sc_hd__or2_1
XTAP_6124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11081_ hold3019/X hold3808/X _11204_/C vssd1 vssd1 vccd1 vccd1 _11082_/B sky130_fd_sc_hd__mux2_1
XTAP_6146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3250 _09901_/X vssd1 vssd1 vccd1 vccd1 _16457_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3261 _16697_/Q vssd1 vssd1 vccd1 vccd1 hold3261/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10032_ _13198_/A _09948_/A _10031_/X vssd1 vssd1 vccd1 vccd1 _10032_/Y sky130_fd_sc_hd__a21oi_1
Xhold3272 _16601_/Q vssd1 vssd1 vccd1 vccd1 hold3272/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3283 _10387_/X vssd1 vssd1 vccd1 vccd1 _16619_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3294 _17376_/Q vssd1 vssd1 vccd1 vccd1 hold3294/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2560 _08320_/X vssd1 vssd1 vccd1 vccd1 _15793_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ _15233_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14840_/X sky130_fd_sc_hd__or2_1
Xhold2571 _16220_/Q vssd1 vssd1 vccd1 vccd1 hold2571/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2582 _15700_/Q vssd1 vssd1 vccd1 vccd1 hold2582/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2593 _17980_/Q vssd1 vssd1 vccd1 vccd1 hold2593/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1870 _15210_/X vssd1 vssd1 vccd1 vccd1 _18387_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1881 _18245_/Q vssd1 vssd1 vccd1 vccd1 hold1881/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14771_ hold2416/X _14774_/B _14770_/Y _15160_/C1 vssd1 vssd1 vccd1 vccd1 _14771_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_216_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11983_ hold4917/X _11798_/B _11982_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _11983_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1892 _14999_/X vssd1 vssd1 vccd1 vccd1 _18285_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16510_ _18393_/CLK _16510_/D vssd1 vssd1 vccd1 vccd1 _16510_/Q sky130_fd_sc_hd__dfxtp_1
X_13722_ _13722_/A _13722_/B vssd1 vssd1 vccd1 vccd1 _13722_/X sky130_fd_sc_hd__or2_1
X_10934_ hold2973/X _16802_/Q _11789_/C vssd1 vssd1 vccd1 vccd1 _10935_/B sky130_fd_sc_hd__mux2_1
X_17490_ _17492_/CLK _17490_/D vssd1 vssd1 vccd1 vccd1 _17490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_1362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16441_ _18380_/CLK _16441_/D vssd1 vssd1 vccd1 vccd1 _16441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13653_ _13788_/A _13653_/B vssd1 vssd1 vccd1 vccd1 _13653_/X sky130_fd_sc_hd__or2_1
X_10865_ hold2804/X hold4616/X _11153_/C vssd1 vssd1 vccd1 vccd1 _10866_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_128_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12604_ hold1499/X hold3263/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12604_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16372_ _18387_/CLK _16372_/D vssd1 vssd1 vccd1 vccd1 _16372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13584_ _13776_/A _13584_/B vssd1 vssd1 vccd1 vccd1 _13584_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ hold2151/X _16756_/Q _11186_/C vssd1 vssd1 vccd1 vccd1 _10797_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_27_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18111_ _18206_/CLK _18111_/D vssd1 vssd1 vccd1 vccd1 _18111_/Q sky130_fd_sc_hd__dfxtp_1
X_15323_ _15490_/A1 _15315_/X _15322_/X _15490_/B1 hold5918/A vssd1 vssd1 vccd1 vccd1
+ _15323_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_143_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ hold1706/X _17356_/Q _12925_/S vssd1 vssd1 vccd1 vccd1 _12535_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15254_ _15254_/A _15254_/B vssd1 vssd1 vccd1 vccd1 _18401_/D sky130_fd_sc_hd__and2_1
XFILLER_0_164_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18042_ _18042_/CLK _18042_/D vssd1 vssd1 vccd1 vccd1 _18042_/Q sky130_fd_sc_hd__dfxtp_1
X_12466_ _17326_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12466_/X sky130_fd_sc_hd__or2_1
XFILLER_0_22_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14205_ hold1231/X _14202_/B _14204_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _14205_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11417_ hold2597/X _16963_/Q _11774_/C vssd1 vssd1 vccd1 vccd1 _11418_/B sky130_fd_sc_hd__mux2_1
X_15185_ _15185_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15185_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_451_wb_clk_i clkbuf_6_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17721_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12397_ hold452/X hold839/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12398_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_22_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14136_ _14529_/A _14140_/B vssd1 vssd1 vccd1 vccd1 _14136_/X sky130_fd_sc_hd__or2_1
X_11348_ hold1658/X hold5293/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11349_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_10_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14067_ hold1233/X _14107_/A2 _14066_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _14067_/X
+ sky130_fd_sc_hd__o211a_1
X_11279_ _17765_/Q hold4384/X _11765_/C vssd1 vssd1 vccd1 vccd1 _11280_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_207_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13018_ hold2378/X _13003_/Y _13017_/X _12984_/A vssd1 vssd1 vccd1 vccd1 _13018_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17826_ _17858_/CLK _17826_/D vssd1 vssd1 vccd1 vccd1 _17826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17757_ _17886_/CLK _17757_/D vssd1 vssd1 vccd1 vccd1 _17757_/Q sky130_fd_sc_hd__dfxtp_1
X_14969_ hold1958/X _15004_/B _14968_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _14969_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16708_ _18073_/CLK _16708_/D vssd1 vssd1 vccd1 vccd1 _16708_/Q sky130_fd_sc_hd__dfxtp_1
X_08490_ _14543_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08490_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17688_ _17720_/CLK _17688_/D vssd1 vssd1 vccd1 vccd1 _17688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16639_ _18197_/CLK _16639_/D vssd1 vssd1 vccd1 vccd1 _16639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09111_ hold1974/X _09102_/B _09110_/X _12984_/A vssd1 vssd1 vccd1 vccd1 _09111_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18309_ _18349_/CLK _18309_/D vssd1 vssd1 vccd1 vccd1 _18309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09042_ hold373/X hold571/X _09060_/S vssd1 vssd1 vccd1 vccd1 _09043_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_192_wb_clk_i clkbuf_6_52_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18376_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold400 hold400/A vssd1 vssd1 vccd1 vccd1 hold400/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_241_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold411 hold411/A vssd1 vssd1 vccd1 vccd1 hold411/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold422 input64/X vssd1 vssd1 vccd1 vccd1 hold422/X sky130_fd_sc_hd__buf_1
Xhold433 hold433/A vssd1 vssd1 vccd1 vccd1 hold433/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_121_wb_clk_i clkbuf_6_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18425_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold444 hold444/A vssd1 vssd1 vccd1 vccd1 hold444/X sky130_fd_sc_hd__clkbuf_4
Xhold455 hold455/A vssd1 vssd1 vccd1 vccd1 hold455/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 hold466/A vssd1 vssd1 vccd1 vccd1 hold466/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold477 hold477/A vssd1 vssd1 vccd1 vccd1 hold477/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold488 hold488/A vssd1 vssd1 vccd1 vccd1 hold488/X sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ hold1821/X hold3880/X _11204_/C vssd1 vssd1 vccd1 vccd1 _09945_/B sky130_fd_sc_hd__mux2_1
Xfanout902 hold1367/X vssd1 vssd1 vccd1 vccd1 hold1368/A sky130_fd_sc_hd__buf_6
Xhold499 hold499/A vssd1 vssd1 vccd1 vccd1 hold499/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 _15173_/A vssd1 vssd1 vccd1 vccd1 _15553_/A sky130_fd_sc_hd__buf_12
XFILLER_0_42_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout924 hold1022/X vssd1 vssd1 vccd1 vccd1 _14970_/A sky130_fd_sc_hd__buf_4
XFILLER_0_239_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout935 hold1183/X vssd1 vssd1 vccd1 vccd1 _15209_/A sky130_fd_sc_hd__clkbuf_8
Xfanout946 hold1193/X vssd1 vssd1 vccd1 vccd1 _14395_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09875_ _18362_/Q _16449_/Q _10475_/S vssd1 vssd1 vccd1 vccd1 _09876_/B sky130_fd_sc_hd__mux2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1100 _08190_/X vssd1 vssd1 vccd1 vccd1 _15731_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 _15090_/X vssd1 vssd1 vccd1 vccd1 _18329_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ hold163/X hold461/X _08860_/S vssd1 vssd1 vccd1 vccd1 hold462/A sky130_fd_sc_hd__mux2_1
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 _09298_/X vssd1 vssd1 vccd1 vccd1 _16259_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1133 _09403_/X vssd1 vssd1 vccd1 vccd1 _16287_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 _08446_/X vssd1 vssd1 vccd1 vccd1 _15853_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1155 _18434_/Q vssd1 vssd1 vccd1 vccd1 hold1155/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1166 _15220_/X vssd1 vssd1 vccd1 vccd1 _18392_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08757_ hold169/X hold412/X _08779_/S vssd1 vssd1 vccd1 vccd1 hold413/A sky130_fd_sc_hd__mux2_1
Xhold1177 _18391_/Q vssd1 vssd1 vccd1 vccd1 hold1177/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1188 _15878_/Q vssd1 vssd1 vccd1 vccd1 hold1188/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1199 _18384_/Q vssd1 vssd1 vccd1 vccd1 hold1199/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08688_ _15244_/A hold415/X vssd1 vssd1 vccd1 vccd1 _15965_/D sky130_fd_sc_hd__and2_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10650_ hold3208/X _10470_/A _10649_/X vssd1 vssd1 vccd1 vccd1 _10650_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_193_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09309_ _14596_/A _09315_/B vssd1 vssd1 vccd1 vccd1 _09309_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10581_ hold3435/X _10530_/A _10580_/X vssd1 vssd1 vccd1 vccd1 _10581_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_181_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ _17264_/Q _12353_/B _13409_/S vssd1 vssd1 vccd1 vccd1 _12320_/X sky130_fd_sc_hd__and3_1
XFILLER_0_90_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_209_wb_clk_i clkbuf_6_55_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18396_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ hold2616/X hold5755/X _12362_/C vssd1 vssd1 vccd1 vccd1 _12252_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11202_ hold3450/X _11106_/A _11201_/X vssd1 vssd1 vccd1 vccd1 _11202_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12182_ hold1678/X _17218_/Q _13748_/S vssd1 vssd1 vccd1 vccd1 _12183_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_102_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11133_ _11637_/A _11133_/B vssd1 vssd1 vccd1 vccd1 _11133_/X sky130_fd_sc_hd__or2_1
X_16990_ _17774_/CLK _16990_/D vssd1 vssd1 vccd1 vccd1 _16990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15941_ _17288_/CLK _15941_/D vssd1 vssd1 vccd1 vccd1 hold769/A sky130_fd_sc_hd__dfxtp_1
X_11064_ _11067_/A _11064_/B vssd1 vssd1 vccd1 vccd1 _11064_/X sky130_fd_sc_hd__or2_1
XFILLER_0_235_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3080 _18357_/Q vssd1 vssd1 vccd1 vccd1 hold3080/X sky130_fd_sc_hd__dlygate4sd3_1
X_10015_ _11203_/A _10015_/B vssd1 vssd1 vccd1 vccd1 _10015_/Y sky130_fd_sc_hd__nor2_1
XTAP_5253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3091 _18004_/Q vssd1 vssd1 vccd1 vccd1 hold3091/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ _17608_/CLK _15872_/D vssd1 vssd1 vccd1 vccd1 _15872_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2390 _18242_/Q vssd1 vssd1 vccd1 vccd1 hold2390/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17611_ _17707_/CLK _17611_/D vssd1 vssd1 vccd1 vccd1 _17611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14823_ hold1754/X _14826_/B _14822_/Y _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14823_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17542_ _18352_/CLK _17542_/D vssd1 vssd1 vccd1 vccd1 _17542_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14754_ _15201_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14754_/X sky130_fd_sc_hd__or2_1
X_11966_ hold1056/X _17146_/Q _13463_/S vssd1 vssd1 vccd1 vccd1 _11967_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_231_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_230_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10917_ _11109_/A _10917_/B vssd1 vssd1 vccd1 vccd1 _10917_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13705_ hold5056/X _13814_/B _13704_/X _13801_/C1 vssd1 vssd1 vccd1 vccd1 _13705_/X
+ sky130_fd_sc_hd__o211a_1
X_14685_ hold1815/X _14720_/B _14684_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14685_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17473_ _17476_/CLK _17473_/D vssd1 vssd1 vccd1 vccd1 _17473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11897_ hold1112/X hold4320/X _13886_/C vssd1 vssd1 vccd1 vccd1 _11898_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16424_ _18373_/CLK _16424_/D vssd1 vssd1 vccd1 vccd1 _16424_/Q sky130_fd_sc_hd__dfxtp_1
X_13636_ hold4823/X _13862_/B _13635_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _13636_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_59_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_59_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_10848_ _11136_/A _10848_/B vssd1 vssd1 vccd1 vccd1 _10848_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16355_ _18298_/CLK _16355_/D vssd1 vssd1 vccd1 vccd1 _16355_/Q sky130_fd_sc_hd__dfxtp_1
X_13567_ hold5283/X _13874_/B _13566_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13567_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10779_ _11010_/A _10779_/B vssd1 vssd1 vccd1 vccd1 _10779_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15306_ _17334_/Q _09362_/C _09362_/D hold858/X vssd1 vssd1 vccd1 vccd1 _15306_/X
+ sky130_fd_sc_hd__a22o_1
X_12518_ hold4477/X _12517_/X _12929_/S vssd1 vssd1 vccd1 vccd1 _12518_/X sky130_fd_sc_hd__mux2_1
X_16286_ _17750_/CLK _16286_/D vssd1 vssd1 vccd1 vccd1 _16286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13498_ hold5595/X _13883_/B _13497_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13498_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18025_ _18222_/CLK _18025_/D vssd1 vssd1 vccd1 vccd1 _18025_/Q sky130_fd_sc_hd__dfxtp_1
X_15237_ _16132_/Q _15487_/A2 _15484_/B1 hold126/X _15236_/X vssd1 vssd1 vccd1 vccd1
+ _15242_/B sky130_fd_sc_hd__a221o_1
X_12449_ hold618/X _12509_/A2 _12501_/A3 _12448_/X _12418_/A vssd1 vssd1 vccd1 vccd1
+ hold135/A sky130_fd_sc_hd__o311a_1
Xhold4709 _17660_/Q vssd1 vssd1 vccd1 vccd1 hold4709/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_65_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15168_ hold2569/X _15167_/B _15167_/Y _15234_/C1 vssd1 vssd1 vccd1 vccd1 _15168_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14119_ hold2384/X _14142_/B _14118_/X _14346_/A vssd1 vssd1 vccd1 vccd1 _14119_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_227_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15099_ _15099_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15099_/X sky130_fd_sc_hd__or2_1
Xfanout209 fanout210/X vssd1 vssd1 vccd1 vccd1 _11792_/B sky130_fd_sc_hd__clkbuf_4
X_07990_ _14732_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07990_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09660_ _09948_/A _09660_/B vssd1 vssd1 vccd1 vccd1 _09660_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08611_ hold29/X hold207/X _08657_/S vssd1 vssd1 vccd1 vccd1 _08612_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_222_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17809_ _17843_/CLK _17809_/D vssd1 vssd1 vccd1 vccd1 _17809_/Q sky130_fd_sc_hd__dfxtp_1
X_09591_ _09957_/A _09591_/B vssd1 vssd1 vccd1 vccd1 _09591_/X sky130_fd_sc_hd__or2_1
XFILLER_0_206_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08542_ hold147/X hold659/X _08592_/S vssd1 vssd1 vccd1 vccd1 _08543_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_179_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08473_ hold1378/X _08486_/B _08472_/X _13765_/C1 vssd1 vssd1 vccd1 vccd1 _08473_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_373_wb_clk_i clkbuf_6_32_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17731_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_302_wb_clk_i clkbuf_6_44_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17898_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_143_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09025_ _15491_/A _09025_/B vssd1 vssd1 vccd1 vccd1 _16129_/D sky130_fd_sc_hd__and2_1
Xhold5900 _18407_/Q vssd1 vssd1 vccd1 vccd1 hold5900/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5911 _18404_/Q vssd1 vssd1 vccd1 vccd1 hold5911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5922 _18416_/Q vssd1 vssd1 vccd1 vccd1 hold5922/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5933 hold5933/A vssd1 vssd1 vccd1 vccd1 hold5933/X sky130_fd_sc_hd__buf_2
XFILLER_0_198_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5944 hold5944/A vssd1 vssd1 vccd1 vccd1 hold5944/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_182_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold230 hold230/A vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5955 hold5955/A vssd1 vssd1 vccd1 vccd1 hold5955/X sky130_fd_sc_hd__clkbuf_4
Xhold241 hold241/A vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 hold49/X vssd1 vssd1 vccd1 vccd1 input13/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5966 _18417_/Q vssd1 vssd1 vccd1 vccd1 hold5966/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5977 _13056_/C vssd1 vssd1 vccd1 vccd1 hold5977/X sky130_fd_sc_hd__buf_1
Xhold263 hold263/A vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5988 _16931_/Q vssd1 vssd1 vccd1 vccd1 hold5988/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 hold274/A vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5999 _16914_/Q vssd1 vssd1 vccd1 vccd1 hold5999/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 hold285/A vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 hold308/X vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__buf_1
Xfanout710 _12394_/A vssd1 vssd1 vccd1 vccd1 _15344_/A sky130_fd_sc_hd__clkbuf_4
Xfanout721 _15176_/C1 vssd1 vssd1 vccd1 vccd1 _14372_/A sky130_fd_sc_hd__buf_4
Xfanout732 _09907_/C1 vssd1 vssd1 vccd1 vccd1 _09003_/A sky130_fd_sc_hd__buf_2
X_09927_ _09981_/A _09927_/B vssd1 vssd1 vccd1 vccd1 _09927_/X sky130_fd_sc_hd__or2_1
XFILLER_0_141_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_217_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout743 fanout843/X vssd1 vssd1 vccd1 vccd1 _13675_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_233_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout754 _13929_/A vssd1 vssd1 vccd1 vccd1 _13933_/A sky130_fd_sc_hd__buf_4
Xfanout765 fanout791/X vssd1 vssd1 vccd1 vccd1 _13765_/C1 sky130_fd_sc_hd__buf_4
Xfanout776 _08149_/A vssd1 vssd1 vccd1 vccd1 _08153_/A sky130_fd_sc_hd__buf_4
X_09858_ _09954_/A _09858_/B vssd1 vssd1 vccd1 vccd1 _09858_/X sky130_fd_sc_hd__or2_1
Xfanout787 fanout791/X vssd1 vssd1 vccd1 vccd1 _13935_/A sky130_fd_sc_hd__buf_4
XFILLER_0_77_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_232_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout798 _15160_/C1 vssd1 vssd1 vccd1 vccd1 _15028_/A sky130_fd_sc_hd__buf_4
XFILLER_0_198_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _12420_/A hold137/X vssd1 vssd1 vccd1 vccd1 _16023_/D sky130_fd_sc_hd__and2_1
XFILLER_0_99_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _09981_/A _09789_/B vssd1 vssd1 vccd1 vccd1 _09789_/X sky130_fd_sc_hd__or2_1
XFILLER_0_38_1227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_103 _13294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11820_ _12210_/A _11820_/B vssd1 vssd1 vccd1 vccd1 _11820_/X sky130_fd_sc_hd__or2_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 hold915/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 _14988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ hold4312/X _11658_/A _11750_/X vssd1 vssd1 vccd1 vccd1 _11751_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_178_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10702_ hold5388/X _11186_/B _10701_/X _14462_/C1 vssd1 vssd1 vccd1 vccd1 _10702_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14470_ hold1487/X _14481_/B _14469_/X _14526_/C1 vssd1 vssd1 vccd1 vccd1 _14470_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11682_ _12285_/A _11682_/B vssd1 vssd1 vccd1 vccd1 _11682_/X sky130_fd_sc_hd__or2_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13421_ hold2979/X _17594_/Q _13721_/S vssd1 vssd1 vccd1 vccd1 _13422_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10633_ _10651_/A _10633_/B vssd1 vssd1 vccd1 vccd1 _16701_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16140_ _17520_/CLK _16140_/D vssd1 vssd1 vccd1 vccd1 hold138/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13352_ hold2899/X _17571_/Q _13766_/S vssd1 vssd1 vccd1 vccd1 _13353_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10564_ hold3893/X _10598_/B _10563_/X _10564_/C1 vssd1 vssd1 vccd1 vccd1 _16678_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_228_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12303_ hold4361/X _13716_/A _12302_/X vssd1 vssd1 vccd1 vccd1 _12303_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16071_ _17319_/CLK _16071_/D vssd1 vssd1 vccd1 vccd1 hold501/A sky130_fd_sc_hd__dfxtp_1
X_13283_ _13282_/X _16928_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13283_/X sky130_fd_sc_hd__mux2_1
X_10495_ _10589_/A _10589_/B _10494_/X _14691_/C1 vssd1 vssd1 vccd1 vccd1 _16655_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15022_ _15030_/A _15022_/B vssd1 vssd1 vccd1 vccd1 _18296_/D sky130_fd_sc_hd__and2_1
X_12234_ _12234_/A _12234_/B vssd1 vssd1 vccd1 vccd1 _12234_/X sky130_fd_sc_hd__or2_1
XFILLER_0_224_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12165_ _13482_/A _12165_/B vssd1 vssd1 vccd1 vccd1 _12165_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11116_ hold5247/X _11753_/B _11115_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11116_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12096_ _13314_/A _12096_/B vssd1 vssd1 vccd1 vccd1 _12096_/X sky130_fd_sc_hd__or2_1
X_16973_ _17853_/CLK _16973_/D vssd1 vssd1 vccd1 vccd1 _16973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15924_ _17300_/CLK _15924_/D vssd1 vssd1 vccd1 vccd1 hold625/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11047_ hold3868/X _11144_/B _11046_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _11047_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 input9/A vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_1
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _15856_/CLK _15855_/D vssd1 vssd1 vccd1 vccd1 _15855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14806_ _15145_/A _14830_/B vssd1 vssd1 vccd1 vccd1 _14806_/X sky130_fd_sc_hd__or2_1
XFILLER_0_188_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15786_ _17703_/CLK _15786_/D vssd1 vssd1 vccd1 vccd1 _15786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12998_ hold4965/X _12997_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12999_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_143_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17525_ _17525_/CLK _17525_/D vssd1 vssd1 vccd1 vccd1 _17525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14737_ hold2033/X _14772_/B _14736_/X _14853_/C1 vssd1 vssd1 vccd1 vccd1 _14737_/X
+ sky130_fd_sc_hd__o211a_1
X_11949_ _12255_/A _11949_/B vssd1 vssd1 vccd1 vccd1 _11949_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17456_ _17456_/CLK _17456_/D vssd1 vssd1 vccd1 vccd1 _17456_/Q sky130_fd_sc_hd__dfxtp_1
X_14668_ _15169_/A _14672_/B vssd1 vssd1 vccd1 vccd1 _14668_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16407_ _18352_/CLK _16407_/D vssd1 vssd1 vccd1 vccd1 _16407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13619_ hold2559/X hold4709/X _13811_/C vssd1 vssd1 vccd1 vccd1 _13620_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_229_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17387_ _18438_/CLK _17387_/D vssd1 vssd1 vccd1 vccd1 _17387_/Q sky130_fd_sc_hd__dfxtp_1
X_14599_ hold2287/X _14610_/B _14598_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14599_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16338_ _18383_/CLK _16338_/D vssd1 vssd1 vccd1 vccd1 _16338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5207 _17656_/Q vssd1 vssd1 vccd1 vccd1 hold5207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5218 _12181_/X vssd1 vssd1 vccd1 vccd1 _17217_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16269_ _17881_/CLK _16269_/D vssd1 vssd1 vccd1 vccd1 _16269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5229 _16676_/Q vssd1 vssd1 vccd1 vccd1 hold5229/X sky130_fd_sc_hd__dlygate4sd3_1
X_18008_ _18072_/CLK _18008_/D vssd1 vssd1 vccd1 vccd1 _18008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4506 _16931_/Q vssd1 vssd1 vccd1 vccd1 hold4506/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4517 _17357_/Q vssd1 vssd1 vccd1 vccd1 hold4517/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4528 _16485_/Q vssd1 vssd1 vccd1 vccd1 hold4528/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4539 _16610_/Q vssd1 vssd1 vccd1 vccd1 hold4539/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3805 _16659_/Q vssd1 vssd1 vccd1 vccd1 hold3805/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3816 _16561_/Q vssd1 vssd1 vccd1 vccd1 hold3816/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3827 _12713_/X vssd1 vssd1 vccd1 vccd1 _12714_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3838 _17603_/Q vssd1 vssd1 vccd1 vccd1 hold3838/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3849 _10468_/X vssd1 vssd1 vccd1 vccd1 _16646_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07973_ hold3053/X _07978_/B _07972_/Y _15502_/A vssd1 vssd1 vccd1 vccd1 _07973_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09712_ hold4693/X _11162_/B _09711_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _09712_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09643_ hold3602/X _10031_/B _09642_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09643_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_223_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09574_ hold3682/X _10052_/B _09573_/X _15019_/C1 vssd1 vssd1 vccd1 vccd1 _09574_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _15491_/A hold765/X vssd1 vssd1 vccd1 vccd1 _15887_/D sky130_fd_sc_hd__and2_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08456_ _14850_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08456_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08387_ _08387_/A _08387_/B vssd1 vssd1 vccd1 vccd1 _15825_/D sky130_fd_sc_hd__and2_1
XFILLER_0_34_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09008_ hold71/X hold280/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09009_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5730 _10017_/Y vssd1 vssd1 vccd1 vccd1 _10018_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10280_ hold2891/X hold3688/X _10571_/C vssd1 vssd1 vccd1 vccd1 _10281_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5741 _17145_/Q vssd1 vssd1 vccd1 vccd1 hold5741/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5752 _12169_/X vssd1 vssd1 vccd1 vccd1 _17213_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5763 _17627_/Q vssd1 vssd1 vccd1 vccd1 hold5763/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5774 _11884_/X vssd1 vssd1 vccd1 vccd1 _17118_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5785 _17182_/Q vssd1 vssd1 vccd1 vccd1 hold5785/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5796 _12133_/X vssd1 vssd1 vccd1 vccd1 _17201_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout540 _08860_/S vssd1 vssd1 vccd1 vccd1 _08866_/S sky130_fd_sc_hd__buf_8
Xfanout551 _08336_/A2 vssd1 vssd1 vccd1 vccd1 _08323_/B sky130_fd_sc_hd__buf_6
Xfanout562 _08048_/Y vssd1 vssd1 vccd1 vccd1 _08097_/A2 sky130_fd_sc_hd__buf_8
Xfanout573 _07871_/B vssd1 vssd1 vccd1 vccd1 _07881_/B sky130_fd_sc_hd__buf_8
X_13970_ _14596_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13970_/X sky130_fd_sc_hd__or2_1
Xfanout584 _13055_/X vssd1 vssd1 vccd1 vccd1 _13308_/S sky130_fd_sc_hd__buf_8
Xfanout595 _12871_/S vssd1 vssd1 vccd1 vccd1 _12850_/S sky130_fd_sc_hd__buf_6
X_12921_ _12924_/A _12921_/B vssd1 vssd1 vccd1 vccd1 _17483_/D sky130_fd_sc_hd__and2_1
XFILLER_0_9_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15640_ _17153_/CLK _15640_/D vssd1 vssd1 vccd1 vccd1 _15640_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _12855_/A _12852_/B vssd1 vssd1 vccd1 vccd1 _17460_/D sky130_fd_sc_hd__and2_1
XFILLER_0_232_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _12337_/A _11803_/B vssd1 vssd1 vccd1 vccd1 _11803_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_295_wb_clk_i clkbuf_6_39_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17964_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12783_ _12786_/A _12783_/B vssd1 vssd1 vccd1 vccd1 _17437_/D sky130_fd_sc_hd__and2_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _17271_/CLK _15571_/D vssd1 vssd1 vccd1 vccd1 _15571_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17310_ _18406_/CLK _17310_/D vssd1 vssd1 vccd1 vccd1 hold514/A sky130_fd_sc_hd__dfxtp_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14522_ hold2981/X _14541_/B _14521_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14522_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _12301_/A _11734_/B vssd1 vssd1 vccd1 vccd1 _17068_/D sky130_fd_sc_hd__nor2_1
X_18290_ _18356_/CLK hold512/X vssd1 vssd1 vccd1 vccd1 _18290_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_224_wb_clk_i clkbuf_6_63_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18197_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17241_ _17743_/CLK _17241_/D vssd1 vssd1 vccd1 vccd1 _17241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14453_ hold911/X _14499_/B vssd1 vssd1 vccd1 vccd1 _14453_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11665_ hold5259/X _11765_/B _11664_/X _14346_/A vssd1 vssd1 vccd1 vccd1 _11665_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10616_ _16696_/Q _10616_/B _11183_/C vssd1 vssd1 vccd1 vccd1 _10616_/X sky130_fd_sc_hd__and3_1
X_13404_ _13788_/A _13404_/B vssd1 vssd1 vccd1 vccd1 _13404_/X sky130_fd_sc_hd__or2_1
XFILLER_0_64_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14384_ _14388_/A _14384_/B vssd1 vssd1 vccd1 vccd1 _17991_/D sky130_fd_sc_hd__and2_1
XFILLER_0_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17172_ _17270_/CLK _17172_/D vssd1 vssd1 vccd1 vccd1 _17172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11596_ hold5257/X _12329_/B _11595_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11596_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16123_ _16147_/CLK _16123_/D vssd1 vssd1 vccd1 vccd1 hold327/A sky130_fd_sc_hd__dfxtp_1
X_13335_ _13722_/A _13335_/B vssd1 vssd1 vccd1 vccd1 _13335_/X sky130_fd_sc_hd__or2_1
XFILLER_0_84_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10547_ _18231_/Q _16673_/Q _10646_/C vssd1 vssd1 vccd1 vccd1 _10548_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16054_ _18401_/CLK _16054_/D vssd1 vssd1 vccd1 vccd1 hold797/A sky130_fd_sc_hd__dfxtp_1
X_13266_ _17584_/Q _17118_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13266_/X sky130_fd_sc_hd__mux2_1
X_10478_ hold2936/X hold4009/X _11186_/C vssd1 vssd1 vccd1 vccd1 _10479_/B sky130_fd_sc_hd__mux2_1
X_15005_ hold1432/X _15004_/B _15004_/Y _15146_/C1 vssd1 vssd1 vccd1 vccd1 _15005_/X
+ sky130_fd_sc_hd__o211a_1
X_12217_ _12311_/A _12217_/A2 _12216_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _12217_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13197_ _13196_/X hold3488/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13197_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_121_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12148_ hold5223/X _11771_/B _12147_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _12148_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_224_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12079_ hold4865/X _11798_/B _12078_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _12079_/X
+ sky130_fd_sc_hd__o211a_1
X_16956_ _17887_/CLK _16956_/D vssd1 vssd1 vccd1 vccd1 _16956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15907_ _16026_/CLK _15907_/D vssd1 vssd1 vccd1 vccd1 hold694/A sky130_fd_sc_hd__dfxtp_1
X_16887_ _18058_/CLK _16887_/D vssd1 vssd1 vccd1 vccd1 _16887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15838_ _17599_/CLK _15838_/D vssd1 vssd1 vccd1 vccd1 _15838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15769_ _17720_/CLK _15769_/D vssd1 vssd1 vccd1 vccd1 _15769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08310_ hold2857/X _08323_/B _08309_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _08310_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17508_ _17509_/CLK _17508_/D vssd1 vssd1 vccd1 vccd1 _17508_/Q sky130_fd_sc_hd__dfxtp_1
X_09290_ hold1242/X _09325_/B _09289_/X _12948_/A vssd1 vssd1 vccd1 vccd1 _09290_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08241_ hold1141/X _08262_/B _08240_/X _13765_/C1 vssd1 vssd1 vccd1 vccd1 _08241_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_14 _13116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17439_ _17446_/CLK _17439_/D vssd1 vssd1 vccd1 vccd1 _17439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_25 _13180_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_36 _13260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_47 _15201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_58 hold484/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ hold444/A hold405/A hold337/A hold509/A vssd1 vssd1 vccd1 vccd1 _15182_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_0_172_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_69 hold579/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5004 _17015_/Q vssd1 vssd1 vccd1 vccd1 hold5004/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5015 _09784_/X vssd1 vssd1 vccd1 vccd1 _16418_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5026 _16873_/Q vssd1 vssd1 vccd1 vccd1 hold5026/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_99_wb_clk_i clkbuf_6_22_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18405_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5037 _12166_/X vssd1 vssd1 vccd1 vccd1 _17212_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5048 _16618_/Q vssd1 vssd1 vccd1 vccd1 hold5048/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput110 hold5944/X vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_12
Xhold4303 _17575_/Q vssd1 vssd1 vccd1 vccd1 hold4303/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4314 _11752_/Y vssd1 vssd1 vccd1 vccd1 _17074_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5059 _10996_/X vssd1 vssd1 vccd1 vccd1 _16822_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput121 hold5957/X vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_12
XFILLER_0_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput132 hold5927/X vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_12
Xhold4325 _12298_/Y vssd1 vssd1 vccd1 vccd1 _17256_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput143 hold5977/X vssd1 vssd1 vccd1 vccd1 load_status[3] sky130_fd_sc_hd__buf_12
Xhold4336 _13819_/Y vssd1 vssd1 vccd1 vccd1 _17726_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_28_wb_clk_i clkbuf_6_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17476_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3602 _16403_/Q vssd1 vssd1 vccd1 vccd1 hold3602/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4347 _16735_/Q vssd1 vssd1 vccd1 vccd1 hold4347/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3613 _09769_/X vssd1 vssd1 vccd1 vccd1 _16413_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4358 _11218_/Y vssd1 vssd1 vccd1 vccd1 _16896_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3624 _17503_/Q vssd1 vssd1 vccd1 vccd1 hold3624/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4369 _13873_/Y vssd1 vssd1 vccd1 vccd1 _17744_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_227_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3635 _10486_/X vssd1 vssd1 vccd1 vccd1 _16652_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2901 _17976_/Q vssd1 vssd1 vccd1 vccd1 hold2901/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3646 _17630_/Q vssd1 vssd1 vccd1 vccd1 hold3646/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3657 _10035_/Y vssd1 vssd1 vccd1 vccd1 _10036_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2912 _15563_/Q vssd1 vssd1 vccd1 vccd1 hold2912/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3668 _16620_/Q vssd1 vssd1 vccd1 vccd1 hold3668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2923 _08428_/X vssd1 vssd1 vccd1 vccd1 _15844_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3679 _09568_/X vssd1 vssd1 vccd1 vccd1 _16346_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2934 _15230_/X vssd1 vssd1 vccd1 vccd1 _18397_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2945 _09322_/X vssd1 vssd1 vccd1 vccd1 _16271_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07956_ _15525_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07956_/X sky130_fd_sc_hd__or2_1
Xhold2956 _15782_/Q vssd1 vssd1 vccd1 vccd1 hold2956/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2967 _17829_/Q vssd1 vssd1 vccd1 vccd1 hold2967/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2978 _14925_/X vssd1 vssd1 vccd1 vccd1 _18249_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2989 _17835_/Q vssd1 vssd1 vccd1 vccd1 hold2989/X sky130_fd_sc_hd__dlygate4sd3_1
X_07887_ hold1562/X _07918_/B _07886_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _07887_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09626_ hold3072/X _16366_/Q _11201_/C vssd1 vssd1 vccd1 vccd1 _09627_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09557_ hold1211/X _13214_/A _10385_/S vssd1 vssd1 vccd1 vccd1 _09558_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_214_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08508_ hold1637/X _08503_/Y _08507_/X _08167_/A vssd1 vssd1 vccd1 vccd1 _08508_/X
+ sky130_fd_sc_hd__o211a_1
X_09488_ _17523_/Q _13035_/D vssd1 vssd1 vccd1 vccd1 _09489_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_182_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08439_ _15553_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08439_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11450_ hold1550/X _16974_/Q _11654_/S vssd1 vssd1 vccd1 vccd1 _11451_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_190_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10401_ _10539_/A _10401_/B vssd1 vssd1 vccd1 vccd1 _10401_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11381_ hold2455/X hold4887/X _11765_/C vssd1 vssd1 vccd1 vccd1 _11382_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ _13113_/X _13119_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17533_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_46_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10332_ _10542_/A _10332_/B vssd1 vssd1 vccd1 vccd1 _10332_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13051_ _13051_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13051_/X sky130_fd_sc_hd__and2_1
Xhold5560 _11827_/X vssd1 vssd1 vccd1 vccd1 _17099_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10263_ _10515_/A _10263_/B vssd1 vssd1 vccd1 vccd1 _10263_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5571 _17220_/Q vssd1 vssd1 vccd1 vccd1 hold5571/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5582 _13756_/X vssd1 vssd1 vccd1 vccd1 _17705_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5593 _17005_/Q vssd1 vssd1 vccd1 vccd1 hold5593/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12002_ hold1427/X hold4873/X _13796_/S vssd1 vssd1 vccd1 vccd1 _12003_/B sky130_fd_sc_hd__mux2_1
Xhold4870 _11068_/X vssd1 vssd1 vccd1 vccd1 _16846_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10194_ _10386_/A _10194_/B vssd1 vssd1 vccd1 vccd1 _10194_/X sky130_fd_sc_hd__or2_1
Xhold4881 _16895_/Q vssd1 vssd1 vccd1 vccd1 hold4881/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4892 _09730_/X vssd1 vssd1 vccd1 vccd1 _16400_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16810_ _17981_/CLK _16810_/D vssd1 vssd1 vccd1 vccd1 _16810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17790_ _17886_/CLK _17790_/D vssd1 vssd1 vccd1 vccd1 _17790_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout370 hold340/X vssd1 vssd1 vccd1 vccd1 hold341/A sky130_fd_sc_hd__buf_6
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout381 hold331/X vssd1 vssd1 vccd1 vccd1 hold332/A sky130_fd_sc_hd__buf_6
Xfanout392 _14672_/B vssd1 vssd1 vccd1 vccd1 _14678_/B sky130_fd_sc_hd__buf_6
X_16741_ _17976_/CLK _16741_/D vssd1 vssd1 vccd1 vccd1 _16741_/Q sky130_fd_sc_hd__dfxtp_1
X_13953_ hold3063/X _13995_/A2 _13952_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _13953_/X
+ sky130_fd_sc_hd__o211a_1
X_12904_ hold2464/X _17479_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12904_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_202_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16672_ _18231_/CLK _16672_/D vssd1 vssd1 vccd1 vccd1 _16672_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_405_wb_clk_i clkbuf_6_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17885_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13884_ hold4488/X _13788_/A _13883_/X vssd1 vssd1 vccd1 vccd1 _13884_/Y sky130_fd_sc_hd__a21oi_1
X_18411_ _18411_/CLK _18411_/D vssd1 vssd1 vccd1 vccd1 _18411_/Q sky130_fd_sc_hd__dfxtp_1
X_15623_ _17187_/CLK _15623_/D vssd1 vssd1 vccd1 vccd1 _15623_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12835_ hold2809/X _17456_/Q _12838_/S vssd1 vssd1 vccd1 vccd1 _12835_/X sky130_fd_sc_hd__mux2_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _18342_/CLK _18342_/D vssd1 vssd1 vccd1 vccd1 _18342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ hold2756/X _15560_/A2 _15553_/X _12843_/A vssd1 vssd1 vccd1 vccd1 _15554_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12766_ hold954/X hold3570/X _12766_/S vssd1 vssd1 vccd1 vccd1 _12766_/X sky130_fd_sc_hd__mux2_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14505_ _14970_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14505_/X sky130_fd_sc_hd__or2_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18273_ _18373_/CLK _18273_/D vssd1 vssd1 vccd1 vccd1 _18273_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11717_ _17063_/Q _11717_/B _11717_/C vssd1 vssd1 vccd1 vccd1 _11717_/X sky130_fd_sc_hd__and3_1
X_15485_ hold300/X _15485_/A2 _15485_/B1 hold256/X vssd1 vssd1 vccd1 vccd1 _15485_/X
+ sky130_fd_sc_hd__a22o_1
X_12697_ hold2564/X hold3793/X _12766_/S vssd1 vssd1 vccd1 vccd1 _12697_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_140_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17224_ _18443_/CLK _17224_/D vssd1 vssd1 vccd1 vccd1 _17224_/Q sky130_fd_sc_hd__dfxtp_1
X_14436_ hold1964/X _14433_/B _14435_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _14436_/X
+ sky130_fd_sc_hd__o211a_1
X_11648_ _17888_/Q hold4040/X _11738_/C vssd1 vssd1 vccd1 vccd1 _11649_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_4_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput12 input12/A vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_6
XFILLER_0_142_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput23 input23/A vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_1
XFILLER_0_226_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput34 input34/A vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput45 input45/A vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_2
X_17155_ _17735_/CLK _17155_/D vssd1 vssd1 vccd1 vccd1 _17155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14367_ _15535_/A hold2015/X _14381_/S vssd1 vssd1 vccd1 vccd1 _14367_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11579_ hold3068/X hold4149/X _12242_/S vssd1 vssd1 vccd1 vccd1 _11580_/B sky130_fd_sc_hd__mux2_1
Xinput56 input56/A vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_2
Xhold807 hold807/A vssd1 vssd1 vccd1 vccd1 hold807/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput67 input67/A vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16106_ _18405_/CLK _16106_/D vssd1 vssd1 vccd1 vccd1 hold398/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold818 hold818/A vssd1 vssd1 vccd1 vccd1 input52/A sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ hold4781/X _12308_/B _13317_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _13318_/X
+ sky130_fd_sc_hd__o211a_1
Xhold829 hold829/A vssd1 vssd1 vccd1 vccd1 hold829/X sky130_fd_sc_hd__dlygate4sd3_1
X_17086_ _17774_/CLK _17086_/D vssd1 vssd1 vccd1 vccd1 _17086_/Q sky130_fd_sc_hd__dfxtp_1
X_14298_ hold423/X _14338_/B vssd1 vssd1 vccd1 vccd1 _14298_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16037_ _17293_/CLK _16037_/D vssd1 vssd1 vccd1 vccd1 hold661/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13249_ _13249_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13249_/X sky130_fd_sc_hd__and2_1
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2208 _14875_/X vssd1 vssd1 vccd1 vccd1 _18226_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2219 _14087_/X vssd1 vssd1 vccd1 vccd1 _17848_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07810_ _15274_/A _17751_/Q vssd1 vssd1 vccd1 vccd1 _07810_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08790_ _15482_/A hold566/X vssd1 vssd1 vccd1 vccd1 _16015_/D sky130_fd_sc_hd__and2_1
Xhold1507 hold6107/X vssd1 vssd1 vccd1 vccd1 _09447_/C sky130_fd_sc_hd__clkbuf_2
Xhold1518 _14494_/X vssd1 vssd1 vccd1 vccd1 _18044_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17988_ _18050_/CLK hold152/X vssd1 vssd1 vccd1 vccd1 _17988_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1529 _13006_/X vssd1 vssd1 vccd1 vccd1 _17511_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16939_ _17883_/CLK _16939_/D vssd1 vssd1 vccd1 vccd1 _16939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_146_wb_clk_i clkbuf_6_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18423_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09411_ _07804_/A _09447_/A _09440_/B _09410_/X vssd1 vssd1 vccd1 vccd1 _09411_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09342_ _09342_/A _09342_/B vssd1 vssd1 vccd1 vccd1 _09342_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_90_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09273_ _15549_/A hold1264/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09274_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08224_ hold1672/X _08209_/B _08223_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _08224_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08155_ _08163_/A _08155_/B vssd1 vssd1 vccd1 vccd1 _15716_/D sky130_fd_sc_hd__and2_1
XFILLER_0_114_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_222_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08086_ _15219_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08086_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_141_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4100 _11038_/X vssd1 vssd1 vccd1 vccd1 _16836_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4111 _16932_/Q vssd1 vssd1 vccd1 vccd1 hold4111/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4122 _10504_/X vssd1 vssd1 vccd1 vccd1 _16658_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4133 hold5926/X vssd1 vssd1 vccd1 vccd1 hold5927/A sky130_fd_sc_hd__buf_4
XTAP_6306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4144 _10864_/X vssd1 vssd1 vccd1 vccd1 _16778_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3410 _10048_/Y vssd1 vssd1 vccd1 vccd1 _16506_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4155 _13504_/X vssd1 vssd1 vccd1 vccd1 _17621_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3421 _10626_/Y vssd1 vssd1 vccd1 vccd1 _10627_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4166 _11428_/X vssd1 vssd1 vccd1 vccd1 _16966_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3432 _16350_/Q vssd1 vssd1 vccd1 vccd1 _13270_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4177 _17063_/Q vssd1 vssd1 vccd1 vccd1 hold4177/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4188 _15303_/X vssd1 vssd1 vccd1 vccd1 _15304_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3443 _11142_/Y vssd1 vssd1 vccd1 vccd1 _11143_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3454 _12345_/Y vssd1 vssd1 vccd1 vccd1 _12346_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4199 hold5900/X vssd1 vssd1 vccd1 vccd1 hold4199/X sky130_fd_sc_hd__clkbuf_4
XTAP_5627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2720 _09093_/X vssd1 vssd1 vccd1 vccd1 _16161_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3465 _16922_/Q vssd1 vssd1 vccd1 vccd1 hold3465/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2731 _17924_/Q vssd1 vssd1 vccd1 vccd1 hold2731/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3476 _16737_/Q vssd1 vssd1 vccd1 vccd1 hold3476/X sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_5649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3487 _10587_/Y vssd1 vssd1 vccd1 vccd1 _10588_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2742 _08414_/X vssd1 vssd1 vccd1 vccd1 _15837_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2753 _15108_/X vssd1 vssd1 vccd1 vccd1 _18338_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08988_ _15314_/A _08988_/B vssd1 vssd1 vccd1 vccd1 _16111_/D sky130_fd_sc_hd__and2_1
Xhold3498 _12367_/Y vssd1 vssd1 vccd1 vccd1 _17279_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2764 _17761_/Q vssd1 vssd1 vccd1 vccd1 hold2764/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2775 _15661_/Q vssd1 vssd1 vccd1 vccd1 hold2775/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07939_ _14735_/A hold355/X vssd1 vssd1 vccd1 vccd1 _07990_/B sky130_fd_sc_hd__or2_4
Xhold2786 _14049_/X vssd1 vssd1 vccd1 vccd1 _17830_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2797 _14420_/X vssd1 vssd1 vccd1 vccd1 _18008_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10950_ _11049_/A _10950_/B vssd1 vssd1 vccd1 vccd1 _10950_/X sky130_fd_sc_hd__or2_1
XFILLER_0_211_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09609_ _09987_/A _09609_/B vssd1 vssd1 vccd1 vccd1 _09609_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10881_ _11649_/A _10881_/B vssd1 vssd1 vccd1 vccd1 _10881_/X sky130_fd_sc_hd__or2_1
XFILLER_0_6_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ _17383_/Q _12619_/X _12626_/S vssd1 vssd1 vccd1 vccd1 _12620_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12551_ hold4552/X _12550_/X _12929_/S vssd1 vssd1 vccd1 vccd1 _12551_/X sky130_fd_sc_hd__mux2_1
XPHY_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11502_ _11694_/A _11502_/B vssd1 vssd1 vccd1 vccd1 _11502_/X sky130_fd_sc_hd__or2_1
X_12482_ _17334_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12482_/X sky130_fd_sc_hd__or2_1
X_15270_ hold666/X _09367_/A _15446_/B1 hold874/X vssd1 vssd1 vccd1 vccd1 _15270_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14221_ hold2163/X _14216_/Y _14220_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _14221_/X
+ sky130_fd_sc_hd__o211a_1
X_11433_ _11622_/A _11433_/B vssd1 vssd1 vccd1 vccd1 _11433_/X sky130_fd_sc_hd__or2_1
XFILLER_0_117_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14152_ hold992/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14152_/X sky130_fd_sc_hd__or2_1
XFILLER_0_145_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11364_ _11556_/A _11364_/B vssd1 vssd1 vccd1 vccd1 _11364_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6080 _18264_/Q vssd1 vssd1 vccd1 vccd1 hold6080/X sky130_fd_sc_hd__dlygate4sd3_1
X_10315_ hold3781/X _10637_/B _10314_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10315_/X
+ sky130_fd_sc_hd__o211a_1
X_13103_ _13199_/A1 _13101_/X _13102_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13103_/X
+ sky130_fd_sc_hd__o211a_1
Xhold6091 _16283_/Q vssd1 vssd1 vccd1 vccd1 hold6091/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14083_ hold2079/X _14094_/B _14082_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _14083_/X
+ sky130_fd_sc_hd__o211a_1
X_11295_ _12243_/A _11295_/B vssd1 vssd1 vccd1 vccd1 _11295_/X sky130_fd_sc_hd__or2_1
X_13034_ hold907/X _13056_/C _17520_/Q _13034_/D vssd1 vssd1 vccd1 vccd1 _13034_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_123_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17911_ _18073_/CLK _17911_/D vssd1 vssd1 vccd1 vccd1 _17911_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5390 _16942_/Q vssd1 vssd1 vccd1 vccd1 hold5390/X sky130_fd_sc_hd__dlygate4sd3_1
X_10246_ hold4456/X _10628_/B _10245_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10246_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17842_ _17874_/CLK _17842_/D vssd1 vssd1 vccd1 vccd1 _17842_/Q sky130_fd_sc_hd__dfxtp_1
X_10177_ hold3550/X _10601_/B _10176_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _10177_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_238_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_234_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17773_ _17774_/CLK _17773_/D vssd1 vssd1 vccd1 vccd1 _17773_/Q sky130_fd_sc_hd__dfxtp_1
X_14985_ hold3102/X _15004_/B _14984_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _14985_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16724_ _17964_/CLK _16724_/D vssd1 vssd1 vccd1 vccd1 _16724_/Q sky130_fd_sc_hd__dfxtp_1
X_13936_ _14330_/A hold1486/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13937_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16655_ _18213_/CLK _16655_/D vssd1 vssd1 vccd1 vccd1 _16655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13867_ _13873_/A _13867_/B vssd1 vssd1 vccd1 vccd1 _13867_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_187_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15606_ _15886_/CLK _15606_/D vssd1 vssd1 vccd1 vccd1 _15606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12818_ hold3380/X _12817_/X _12839_/S vssd1 vssd1 vccd1 vccd1 _12819_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_158_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16586_ _18176_/CLK _16586_/D vssd1 vssd1 vccd1 vccd1 _16586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ hold4743/X _12308_/B _13797_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _13798_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18325_ _18325_/CLK _18325_/D vssd1 vssd1 vccd1 vccd1 _18325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15537_ _15537_/A _15549_/B vssd1 vssd1 vccd1 vccd1 _15537_/X sky130_fd_sc_hd__or2_1
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ hold3175/X _12748_/X _12749_/S vssd1 vssd1 vccd1 vccd1 _12749_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18256_ _18384_/CLK _18256_/D vssd1 vssd1 vccd1 vccd1 _18256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15468_ hold302/X _09367_/A _09362_/C hold136/X vssd1 vssd1 vccd1 vccd1 _15468_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_231_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17207_ _17271_/CLK _17207_/D vssd1 vssd1 vccd1 vccd1 _17207_/Q sky130_fd_sc_hd__dfxtp_1
X_14419_ _15099_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14419_/X sky130_fd_sc_hd__or2_1
XFILLER_0_115_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18187_ _18233_/CLK _18187_/D vssd1 vssd1 vccd1 vccd1 _18187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15399_ hold634/X _09365_/B _09392_/C hold773/X _15398_/X vssd1 vssd1 vccd1 vccd1
+ _15402_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_25_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold604 hold604/A vssd1 vssd1 vccd1 vccd1 hold604/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17138_ _17209_/CLK _17138_/D vssd1 vssd1 vccd1 vccd1 _17138_/Q sky130_fd_sc_hd__dfxtp_1
Xhold615 data_in[1] vssd1 vssd1 vccd1 vccd1 hold615/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 hold626/A vssd1 vssd1 vccd1 vccd1 hold626/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold637 hold637/A vssd1 vssd1 vccd1 vccd1 hold637/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 hold648/A vssd1 vssd1 vccd1 vccd1 hold648/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold659 hold659/A vssd1 vssd1 vccd1 vccd1 hold659/X sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ _10482_/A _09960_/B vssd1 vssd1 vccd1 vccd1 _09960_/X sky130_fd_sc_hd__or2_1
X_17069_ _17885_/CLK _17069_/D vssd1 vssd1 vccd1 vccd1 _17069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08911_ _15434_/A hold284/X vssd1 vssd1 vccd1 vccd1 _16073_/D sky130_fd_sc_hd__and2_1
XFILLER_0_228_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09891_ _09987_/A _09891_/B vssd1 vssd1 vccd1 vccd1 _09891_/X sky130_fd_sc_hd__or2_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_398_wb_clk_i clkbuf_6_36_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17838_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2005 _14263_/X vssd1 vssd1 vccd1 vccd1 _17932_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2016 _14367_/X vssd1 vssd1 vccd1 vccd1 _14368_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2027 _18198_/Q vssd1 vssd1 vccd1 vccd1 hold2027/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08842_ hold215/X hold601/X _08866_/S vssd1 vssd1 vccd1 vccd1 _08843_/B sky130_fd_sc_hd__mux2_1
Xhold2038 _15134_/X vssd1 vssd1 vccd1 vccd1 _18350_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1304 _08018_/X vssd1 vssd1 vccd1 vccd1 _15650_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_327_wb_clk_i clkbuf_6_44_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17873_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2049 _18147_/Q vssd1 vssd1 vccd1 vccd1 hold2049/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1315 _18255_/Q vssd1 vssd1 vccd1 vccd1 hold1315/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1326 _07874_/X vssd1 vssd1 vccd1 vccd1 _15582_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_236_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08773_ hold373/X hold400/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08774_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1337 _07941_/X vssd1 vssd1 vccd1 vccd1 _15613_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1348 _18039_/Q vssd1 vssd1 vccd1 vccd1 hold1348/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1359 _08044_/X vssd1 vssd1 vccd1 vccd1 _15663_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09325_ _14952_/A _09325_/B vssd1 vssd1 vccd1 vccd1 _09325_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_164_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09256_ _12753_/A _09256_/B vssd1 vssd1 vccd1 vccd1 _16239_/D sky130_fd_sc_hd__and2_1
XFILLER_0_209_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08207_ _15215_/A _08209_/B vssd1 vssd1 vccd1 vccd1 _08207_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_105_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_43_wb_clk_i clkbuf_6_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17884_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_106_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09187_ hold3000/X _09218_/B _09186_/X _12843_/A vssd1 vssd1 vccd1 vccd1 _09187_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08138_ hold597/X hold622/X hold108/X vssd1 vssd1 vccd1 vccd1 hold623/A sky130_fd_sc_hd__mux2_1
XFILLER_0_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08069_ hold2662/X _08097_/A2 _08068_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _08069_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10100_ hold1730/X hold3435/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10101_/B sky130_fd_sc_hd__mux2_1
XTAP_6114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11080_ hold4957/X _11753_/B _11079_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _11080_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3240 _16587_/Q vssd1 vssd1 vccd1 vccd1 hold3240/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10031_ _16501_/Q _10031_/B _10031_/C vssd1 vssd1 vccd1 vccd1 _10031_/X sky130_fd_sc_hd__and3_1
Xhold3251 _16667_/Q vssd1 vssd1 vccd1 vccd1 hold3251/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3262 _10525_/X vssd1 vssd1 vccd1 vccd1 _16665_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3273 _10237_/X vssd1 vssd1 vccd1 vccd1 _16569_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3284 _16619_/Q vssd1 vssd1 vccd1 vccd1 hold3284/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2550 _18366_/Q vssd1 vssd1 vccd1 vccd1 hold2550/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3295 _17373_/Q vssd1 vssd1 vccd1 vccd1 hold3295/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2561 _18306_/Q vssd1 vssd1 vccd1 vccd1 hold2561/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2572 _09217_/X vssd1 vssd1 vccd1 vccd1 _16220_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2583 _18182_/Q vssd1 vssd1 vccd1 vccd1 hold2583/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2594 _18099_/Q vssd1 vssd1 vccd1 vccd1 hold2594/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1860 _14021_/X vssd1 vssd1 vccd1 vccd1 _17816_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1871 _18149_/Q vssd1 vssd1 vccd1 vccd1 hold1871/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14770_ _15163_/A _14774_/B vssd1 vssd1 vccd1 vccd1 _14770_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1882 _14917_/X vssd1 vssd1 vccd1 vccd1 _18245_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ _12174_/A _11982_/B vssd1 vssd1 vccd1 vccd1 _11982_/X sky130_fd_sc_hd__or2_1
Xhold1893 _18072_/Q vssd1 vssd1 vccd1 vccd1 hold1893/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13721_ hold1471/X _17694_/Q _13721_/S vssd1 vssd1 vccd1 vccd1 _13722_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10933_ hold4705/X _11765_/B _10932_/X _14346_/A vssd1 vssd1 vccd1 vccd1 _10933_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_1374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16440_ _18321_/CLK _16440_/D vssd1 vssd1 vccd1 vccd1 _16440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13652_ hold1935/X _17671_/Q _13874_/C vssd1 vssd1 vccd1 vccd1 _13653_/B sky130_fd_sc_hd__mux2_1
X_10864_ hold4143/X _11723_/B _10863_/X _14364_/A vssd1 vssd1 vccd1 vccd1 _10864_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_49_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_49_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ _12612_/A _12603_/B vssd1 vssd1 vccd1 vccd1 _17377_/D sky130_fd_sc_hd__and2_1
X_16371_ _18342_/CLK _16371_/D vssd1 vssd1 vccd1 vccd1 _16371_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ hold4945/X _11171_/B _10794_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _10795_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ hold1049/X hold5150/X _13865_/C vssd1 vssd1 vccd1 vccd1 _13584_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18110_ _18265_/CLK _18110_/D vssd1 vssd1 vccd1 vccd1 _18110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15322_ _15489_/A _15322_/B _15322_/C _15322_/D vssd1 vssd1 vccd1 vccd1 _15322_/X
+ sky130_fd_sc_hd__or4_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _12948_/A _12534_/B vssd1 vssd1 vccd1 vccd1 _17354_/D sky130_fd_sc_hd__and2_1
XFILLER_0_26_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18041_ _18041_/CLK _18041_/D vssd1 vssd1 vccd1 vccd1 _18041_/Q sky130_fd_sc_hd__dfxtp_1
X_15253_ _15490_/A1 _15245_/X _15252_/X _15490_/B1 hold5916/A vssd1 vssd1 vccd1 vccd1
+ _15253_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_41_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12465_ hold673/X _08597_/Y _12501_/A3 _12464_/X _12420_/A vssd1 vssd1 vccd1 vccd1
+ hold75/A sky130_fd_sc_hd__o311a_1
XFILLER_0_227_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14204_ _14543_/A _14204_/B vssd1 vssd1 vccd1 vccd1 _14204_/X sky130_fd_sc_hd__or2_1
X_11416_ hold4789/X _11798_/B _11415_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _11416_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15184_ hold1968/X _15219_/B _15183_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _15184_/X
+ sky130_fd_sc_hd__o211a_1
X_12396_ _15274_/A hold889/X vssd1 vssd1 vccd1 vccd1 _17291_/D sky130_fd_sc_hd__and2_1
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14135_ hold1558/X _14142_/B _14134_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _14135_/X
+ sky130_fd_sc_hd__o211a_1
X_11347_ hold5191/X _11726_/B _11346_/X _13895_/A vssd1 vssd1 vccd1 vccd1 _11347_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14066_ _15085_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14066_/X sky130_fd_sc_hd__or2_1
X_11278_ hold5633/X _11786_/B _11277_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _11278_/X
+ sky130_fd_sc_hd__o211a_1
X_10229_ hold2689/X hold3328/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10230_/B sky130_fd_sc_hd__mux2_1
X_13017_ _14980_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13017_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_420_wb_clk_i clkbuf_6_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17157_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17825_ _17825_/CLK _17825_/D vssd1 vssd1 vccd1 vccd1 _17825_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_234_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17756_ _17820_/CLK _17756_/D vssd1 vssd1 vccd1 vccd1 _17756_/Q sky130_fd_sc_hd__dfxtp_1
X_14968_ hold927/X _15018_/B vssd1 vssd1 vccd1 vccd1 _14968_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16707_ _18233_/CLK _16707_/D vssd1 vssd1 vccd1 vccd1 _16707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13919_ _13935_/A _13919_/B vssd1 vssd1 vccd1 vccd1 _13919_/X sky130_fd_sc_hd__and2_1
X_17687_ _17719_/CLK _17687_/D vssd1 vssd1 vccd1 vccd1 _17687_/Q sky130_fd_sc_hd__dfxtp_1
X_14899_ hold2177/X _14896_/Y _14898_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _14899_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16638_ _18228_/CLK _16638_/D vssd1 vssd1 vccd1 vccd1 _16638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16569_ _18191_/CLK _16569_/D vssd1 vssd1 vccd1 vccd1 _16569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09110_ hold992/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09110_/X sky130_fd_sc_hd__or2_1
X_18308_ _18308_/CLK _18308_/D vssd1 vssd1 vccd1 vccd1 _18308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09041_ _12438_/A _09041_/B vssd1 vssd1 vccd1 vccd1 _16137_/D sky130_fd_sc_hd__and2_1
X_18239_ _18411_/CLK _18239_/D vssd1 vssd1 vccd1 vccd1 _18239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold401 hold401/A vssd1 vssd1 vccd1 vccd1 hold401/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold412 hold412/A vssd1 vssd1 vccd1 vccd1 hold412/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold423 hold423/A vssd1 vssd1 vccd1 vccd1 hold423/X sky130_fd_sc_hd__buf_6
Xhold434 hold434/A vssd1 vssd1 vccd1 vccd1 hold434/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold445 hold445/A vssd1 vssd1 vccd1 vccd1 hold445/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold456 hold456/A vssd1 vssd1 vccd1 vccd1 hold456/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold467 hold467/A vssd1 vssd1 vccd1 vccd1 hold467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 hold478/A vssd1 vssd1 vccd1 vccd1 hold478/X sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ hold3632/X _10049_/B _09942_/X _15212_/C1 vssd1 vssd1 vccd1 vccd1 _09943_/X
+ sky130_fd_sc_hd__o211a_1
Xhold489 hold489/A vssd1 vssd1 vccd1 vccd1 hold489/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout903 hold1367/X vssd1 vssd1 vccd1 vccd1 _15187_/A sky130_fd_sc_hd__buf_4
XFILLER_0_106_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout914 _15173_/A vssd1 vssd1 vccd1 vccd1 _14726_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout925 hold1022/X vssd1 vssd1 vccd1 vccd1 hold915/A sky130_fd_sc_hd__buf_6
XFILLER_0_238_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout936 _15207_/A vssd1 vssd1 vccd1 vccd1 _15533_/A sky130_fd_sc_hd__buf_12
XFILLER_0_42_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09874_ hold3950/X _10046_/B _09873_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09874_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_161_wb_clk_i clkbuf_6_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18411_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout947 hold1193/X vssd1 vssd1 vccd1 vccd1 hold927/A sky130_fd_sc_hd__buf_6
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 _17948_/Q vssd1 vssd1 vccd1 vccd1 hold1101/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1112 _15715_/Q vssd1 vssd1 vccd1 vccd1 hold1112/X sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ _15344_/A _08825_/B vssd1 vssd1 vccd1 vccd1 _16031_/D sky130_fd_sc_hd__and2_1
Xhold1123 _15729_/Q vssd1 vssd1 vccd1 vccd1 hold1123/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1134 _15825_/Q vssd1 vssd1 vccd1 vccd1 hold1134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 la_data_in[12] vssd1 vssd1 vccd1 vccd1 hold1145/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1156 _15512_/X vssd1 vssd1 vccd1 vccd1 _18434_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1167 _17812_/Q vssd1 vssd1 vccd1 vccd1 hold1167/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08756_ _15414_/A _08756_/B vssd1 vssd1 vccd1 vccd1 _15998_/D sky130_fd_sc_hd__and2_1
Xhold1178 _15218_/X vssd1 vssd1 vccd1 vccd1 _18391_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1189 _08499_/X vssd1 vssd1 vccd1 vccd1 _15878_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ hold163/X hold414/X _08721_/S vssd1 vssd1 vccd1 vccd1 hold415/A sky130_fd_sc_hd__mux2_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09308_ hold2767/X _09323_/B _09307_/X _14358_/A vssd1 vssd1 vccd1 vccd1 _09308_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10580_ _16684_/Q _10625_/B _10625_/C vssd1 vssd1 vccd1 vccd1 _10580_/X sky130_fd_sc_hd__and3_1
XFILLER_0_10_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09239_ _15515_/A hold2524/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09240_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12250_ hold4987/X _12374_/B _12249_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _12250_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11201_ _16891_/Q _11201_/B _11201_/C vssd1 vssd1 vccd1 vccd1 _11201_/X sky130_fd_sc_hd__and3_1
X_12181_ hold5217/X _12374_/B _12180_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _12181_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_249_wb_clk_i clkbuf_6_59_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18166_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11132_ _18071_/Q hold4099/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11133_/B sky130_fd_sc_hd__mux2_1
Xhold990 input50/X vssd1 vssd1 vccd1 vccd1 hold990/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_102_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15940_ _18410_/CLK _15940_/D vssd1 vssd1 vccd1 vccd1 hold539/A sky130_fd_sc_hd__dfxtp_1
XTAP_5210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11063_ hold2133/X _16845_/Q _11162_/C vssd1 vssd1 vccd1 vccd1 _11064_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_229_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3070 _16157_/Q vssd1 vssd1 vccd1 vccd1 hold3070/X sky130_fd_sc_hd__dlygate4sd3_1
X_10014_ _13150_/A _11061_/A _10013_/X vssd1 vssd1 vccd1 vccd1 _10014_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3081 _15148_/X vssd1 vssd1 vccd1 vccd1 _18357_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3092 _14412_/X vssd1 vssd1 vccd1 vccd1 _18004_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15871_ _17584_/CLK _15871_/D vssd1 vssd1 vccd1 vccd1 _15871_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2380 _18100_/Q vssd1 vssd1 vccd1 vccd1 hold2380/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ _17738_/CLK _17610_/D vssd1 vssd1 vccd1 vccd1 _17610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14822_ _15161_/A _14826_/B vssd1 vssd1 vccd1 vccd1 _14822_/Y sky130_fd_sc_hd__nand2_1
XTAP_5298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2391 _14909_/X vssd1 vssd1 vccd1 vccd1 _18242_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17541_ _18386_/CLK _17541_/D vssd1 vssd1 vccd1 vccd1 _17541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1690 _16197_/Q vssd1 vssd1 vccd1 vccd1 hold1690/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14753_ hold2236/X _14774_/B _14752_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14753_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ hold5765/X _12350_/B _11964_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _11965_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13704_ _13800_/A _13704_/B vssd1 vssd1 vccd1 vccd1 _13704_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10916_ hold3169/X hold4819/X _11204_/C vssd1 vssd1 vccd1 vccd1 _10917_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_86_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17472_ _17477_/CLK _17472_/D vssd1 vssd1 vccd1 vccd1 _17472_/Q sky130_fd_sc_hd__dfxtp_1
X_14684_ _15185_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14684_/X sky130_fd_sc_hd__or2_1
XFILLER_0_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11896_ hold5331/X _12374_/B _11895_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _11896_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16423_ _18398_/CLK _16423_/D vssd1 vssd1 vccd1 vccd1 _16423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_1299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ _13737_/A _13635_/B vssd1 vssd1 vccd1 vccd1 _13635_/X sky130_fd_sc_hd__or2_1
XFILLER_0_89_1318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10847_ hold2901/X hold4995/X _11153_/C vssd1 vssd1 vccd1 vccd1 _10848_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_172_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16354_ _18395_/CLK _16354_/D vssd1 vssd1 vccd1 vccd1 _16354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13566_ _13758_/A _13566_/B vssd1 vssd1 vccd1 vccd1 _13566_/X sky130_fd_sc_hd__or2_1
XFILLER_0_41_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10778_ hold1674/X _16750_/Q _11171_/C vssd1 vssd1 vccd1 vccd1 _10779_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_125_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15305_ hold877/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15305_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12517_ hold1811/X _17350_/Q _12925_/S vssd1 vssd1 vccd1 vccd1 _12517_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16285_ _17750_/CLK _16285_/D vssd1 vssd1 vccd1 vccd1 _16285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13497_ _13788_/A _13497_/B vssd1 vssd1 vccd1 vccd1 _13497_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18024_ _18024_/CLK _18024_/D vssd1 vssd1 vccd1 vccd1 _18024_/Q sky130_fd_sc_hd__dfxtp_1
X_15236_ _17327_/Q _15486_/B1 _15485_/B1 _16104_/Q vssd1 vssd1 vccd1 vccd1 _15236_/X
+ sky130_fd_sc_hd__a22o_1
X_12448_ _17317_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12448_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15167_ _15547_/A _15167_/B vssd1 vssd1 vccd1 vccd1 _15167_/Y sky130_fd_sc_hd__nand2_1
X_12379_ _13888_/A _12379_/B vssd1 vssd1 vccd1 vccd1 _12379_/Y sky130_fd_sc_hd__nor2_1
X_14118_ _14457_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14118_/X sky130_fd_sc_hd__or2_1
X_15098_ hold2191/X hold340/X _15097_/X _15202_/C1 vssd1 vssd1 vccd1 vccd1 _15098_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_197_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14049_ hold2785/X _14040_/B _14048_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14049_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08610_ _12420_/A _08610_/B vssd1 vssd1 vccd1 vccd1 _15927_/D sky130_fd_sc_hd__and2_1
XFILLER_0_179_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09590_ hold1299/X _13302_/A _10040_/C vssd1 vssd1 vccd1 vccd1 _09591_/B sky130_fd_sc_hd__mux2_1
X_17808_ _17840_/CLK _17808_/D vssd1 vssd1 vccd1 vccd1 _17808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_234_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08541_ _09057_/A _08541_/B vssd1 vssd1 vccd1 vccd1 _15894_/D sky130_fd_sc_hd__and2_1
X_17739_ _17739_/CLK _17739_/D vssd1 vssd1 vccd1 vccd1 _17739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08472_ _15531_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08472_/X sky130_fd_sc_hd__or2_1
XFILLER_0_159_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09024_ hold77/X hold256/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09025_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_143_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5901 hold6036/X vssd1 vssd1 vccd1 vccd1 _13051_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_60_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5912 hold5912/A vssd1 vssd1 vccd1 vccd1 hold5912/X sky130_fd_sc_hd__buf_2
XFILLER_0_108_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5923 hold5923/A vssd1 vssd1 vccd1 vccd1 hold5923/X sky130_fd_sc_hd__buf_2
XFILLER_0_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5934 _18405_/Q vssd1 vssd1 vccd1 vccd1 hold5934/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold220 hold220/A vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__buf_6
XFILLER_0_41_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5945 _18409_/Q vssd1 vssd1 vccd1 vccd1 hold5945/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5956 _18422_/Q vssd1 vssd1 vccd1 vccd1 hold5956/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold231 hold231/A vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_342_wb_clk_i clkbuf_6_42_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17703_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold242 hold242/A vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5967 hold5967/A vssd1 vssd1 vccd1 vccd1 hold5967/X sky130_fd_sc_hd__clkbuf_4
Xhold253 input13/X vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5978 _18459_/Q vssd1 vssd1 vccd1 vccd1 hold5978/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 hold264/A vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5989 _16310_/Q vssd1 vssd1 vccd1 vccd1 hold5989/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 hold275/A vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout700 _08851_/A vssd1 vssd1 vccd1 vccd1 _09440_/B sky130_fd_sc_hd__buf_4
Xhold286 hold286/A vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 hold297/A vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__clkbuf_16
Xfanout711 fanout739/X vssd1 vssd1 vccd1 vccd1 _12394_/A sky130_fd_sc_hd__buf_2
Xfanout722 _15404_/A vssd1 vssd1 vccd1 vccd1 _15394_/A sky130_fd_sc_hd__buf_4
X_09926_ hold2948/X hold4849/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09927_/B sky130_fd_sc_hd__mux2_1
Xfanout733 _08954_/A vssd1 vssd1 vccd1 vccd1 _15482_/A sky130_fd_sc_hd__buf_4
Xfanout744 _08111_/A vssd1 vssd1 vccd1 vccd1 _08139_/A sky130_fd_sc_hd__buf_4
Xfanout755 _14131_/C1 vssd1 vssd1 vccd1 vccd1 _13929_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout766 fanout791/X vssd1 vssd1 vccd1 vccd1 _08391_/A sky130_fd_sc_hd__buf_2
X_09857_ hold2259/X _16443_/Q _10049_/C vssd1 vssd1 vccd1 vccd1 _09858_/B sky130_fd_sc_hd__mux2_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout777 fanout791/X vssd1 vssd1 vccd1 vccd1 _08149_/A sky130_fd_sc_hd__clkbuf_4
Xfanout788 fanout791/X vssd1 vssd1 vccd1 vccd1 _14546_/C1 sky130_fd_sc_hd__buf_2
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout799 _15160_/C1 vssd1 vssd1 vccd1 vccd1 _14388_/A sky130_fd_sc_hd__buf_4
XFILLER_0_137_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ hold131/X hold136/X _08866_/S vssd1 vssd1 vccd1 vccd1 hold137/A sky130_fd_sc_hd__mux2_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09788_ hold2191/X hold4042/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09789_/B sky130_fd_sc_hd__mux2_1
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ hold71/X hold300/X _08779_/S vssd1 vssd1 vccd1 vccd1 _08740_/B sky130_fd_sc_hd__mux2_1
XANTENNA_104 _13294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 hold915/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_126 hold915/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _17074_/Q _11753_/B _11753_/C vssd1 vssd1 vccd1 vccd1 _11750_/X sky130_fd_sc_hd__and3_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10701_ _11661_/A _10701_/B vssd1 vssd1 vccd1 vccd1 _10701_/X sky130_fd_sc_hd__or2_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ hold1362/X _17051_/Q _12317_/C vssd1 vssd1 vccd1 vccd1 _11682_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_37_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13420_ hold4831/X _13814_/B _13419_/X _08361_/A vssd1 vssd1 vccd1 vccd1 _13420_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10632_ hold3463/X _10536_/A _10631_/X vssd1 vssd1 vccd1 vccd1 _10632_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_193_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10563_ _10563_/A _10563_/B vssd1 vssd1 vccd1 vccd1 _10563_/X sky130_fd_sc_hd__or2_1
XFILLER_0_148_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13351_ hold4664/X _13829_/B _13350_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13351_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12302_ _17258_/Q _13811_/B _13811_/C vssd1 vssd1 vccd1 vccd1 _12302_/X sky130_fd_sc_hd__and3_1
XFILLER_0_228_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16070_ _18417_/CLK _16070_/D vssd1 vssd1 vccd1 vccd1 hold426/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_1368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10494_ _10554_/A _10494_/B vssd1 vssd1 vccd1 vccd1 _10494_/X sky130_fd_sc_hd__or2_1
X_13282_ _17586_/Q _17120_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13282_/X sky130_fd_sc_hd__mux2_1
X_15021_ _15183_/A hold1483/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15022_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12233_ hold2426/X hold5675/X _12242_/S vssd1 vssd1 vccd1 vccd1 _12234_/B sky130_fd_sc_hd__mux2_1
X_12164_ hold2840/X hold4749/X _13481_/S vssd1 vssd1 vccd1 vccd1 _12165_/B sky130_fd_sc_hd__mux2_1
X_11115_ _11658_/A _11115_/B vssd1 vssd1 vccd1 vccd1 _11115_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12095_ hold2828/X hold4970/X _13409_/S vssd1 vssd1 vccd1 vccd1 _12096_/B sky130_fd_sc_hd__mux2_1
X_16972_ _17884_/CLK _16972_/D vssd1 vssd1 vccd1 vccd1 _16972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15923_ _16090_/CLK _15923_/D vssd1 vssd1 vccd1 vccd1 hold767/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11046_ _11049_/A _11046_/B vssd1 vssd1 vccd1 vccd1 _11046_/X sky130_fd_sc_hd__or2_1
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _17630_/CLK _15854_/D vssd1 vssd1 vccd1 vccd1 _15854_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14805_ hold1265/X _14828_/B _14804_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14805_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15785_ _17716_/CLK _15785_/D vssd1 vssd1 vccd1 vccd1 _15785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12997_ hold2060/X hold4760/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12997_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17524_ _17525_/CLK hold924/X vssd1 vssd1 vccd1 vccd1 _17524_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ _15183_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14736_/X sky130_fd_sc_hd__or2_1
XFILLER_0_143_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11948_ hold1544/X _17140_/Q _13463_/S vssd1 vssd1 vccd1 vccd1 _11949_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17455_ _17456_/CLK _17455_/D vssd1 vssd1 vccd1 vccd1 _17455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ hold2351/X _14666_/B _14666_/Y _14344_/A vssd1 vssd1 vccd1 vccd1 _14667_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11879_ _15709_/Q hold5708/X _12362_/C vssd1 vssd1 vccd1 vccd1 _11880_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_184_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16406_ _18383_/CLK _16406_/D vssd1 vssd1 vccd1 vccd1 _16406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13618_ hold4660/X _13814_/B _13617_/X _12753_/A vssd1 vssd1 vccd1 vccd1 _13618_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17386_ _18438_/CLK _17386_/D vssd1 vssd1 vccd1 vccd1 _17386_/Q sky130_fd_sc_hd__dfxtp_1
X_14598_ _15099_/A _14622_/B vssd1 vssd1 vccd1 vccd1 _14598_/X sky130_fd_sc_hd__or2_1
XFILLER_0_172_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16337_ _18378_/CLK _16337_/D vssd1 vssd1 vccd1 vccd1 _16337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13549_ hold5319/X _13856_/B _13548_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13549_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16268_ _18013_/CLK _16268_/D vssd1 vssd1 vccd1 vccd1 _16268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5208 _13513_/X vssd1 vssd1 vccd1 vccd1 _17624_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5219 _16859_/Q vssd1 vssd1 vccd1 vccd1 hold5219/X sky130_fd_sc_hd__dlygate4sd3_1
X_18007_ _18039_/CLK _18007_/D vssd1 vssd1 vccd1 vccd1 _18007_/Q sky130_fd_sc_hd__dfxtp_1
X_15219_ _15219_/A _15219_/B vssd1 vssd1 vccd1 vccd1 _15219_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_207_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4507 _11802_/Y vssd1 vssd1 vccd1 vccd1 _11803_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4518 _12542_/X vssd1 vssd1 vccd1 vccd1 _12543_/B sky130_fd_sc_hd__dlygate4sd3_1
X_16199_ _17484_/CLK _16199_/D vssd1 vssd1 vccd1 vccd1 _16199_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4529 _09889_/X vssd1 vssd1 vccd1 vccd1 _16453_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3806 _10411_/X vssd1 vssd1 vccd1 vccd1 _16627_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3817 _10117_/X vssd1 vssd1 vccd1 vccd1 _16529_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3828 _16744_/Q vssd1 vssd1 vccd1 vccd1 hold3828/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3839 _13354_/X vssd1 vssd1 vccd1 vccd1 _17571_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07972_ _15541_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _07972_/Y sky130_fd_sc_hd__nand2_1
X_09711_ _11067_/A _09711_/B vssd1 vssd1 vccd1 vccd1 _09711_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09642_ _09948_/A _09642_/B vssd1 vssd1 vccd1 vccd1 _09642_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09573_ _09957_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09573_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ hold226/X hold764/X _08528_/S vssd1 vssd1 vccd1 vccd1 hold765/A sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08455_ hold2983/X _08488_/B _08454_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _08455_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08386_ _14960_/A hold1134/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08386_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_107_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09007_ _12440_/A hold836/X vssd1 vssd1 vccd1 vccd1 _16120_/D sky130_fd_sc_hd__and2_1
Xhold5720 _17562_/Q vssd1 vssd1 vccd1 vccd1 hold5720/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5731 _17170_/Q vssd1 vssd1 vccd1 vccd1 hold5731/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5742 _11869_/X vssd1 vssd1 vccd1 vccd1 _17113_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5753 _16338_/Q vssd1 vssd1 vccd1 vccd1 _13174_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5764 _13426_/X vssd1 vssd1 vccd1 vccd1 _17595_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5775 _17210_/Q vssd1 vssd1 vccd1 vccd1 hold5775/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5786 _11980_/X vssd1 vssd1 vccd1 vccd1 _17150_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5797 _17689_/Q vssd1 vssd1 vccd1 vccd1 hold5797/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout530 _09218_/B vssd1 vssd1 vccd1 vccd1 _09214_/B sky130_fd_sc_hd__clkbuf_8
Xfanout541 _08858_/S vssd1 vssd1 vccd1 vccd1 _08860_/S sky130_fd_sc_hd__buf_8
X_09909_ _09984_/A _09909_/B vssd1 vssd1 vccd1 vccd1 _09909_/X sky130_fd_sc_hd__or2_1
Xfanout552 _08283_/Y vssd1 vssd1 vccd1 vccd1 _08336_/A2 sky130_fd_sc_hd__buf_8
Xfanout563 _08048_/Y vssd1 vssd1 vccd1 vccd1 _08088_/B sky130_fd_sc_hd__clkbuf_8
Xfanout574 _07829_/Y vssd1 vssd1 vccd1 vccd1 _07865_/B sky130_fd_sc_hd__buf_6
Xfanout585 _13294_/B vssd1 vssd1 vccd1 vccd1 _13302_/B sky130_fd_sc_hd__buf_6
Xfanout596 _12871_/S vssd1 vssd1 vccd1 vccd1 _12916_/S sky130_fd_sc_hd__buf_6
X_12920_ hold3355/X _12919_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12921_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_88_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ hold3149/X _12850_/X _12851_/S vssd1 vssd1 vccd1 vccd1 _12851_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_197_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ hold4506/X _12240_/A _11801_/X vssd1 vssd1 vccd1 vccd1 _11802_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _17204_/CLK _15570_/D vssd1 vssd1 vccd1 vccd1 _15570_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ hold4036/X _12781_/X _12839_/S vssd1 vssd1 vccd1 vccd1 _12783_/B sky130_fd_sc_hd__mux2_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14521_ _15201_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14521_/X sky130_fd_sc_hd__or2_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11733_ hold4419/X _11637_/A _11732_/X vssd1 vssd1 vccd1 vccd1 _11733_/Y sky130_fd_sc_hd__a21oi_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17240_ _17272_/CLK _17240_/D vssd1 vssd1 vccd1 vccd1 _17240_/Q sky130_fd_sc_hd__dfxtp_1
X_14452_ hold2066/X _14481_/B _14451_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _14452_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11664_ _11670_/A _11664_/B vssd1 vssd1 vccd1 vccd1 _11664_/X sky130_fd_sc_hd__or2_1
XFILLER_0_83_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13403_ hold1497/X hold4488/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13404_/B sky130_fd_sc_hd__mux2_1
X_10615_ _10651_/A _10615_/B vssd1 vssd1 vccd1 vccd1 _16695_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_3_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17171_ _17897_/CLK _17171_/D vssd1 vssd1 vccd1 vccd1 _17171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_264_wb_clk_i clkbuf_6_56_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18057_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14383_ _15225_/A hold1955/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14384_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_37_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11595_ _12234_/A _11595_/B vssd1 vssd1 vccd1 vccd1 _11595_/X sky130_fd_sc_hd__or2_1
X_16122_ _17341_/CLK _16122_/D vssd1 vssd1 vccd1 vccd1 hold665/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13334_ hold1647/X _17565_/Q _13721_/S vssd1 vssd1 vccd1 vccd1 _13335_/B sky130_fd_sc_hd__mux2_1
X_10546_ hold4579/X _10649_/B _10545_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _10546_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16053_ _17284_/CLK _16053_/D vssd1 vssd1 vccd1 vccd1 hold647/A sky130_fd_sc_hd__dfxtp_1
X_13265_ _13265_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13265_/X sky130_fd_sc_hd__and2_1
XFILLER_0_165_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10477_ _10571_/A _10568_/B _10476_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _10477_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15004_ _15219_/A _15004_/B vssd1 vssd1 vccd1 vccd1 _15004_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_121_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12216_ _12216_/A _12216_/B vssd1 vssd1 vccd1 vccd1 _12216_/X sky130_fd_sc_hd__or2_1
X_13196_ hold3490/X _13195_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13196_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_62_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12147_ _12243_/A _12147_/B vssd1 vssd1 vccd1 vccd1 _12147_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_236_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12078_ _12174_/A _12078_/B vssd1 vssd1 vccd1 vccd1 _12078_/X sky130_fd_sc_hd__or2_1
X_16955_ _17823_/CLK _16955_/D vssd1 vssd1 vccd1 vccd1 _16955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_236_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15906_ _17324_/CLK _15906_/D vssd1 vssd1 vccd1 vccd1 hold745/A sky130_fd_sc_hd__dfxtp_1
X_11029_ hold3858/X _11765_/B _11028_/X _14346_/A vssd1 vssd1 vccd1 vccd1 _11029_/X
+ sky130_fd_sc_hd__o211a_1
X_16886_ _17929_/CLK _16886_/D vssd1 vssd1 vccd1 vccd1 _16886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_8_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_8_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15837_ _17728_/CLK _15837_/D vssd1 vssd1 vccd1 vccd1 _15837_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_232_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_235_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15768_ _17718_/CLK _15768_/D vssd1 vssd1 vccd1 vccd1 _15768_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14719_ hold2587/X _14718_/B _14718_/Y _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14719_/X
+ sky130_fd_sc_hd__o211a_1
X_17507_ _18400_/CLK _17507_/D vssd1 vssd1 vccd1 vccd1 _17507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15699_ _17107_/CLK _15699_/D vssd1 vssd1 vccd1 vccd1 _15699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08240_ _15085_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08240_/X sky130_fd_sc_hd__or2_1
X_17438_ _17446_/CLK _17438_/D vssd1 vssd1 vccd1 vccd1 _17438_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_15 _13116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 _13180_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_37 _13260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08171_ _08171_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _15723_/D sky130_fd_sc_hd__and2_1
XANTENNA_48 _15525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17369_ _18013_/CLK _17369_/D vssd1 vssd1 vccd1 vccd1 _17369_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_59 hold484/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5005 _11479_/X vssd1 vssd1 vccd1 vccd1 _16983_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5016 _17090_/Q vssd1 vssd1 vccd1 vccd1 hold5016/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5027 _11053_/X vssd1 vssd1 vccd1 vccd1 _16841_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput100 _13105_/A vssd1 vssd1 vccd1 vccd1 hold5876/A sky130_fd_sc_hd__buf_6
Xhold5038 _16881_/Q vssd1 vssd1 vccd1 vccd1 hold5038/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5049 _10288_/X vssd1 vssd1 vccd1 vccd1 _16586_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput111 hold5972/X vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_12
Xhold4304 _13845_/Y vssd1 vssd1 vccd1 vccd1 _13846_/B sky130_fd_sc_hd__dlygate4sd3_1
Xoutput122 hold5968/X vssd1 vssd1 vccd1 vccd1 hold5969/A sky130_fd_sc_hd__buf_6
Xhold4315 _17103_/Q vssd1 vssd1 vccd1 vccd1 hold4315/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4326 _16732_/Q vssd1 vssd1 vccd1 vccd1 hold4326/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput133 hold5912/X vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_12
XFILLER_0_203_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4337 _16919_/Q vssd1 vssd1 vccd1 vccd1 hold4337/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput144 hold907/X vssd1 vssd1 vccd1 vccd1 load_status[4] sky130_fd_sc_hd__buf_12
Xhold3603 _09643_/X vssd1 vssd1 vccd1 vccd1 _16371_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4348 _11214_/Y vssd1 vssd1 vccd1 vccd1 _11215_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3614 _16442_/Q vssd1 vssd1 vccd1 vccd1 hold3614/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4359 hold5922/X vssd1 vssd1 vccd1 vccd1 hold5923/A sky130_fd_sc_hd__buf_4
Xhold3625 _12980_/X vssd1 vssd1 vccd1 vccd1 _12981_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3636 _17365_/Q vssd1 vssd1 vccd1 vccd1 hold3636/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3647 _13435_/X vssd1 vssd1 vccd1 vccd1 _17598_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2902 _15701_/Q vssd1 vssd1 vccd1 vccd1 hold2902/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2913 _07836_/X vssd1 vssd1 vccd1 vccd1 _15563_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3658 _16487_/Q vssd1 vssd1 vccd1 vccd1 hold3658/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3669 _10294_/X vssd1 vssd1 vccd1 vccd1 _16588_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2924 _16178_/Q vssd1 vssd1 vccd1 vccd1 hold2924/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_68_wb_clk_i clkbuf_6_19_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18460_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2935 _16236_/Q vssd1 vssd1 vccd1 vccd1 hold2935/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2946 _15756_/Q vssd1 vssd1 vccd1 vccd1 hold2946/X sky130_fd_sc_hd__dlygate4sd3_1
X_07955_ hold1170/X _07991_/A2 _07954_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _07955_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2957 _08298_/X vssd1 vssd1 vccd1 vccd1 _15782_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2968 _14047_/X vssd1 vssd1 vccd1 vccd1 _17829_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2979 _15831_/Q vssd1 vssd1 vccd1 vccd1 hold2979/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07886_ _14395_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07886_/X sky130_fd_sc_hd__or2_1
X_09625_ hold4691/X _10031_/B _09624_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09625_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09556_ hold3726/X _10052_/B _09555_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _09556_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08507_ _14166_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08507_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09487_ _13056_/C hold935/X _13034_/D hold907/X vssd1 vssd1 vccd1 vccd1 _13035_/D
+ sky130_fd_sc_hd__a31o_1
X_08438_ hold1436/X _08433_/B _08437_/X _13765_/C1 vssd1 vssd1 vccd1 vccd1 _08438_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_230_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08369_ _08373_/A _08369_/B vssd1 vssd1 vccd1 vccd1 _15816_/D sky130_fd_sc_hd__and2_1
XFILLER_0_18_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10400_ hold2583/X _16624_/Q _10538_/S vssd1 vssd1 vccd1 vccd1 _10401_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_116_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11380_ hold4883/X _11195_/B _11379_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _11380_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10331_ hold2033/X hold3272/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10332_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5550 _10816_/X vssd1 vssd1 vccd1 vccd1 _16762_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13050_ hold5938/X hold907/X _13055_/C vssd1 vssd1 vccd1 vccd1 _13225_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_225_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10262_ hold3106/X _16578_/Q _10628_/C vssd1 vssd1 vccd1 vccd1 _10263_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_30_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5561 _16957_/Q vssd1 vssd1 vccd1 vccd1 hold5561/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5572 _12094_/X vssd1 vssd1 vccd1 vccd1 _17188_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5583 _17069_/Q vssd1 vssd1 vccd1 vccd1 hold5583/X sky130_fd_sc_hd__dlygate4sd3_1
X_12001_ hold4970/X _12308_/B _12000_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _12001_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5594 _11449_/X vssd1 vssd1 vccd1 vccd1 _16973_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4860 _12202_/X vssd1 vssd1 vccd1 vccd1 _17224_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10193_ hold2721/X _16555_/Q _10385_/S vssd1 vssd1 vccd1 vccd1 _10194_/B sky130_fd_sc_hd__mux2_1
Xhold4871 _17266_/Q vssd1 vssd1 vccd1 vccd1 hold4871/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4882 _11119_/X vssd1 vssd1 vccd1 vccd1 _16863_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4893 _17232_/Q vssd1 vssd1 vccd1 vccd1 hold4893/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout360 _15549_/B vssd1 vssd1 vccd1 vccd1 _15559_/B sky130_fd_sc_hd__buf_4
Xfanout371 hold339/X vssd1 vssd1 vccd1 vccd1 hold340/A sky130_fd_sc_hd__buf_6
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout382 hold331/X vssd1 vssd1 vccd1 vccd1 _14880_/B sky130_fd_sc_hd__buf_6
X_16740_ _18039_/CLK _16740_/D vssd1 vssd1 vccd1 vccd1 _16740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout393 _14666_/B vssd1 vssd1 vccd1 vccd1 _14664_/B sky130_fd_sc_hd__buf_6
X_13952_ _15513_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13952_/X sky130_fd_sc_hd__or2_1
XFILLER_0_233_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12903_ _12906_/A _12903_/B vssd1 vssd1 vccd1 vccd1 _17477_/D sky130_fd_sc_hd__and2_1
X_16671_ _18229_/CLK _16671_/D vssd1 vssd1 vccd1 vccd1 _16671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13883_ _17748_/Q _13883_/B _13883_/C vssd1 vssd1 vccd1 vccd1 _13883_/X sky130_fd_sc_hd__and3_1
XFILLER_0_232_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18410_ _18410_/CLK _18410_/D vssd1 vssd1 vccd1 vccd1 _18410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15622_ _17154_/CLK _15622_/D vssd1 vssd1 vccd1 vccd1 _15622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12834_ _12837_/A _12834_/B vssd1 vssd1 vccd1 vccd1 _17454_/D sky130_fd_sc_hd__and2_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18341_ _18369_/CLK _18341_/D vssd1 vssd1 vccd1 vccd1 _18341_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _15553_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15553_/X sky130_fd_sc_hd__or2_1
X_12765_ _12786_/A _12765_/B vssd1 vssd1 vccd1 vccd1 _17431_/D sky130_fd_sc_hd__and2_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_445_wb_clk_i clkbuf_6_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17190_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ hold2133/X _14537_/B _14503_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _14504_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18272_ _18418_/CLK _18272_/D vssd1 vssd1 vccd1 vccd1 _18272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ hold5547/X _12305_/B _11715_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _11716_/X
+ sky130_fd_sc_hd__o211a_1
X_15484_ hold865/X _15484_/A2 _15484_/B1 hold745/X vssd1 vssd1 vccd1 vccd1 _15489_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12696_ _12843_/A _12696_/B vssd1 vssd1 vccd1 vccd1 _17408_/D sky130_fd_sc_hd__and2_1
XFILLER_0_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17223_ _18445_/CLK _17223_/D vssd1 vssd1 vccd1 vccd1 _17223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14435_ _15169_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14435_/X sky130_fd_sc_hd__or2_1
XFILLER_0_115_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11647_ hold5480/X _12323_/B _11646_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11647_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 input13/A vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_1
XFILLER_0_154_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput24 hold80/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__buf_6
X_17154_ _17154_/CLK _17154_/D vssd1 vssd1 vccd1 vccd1 _17154_/Q sky130_fd_sc_hd__dfxtp_1
Xinput35 input35/A vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14366_ _14368_/A _14366_/B vssd1 vssd1 vccd1 vccd1 _17982_/D sky130_fd_sc_hd__and2_1
XFILLER_0_135_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput46 input46/A vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__buf_6
X_11578_ hold5133/X _11789_/B _11577_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _11578_/X
+ sky130_fd_sc_hd__o211a_1
Xinput57 input57/A vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__buf_6
X_16105_ _17293_/CLK _16105_/D vssd1 vssd1 vccd1 vccd1 hold541/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput68 input68/A vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_1
Xhold808 hold808/A vssd1 vssd1 vccd1 vccd1 hold808/X sky130_fd_sc_hd__dlygate4sd3_1
X_13317_ _13797_/A _13317_/B vssd1 vssd1 vccd1 vccd1 _13317_/X sky130_fd_sc_hd__or2_1
X_10529_ hold1714/X hold3251/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10530_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold819 input52/X vssd1 vssd1 vccd1 vccd1 hold819/X sky130_fd_sc_hd__buf_1
X_17085_ _17901_/CLK _17085_/D vssd1 vssd1 vccd1 vccd1 _17085_/Q sky130_fd_sc_hd__dfxtp_1
X_14297_ hold1101/X _14333_/A2 _14296_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _14297_/X
+ sky130_fd_sc_hd__o211a_1
X_16036_ _17301_/CLK _16036_/D vssd1 vssd1 vccd1 vccd1 hold590/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13248_ _13241_/X _13247_/X _13296_/B1 vssd1 vssd1 vccd1 vccd1 _17549_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_204_1338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13179_ _13178_/X hold4751/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13179_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_209_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2209 _17808_/Q vssd1 vssd1 vccd1 vccd1 hold2209/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1508 _09407_/X vssd1 vssd1 vccd1 vccd1 _16289_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17987_ _18051_/CLK _17987_/D vssd1 vssd1 vccd1 vccd1 hold786/A sky130_fd_sc_hd__dfxtp_1
Xhold1519 _18131_/Q vssd1 vssd1 vccd1 vccd1 hold1519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16938_ _18432_/CLK _16938_/D vssd1 vssd1 vccd1 vccd1 _16938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16869_ _18072_/CLK _16869_/D vssd1 vssd1 vccd1 vccd1 _16869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09410_ _09438_/B _16291_/Q vssd1 vssd1 vccd1 vccd1 _09410_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09341_ _07809_/B _07802_/B _15481_/A1 vssd1 vssd1 vccd1 vccd1 _09342_/B sky130_fd_sc_hd__o21bai_4
Xclkbuf_leaf_186_wb_clk_i clkbuf_6_54_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18394_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09272_ _09272_/A hold272/X vssd1 vssd1 vccd1 vccd1 hold273/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_115_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16129_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08223_ _15557_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08223_/X sky130_fd_sc_hd__or2_1
XFILLER_0_56_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08154_ _15559_/A hold1241/X hold108/X vssd1 vssd1 vccd1 vccd1 _08155_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08085_ hold2293/X _08088_/B _08084_/Y _13925_/A vssd1 vssd1 vccd1 vccd1 _08085_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4101 _16988_/Q vssd1 vssd1 vccd1 vccd1 hold4101/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4112 _11230_/X vssd1 vssd1 vccd1 vccd1 _16900_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4123 _17618_/Q vssd1 vssd1 vccd1 vccd1 hold4123/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4134 _15273_/X vssd1 vssd1 vccd1 vccd1 _15274_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4145 _16398_/Q vssd1 vssd1 vccd1 vccd1 hold4145/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3400 _17418_/Q vssd1 vssd1 vccd1 vccd1 hold3400/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3411 _16331_/Q vssd1 vssd1 vccd1 vccd1 _13118_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4156 _16985_/Q vssd1 vssd1 vccd1 vccd1 hold4156/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3422 _10627_/Y vssd1 vssd1 vccd1 vccd1 _16699_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4167 _16816_/Q vssd1 vssd1 vccd1 vccd1 hold4167/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3433 _10059_/Y vssd1 vssd1 vccd1 vccd1 _10060_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4178 _11623_/X vssd1 vssd1 vccd1 vccd1 _17031_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4189 hold5934/X vssd1 vssd1 vccd1 vccd1 hold5935/A sky130_fd_sc_hd__buf_4
XTAP_5606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3444 _11143_/Y vssd1 vssd1 vccd1 vccd1 _16871_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2710 _15120_/X vssd1 vssd1 vccd1 vccd1 _18344_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3455 _12346_/Y vssd1 vssd1 vccd1 vccd1 _17272_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2721 _18113_/Q vssd1 vssd1 vccd1 vccd1 hold2721/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3466 _11775_/Y vssd1 vssd1 vccd1 vccd1 _11776_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2732 _14247_/X vssd1 vssd1 vccd1 vccd1 _17924_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08987_ hold315/X hold858/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08988_/B sky130_fd_sc_hd__mux2_1
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3477 _11220_/Y vssd1 vssd1 vccd1 vccd1 _11221_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3488 _16533_/Q vssd1 vssd1 vccd1 vccd1 hold3488/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2743 _18169_/Q vssd1 vssd1 vccd1 vccd1 hold2743/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3499 _16529_/Q vssd1 vssd1 vccd1 vccd1 hold3499/X sky130_fd_sc_hd__clkbuf_2
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2754 _16219_/Q vssd1 vssd1 vccd1 vccd1 hold2754/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2765 _18110_/Q vssd1 vssd1 vccd1 vccd1 hold2765/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07938_ _14735_/A hold355/X vssd1 vssd1 vccd1 vccd1 _07938_/Y sky130_fd_sc_hd__nor2_1
Xhold2776 _08040_/X vssd1 vssd1 vccd1 vccd1 _15661_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2787 _15697_/Q vssd1 vssd1 vccd1 vccd1 hold2787/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2798 _17797_/Q vssd1 vssd1 vccd1 vccd1 hold2798/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07869_ _15221_/A _07869_/B vssd1 vssd1 vccd1 vccd1 _07869_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_196_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09608_ _18273_/Q hold4677/X _09992_/C vssd1 vssd1 vccd1 vccd1 _09609_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10880_ hold786/X hold4138/X _11168_/C vssd1 vssd1 vccd1 vccd1 _10881_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_211_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_39_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_39_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09539_ _18250_/Q _16337_/Q _10004_/C vssd1 vssd1 vccd1 vccd1 _09540_/B sky130_fd_sc_hd__mux2_1
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12550_ hold1121/X _17361_/Q _12925_/S vssd1 vssd1 vccd1 vccd1 _12550_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11501_ hold2985/X _16991_/Q _12173_/S vssd1 vssd1 vccd1 vccd1 _11502_/B sky130_fd_sc_hd__mux2_1
X_12481_ hold50/X _12509_/A2 _12501_/A3 _12480_/X _12440_/A vssd1 vssd1 vccd1 vccd1
+ hold51/A sky130_fd_sc_hd__o311a_1
XFILLER_0_65_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14220_ _14970_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14220_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11432_ hold1859/X _16968_/Q _11717_/C vssd1 vssd1 vccd1 vccd1 _11433_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_149_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14151_ hold2056/X _14148_/B _14150_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _14151_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11363_ hold1289/X _16945_/Q _11654_/S vssd1 vssd1 vccd1 vccd1 _11364_/B sky130_fd_sc_hd__mux2_1
Xhold6070 data_in[31] vssd1 vssd1 vccd1 vccd1 hold275/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13102_ _13102_/A _13294_/B vssd1 vssd1 vccd1 vccd1 _13102_/X sky130_fd_sc_hd__or2_1
XFILLER_0_238_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10314_ _10542_/A _10314_/B vssd1 vssd1 vccd1 vccd1 _10314_/X sky130_fd_sc_hd__or2_1
Xhold6081 _18231_/Q vssd1 vssd1 vccd1 vccd1 hold6081/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6092 data_in[6] vssd1 vssd1 vccd1 vccd1 hold194/A sky130_fd_sc_hd__dlygate4sd3_1
X_14082_ _15535_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14082_/X sky130_fd_sc_hd__or2_1
XFILLER_0_225_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11294_ hold1505/X hold3465/X _12242_/S vssd1 vssd1 vccd1 vccd1 _11295_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_162_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_237_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5380 _17135_/Q vssd1 vssd1 vccd1 vccd1 hold5380/X sky130_fd_sc_hd__dlygate4sd3_1
X_13033_ _13056_/C hold896/X _13032_/Y vssd1 vssd1 vccd1 vccd1 hold897/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17910_ _17910_/CLK _17910_/D vssd1 vssd1 vccd1 vccd1 _17910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10245_ _10515_/A _10245_/B vssd1 vssd1 vccd1 vccd1 _10245_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5391 _11260_/X vssd1 vssd1 vccd1 vccd1 _16910_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4690 _13531_/X vssd1 vssd1 vccd1 vccd1 _17630_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_238_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10176_ _10482_/A _10176_/B vssd1 vssd1 vccd1 vccd1 _10176_/X sky130_fd_sc_hd__or2_1
X_17841_ _17873_/CLK _17841_/D vssd1 vssd1 vccd1 vccd1 _17841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_234_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14984_ _15199_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14984_/X sky130_fd_sc_hd__or2_1
X_17772_ _17838_/CLK hold555/X vssd1 vssd1 vccd1 vccd1 _17772_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout190 fanout210/X vssd1 vssd1 vccd1 vccd1 _12332_/B sky130_fd_sc_hd__clkbuf_4
X_16723_ _17967_/CLK _16723_/D vssd1 vssd1 vccd1 vccd1 _16723_/Q sky130_fd_sc_hd__dfxtp_1
X_13935_ _13935_/A _13935_/B vssd1 vssd1 vccd1 vccd1 _17775_/D sky130_fd_sc_hd__and2_1
XFILLER_0_233_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16654_ _18212_/CLK _16654_/D vssd1 vssd1 vccd1 vccd1 _16654_/Q sky130_fd_sc_hd__dfxtp_1
X_13866_ hold4442/X _13776_/A _13865_/X vssd1 vssd1 vccd1 vccd1 _13866_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15605_ _17590_/CLK _15605_/D vssd1 vssd1 vccd1 vccd1 _15605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12817_ hold2954/X hold3136/X _12844_/S vssd1 vssd1 vccd1 vccd1 _12817_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16585_ _18205_/CLK _16585_/D vssd1 vssd1 vccd1 vccd1 _16585_/Q sky130_fd_sc_hd__dfxtp_1
X_13797_ _13797_/A _13797_/B vssd1 vssd1 vccd1 vccd1 _13797_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18324_ _18324_/CLK _18324_/D vssd1 vssd1 vccd1 vccd1 _18324_/Q sky130_fd_sc_hd__dfxtp_1
X_15536_ hold2155/X _15547_/B _15535_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _15536_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _16247_/Q _17427_/Q _12811_/S vssd1 vssd1 vccd1 vccd1 _12748_/X sky130_fd_sc_hd__mux2_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18255_ _18327_/CLK _18255_/D vssd1 vssd1 vccd1 vccd1 _18255_/Q sky130_fd_sc_hd__dfxtp_1
X_15467_ _15988_/Q _09365_/B _15485_/B1 hold326/X vssd1 vssd1 vccd1 vccd1 _15467_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12679_ hold2756/X hold3376/X _12844_/S vssd1 vssd1 vccd1 vccd1 _12679_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17206_ _17898_/CLK _17206_/D vssd1 vssd1 vccd1 vccd1 _17206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14418_ hold1897/X _14446_/A2 _14417_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _14418_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18186_ _18218_/CLK _18186_/D vssd1 vssd1 vccd1 vccd1 _18186_/Q sky130_fd_sc_hd__dfxtp_1
X_15398_ hold861/X _09386_/A _15441_/A2 hold800/X vssd1 vssd1 vccd1 vccd1 _15398_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17137_ _17902_/CLK _17137_/D vssd1 vssd1 vccd1 vccd1 _17137_/Q sky130_fd_sc_hd__dfxtp_1
X_14349_ _14457_/A hold2292/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14350_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold605 hold605/A vssd1 vssd1 vccd1 vccd1 input10/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 hold616/A vssd1 vssd1 vccd1 vccd1 input16/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold627 hold627/A vssd1 vssd1 vccd1 vccd1 hold627/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 hold638/A vssd1 vssd1 vccd1 vccd1 hold638/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold649 hold649/A vssd1 vssd1 vccd1 vccd1 hold649/X sky130_fd_sc_hd__dlygate4sd3_1
X_17068_ _17884_/CLK _17068_/D vssd1 vssd1 vccd1 vccd1 _17068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16019_ _16120_/CLK _16019_/D vssd1 vssd1 vccd1 vccd1 hold803/A sky130_fd_sc_hd__dfxtp_1
X_08910_ hold5/X hold283/X _08910_/S vssd1 vssd1 vccd1 vccd1 hold284/A sky130_fd_sc_hd__mux2_1
XFILLER_0_228_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09890_ hold2569/X _16454_/Q _09992_/C vssd1 vssd1 vccd1 vccd1 _09891_/B sky130_fd_sc_hd__mux2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2006 _18454_/Q vssd1 vssd1 vccd1 vccd1 hold2006/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_237_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08841_ _12412_/A _08841_/B vssd1 vssd1 vccd1 vccd1 _16039_/D sky130_fd_sc_hd__and2_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2017 _15737_/Q vssd1 vssd1 vccd1 vccd1 hold2017/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2028 _14817_/X vssd1 vssd1 vccd1 vccd1 _18198_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2039 _17781_/Q vssd1 vssd1 vccd1 vccd1 hold2039/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1305 _15692_/Q vssd1 vssd1 vccd1 vccd1 hold1305/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1316 _14937_/X vssd1 vssd1 vccd1 vccd1 _18255_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1327 _15771_/Q vssd1 vssd1 vccd1 vccd1 hold1327/X sky130_fd_sc_hd__dlygate4sd3_1
X_08772_ _15374_/A hold123/X vssd1 vssd1 vccd1 vccd1 _16006_/D sky130_fd_sc_hd__and2_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1338 _16185_/Q vssd1 vssd1 vccd1 vccd1 hold1338/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1349 _14484_/X vssd1 vssd1 vccd1 vccd1 _18039_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_367_wb_clk_i clkbuf_6_34_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17702_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09324_ hold2495/X _09323_/B _09323_/Y _12597_/A vssd1 vssd1 vccd1 vccd1 _09324_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09255_ _15531_/A hold1069/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09256_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08206_ hold1680/X _08209_/B _08205_/X _13675_/C1 vssd1 vssd1 vccd1 vccd1 _08206_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09186_ _15515_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09186_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08137_ _08137_/A hold536/X vssd1 vssd1 vccd1 vccd1 _15707_/D sky130_fd_sc_hd__and2_1
XFILLER_0_146_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_83_wb_clk_i clkbuf_6_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17492_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08068_ _14413_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08068_/X sky130_fd_sc_hd__or2_1
XFILLER_0_222_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_12_wb_clk_i clkbuf_6_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18448_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3230 _17446_/Q vssd1 vssd1 vccd1 vccd1 hold3230/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3241 _10195_/X vssd1 vssd1 vccd1 vccd1 _16555_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10030_ _11203_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _10030_/Y sky130_fd_sc_hd__nor2_1
XTAP_5414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3252 _10435_/X vssd1 vssd1 vccd1 vccd1 _16635_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3263 _17379_/Q vssd1 vssd1 vccd1 vccd1 hold3263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3274 _16553_/Q vssd1 vssd1 vccd1 vccd1 hold3274/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3285 _10291_/X vssd1 vssd1 vccd1 vccd1 _16587_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2540 _07852_/X vssd1 vssd1 vccd1 vccd1 _15571_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3296 _16665_/Q vssd1 vssd1 vccd1 vccd1 hold3296/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2551 _15166_/X vssd1 vssd1 vccd1 vccd1 _18366_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2562 _16193_/Q vssd1 vssd1 vccd1 vccd1 hold2562/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2573 _18041_/Q vssd1 vssd1 vccd1 vccd1 hold2573/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2584 _14783_/X vssd1 vssd1 vccd1 vccd1 _18182_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2595 _14611_/X vssd1 vssd1 vccd1 vccd1 _18099_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1850 _14115_/X vssd1 vssd1 vccd1 vccd1 _17861_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1861 _18286_/Q vssd1 vssd1 vccd1 vccd1 hold1861/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1872 _14715_/X vssd1 vssd1 vccd1 vccd1 _18149_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ hold1600/X _17151_/Q _12173_/S vssd1 vssd1 vccd1 vccd1 _11982_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_215_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1883 _15717_/Q vssd1 vssd1 vccd1 vccd1 hold1883/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1894 _14552_/X vssd1 vssd1 vccd1 vccd1 _18072_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13720_ hold5809/X _13808_/B _13719_/X _12753_/A vssd1 vssd1 vccd1 vccd1 _13720_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10932_ _11670_/A _10932_/B vssd1 vssd1 vccd1 vccd1 _10932_/X sky130_fd_sc_hd__or2_1
XFILLER_0_211_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13651_ hold5579/X _13847_/B _13650_/X _13765_/C1 vssd1 vssd1 vccd1 vccd1 _13651_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_1386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10863_ _11043_/A _10863_/B vssd1 vssd1 vccd1 vccd1 _10863_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12602_ hold3286/X _12601_/X _12923_/S vssd1 vssd1 vccd1 vccd1 _12602_/X sky130_fd_sc_hd__mux2_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _18315_/CLK _16370_/D vssd1 vssd1 vccd1 vccd1 _16370_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ hold3989/X _13868_/B _13581_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _13582_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10794_ _11010_/A _10794_/B vssd1 vssd1 vccd1 vccd1 _10794_/X sky130_fd_sc_hd__or2_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15321_ _16296_/Q _15477_/A2 _15487_/B1 hold649/X _15320_/X vssd1 vssd1 vccd1 vccd1
+ _15322_/D sky130_fd_sc_hd__a221o_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12533_ hold4519/X _12532_/X _12929_/S vssd1 vssd1 vccd1 vccd1 _12533_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18040_ _18072_/CLK _18040_/D vssd1 vssd1 vccd1 vccd1 _18040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15252_ _15489_/A _15252_/B _15252_/C _15252_/D vssd1 vssd1 vccd1 vccd1 _15252_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_136_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12464_ _17325_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12464_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14203_ hold2603/X _14202_/B _14202_/Y _08125_/A vssd1 vssd1 vccd1 vccd1 _14203_/X
+ sky130_fd_sc_hd__o211a_1
X_11415_ _12174_/A _11415_/B vssd1 vssd1 vccd1 vccd1 _11415_/X sky130_fd_sc_hd__or2_1
X_15183_ _15183_/A _15227_/B vssd1 vssd1 vccd1 vccd1 _15183_/X sky130_fd_sc_hd__or2_1
X_12395_ hold679/X hold888/X _12441_/S vssd1 vssd1 vccd1 vccd1 hold889/A sky130_fd_sc_hd__mux2_1
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14134_ _15207_/A _14140_/B vssd1 vssd1 vccd1 vccd1 _14134_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11346_ _11631_/A _11346_/B vssd1 vssd1 vccd1 vccd1 _11346_/X sky130_fd_sc_hd__or2_1
XFILLER_0_61_1419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_240_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14065_ hold2577/X _14107_/A2 _14064_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _14065_/X
+ sky130_fd_sc_hd__o211a_1
X_11277_ _12243_/A _11277_/B vssd1 vssd1 vccd1 vccd1 _11277_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13016_ hold1062/X _13003_/Y _13015_/X _12984_/A vssd1 vssd1 vccd1 vccd1 _13016_/X
+ sky130_fd_sc_hd__o211a_1
X_10228_ hold4555/X _10604_/B _10227_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10228_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17824_ _17888_/CLK _17824_/D vssd1 vssd1 vccd1 vccd1 _17824_/Q sky130_fd_sc_hd__dfxtp_1
X_10159_ hold3322/X _10619_/B _10158_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10159_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__buf_1
XTAP_5970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14967_ hold445/X _15182_/B vssd1 vssd1 vccd1 vccd1 hold510/A sky130_fd_sc_hd__or2_4
X_17755_ _17949_/CLK _17755_/D vssd1 vssd1 vccd1 vccd1 _17755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_460_wb_clk_i clkbuf_6_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17754_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16706_ _18200_/CLK _16706_/D vssd1 vssd1 vccd1 vccd1 _16706_/Q sky130_fd_sc_hd__dfxtp_1
X_13918_ _15207_/A _17767_/Q hold297/X vssd1 vssd1 vccd1 vccd1 _13918_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_221_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14898_ hold927/X _14910_/B vssd1 vssd1 vccd1 vccd1 _14898_/X sky130_fd_sc_hd__or2_1
X_17686_ _17686_/CLK _17686_/D vssd1 vssd1 vccd1 vccd1 _17686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16637_ _18227_/CLK _16637_/D vssd1 vssd1 vccd1 vccd1 _16637_/Q sky130_fd_sc_hd__dfxtp_1
X_13849_ _13873_/A _13849_/B vssd1 vssd1 vccd1 vccd1 _13849_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_231_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16568_ _18126_/CLK _16568_/D vssd1 vssd1 vccd1 vccd1 _16568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18307_ _18307_/CLK _18307_/D vssd1 vssd1 vccd1 vccd1 _18307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15519_ _15519_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15519_/X sky130_fd_sc_hd__or2_1
X_16499_ _18380_/CLK _16499_/D vssd1 vssd1 vccd1 vccd1 _16499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09040_ hold5/X hold156/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09041_/B sky130_fd_sc_hd__mux2_1
X_18238_ _18242_/CLK _18238_/D vssd1 vssd1 vccd1 vccd1 _18238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18169_ _18224_/CLK _18169_/D vssd1 vssd1 vccd1 vccd1 _18169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold402 la_data_in[27] vssd1 vssd1 vccd1 vccd1 hold402/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold413 hold413/A vssd1 vssd1 vccd1 vccd1 hold413/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold424 hold424/A vssd1 vssd1 vccd1 vccd1 hold424/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 hold435/A vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold446 hold446/A vssd1 vssd1 vccd1 vccd1 hold446/X sky130_fd_sc_hd__clkbuf_2
Xhold457 hold457/A vssd1 vssd1 vccd1 vccd1 hold457/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold468 hold468/A vssd1 vssd1 vccd1 vccd1 hold468/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09942_ _09954_/A _09942_/B vssd1 vssd1 vccd1 vccd1 _09942_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold479 hold479/A vssd1 vssd1 vccd1 vccd1 hold479/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout904 hold579/X vssd1 vssd1 vccd1 vccd1 _15559_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout915 _15173_/A vssd1 vssd1 vccd1 vccd1 _15227_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout926 hold1022/X vssd1 vssd1 vccd1 vccd1 _15185_/A sky130_fd_sc_hd__buf_4
XFILLER_0_96_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09873_ _09978_/A _09873_/B vssd1 vssd1 vccd1 vccd1 _09873_/X sky130_fd_sc_hd__or2_1
Xfanout937 _15207_/A vssd1 vssd1 vccd1 vccd1 _15099_/A sky130_fd_sc_hd__buf_12
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout948 hold1193/X vssd1 vssd1 vccd1 vccd1 _15183_/A sky130_fd_sc_hd__clkbuf_4
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08824_ hold23/X hold527/X _08866_/S vssd1 vssd1 vccd1 vccd1 _08825_/B sky130_fd_sc_hd__mux2_1
Xhold1102 _14297_/X vssd1 vssd1 vccd1 vccd1 _17948_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 _18166_/Q vssd1 vssd1 vccd1 vccd1 hold1113/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1124 _08186_/X vssd1 vssd1 vccd1 vccd1 _15729_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 _08386_/X vssd1 vssd1 vccd1 vccd1 _08387_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 hold1146/A vssd1 vssd1 vccd1 vccd1 input40/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ hold77/X hold766/X _08779_/S vssd1 vssd1 vccd1 vccd1 _08756_/B sky130_fd_sc_hd__mux2_1
Xhold1157 _18282_/Q vssd1 vssd1 vccd1 vccd1 hold1157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1168 _14013_/X vssd1 vssd1 vccd1 vccd1 _17812_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 _18316_/Q vssd1 vssd1 vccd1 vccd1 hold1179/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _12418_/A _08686_/B vssd1 vssd1 vccd1 vccd1 _15964_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_130_wb_clk_i clkbuf_6_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17319_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_240_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09307_ _14988_/A _09315_/B vssd1 vssd1 vccd1 vccd1 _09307_/X sky130_fd_sc_hd__or2_1
XFILLER_0_118_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09238_ _12786_/A _09238_/B vssd1 vssd1 vccd1 vccd1 _16230_/D sky130_fd_sc_hd__and2_1
XFILLER_0_185_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09169_ hold1690/X _09177_/A2 _09168_/X _12906_/A vssd1 vssd1 vccd1 vccd1 _09169_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11200_ _12331_/A _11200_/B vssd1 vssd1 vccd1 vccd1 _11200_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_32_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12180_ _13749_/A _12180_/B vssd1 vssd1 vccd1 vccd1 _12180_/X sky130_fd_sc_hd__or2_1
X_11131_ hold4766/X _11765_/B _11130_/X _14346_/A vssd1 vssd1 vccd1 vccd1 _11131_/X
+ sky130_fd_sc_hd__o211a_1
Xhold980 hold980/A vssd1 vssd1 vccd1 vccd1 hold980/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold991 hold991/A vssd1 vssd1 vccd1 vccd1 hold991/X sky130_fd_sc_hd__buf_6
XTAP_5200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11062_ hold3991/X _10013_/B _11061_/X _14552_/C1 vssd1 vssd1 vccd1 vccd1 _11062_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_289_wb_clk_i clkbuf_6_37_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18020_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold3060 _13965_/X vssd1 vssd1 vccd1 vccd1 _17789_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10013_ _16495_/Q _10013_/B _10964_/S vssd1 vssd1 vccd1 vccd1 _10013_/X sky130_fd_sc_hd__and3_1
XFILLER_0_194_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3071 _09085_/X vssd1 vssd1 vccd1 vccd1 _16157_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3082 _18141_/Q vssd1 vssd1 vccd1 vccd1 hold3082/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15870_ _17244_/CLK _15870_/D vssd1 vssd1 vccd1 vccd1 _15870_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_218_wb_clk_i clkbuf_6_61_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18211_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3093 _18056_/Q vssd1 vssd1 vccd1 vccd1 hold3093/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2370 _14923_/X vssd1 vssd1 vccd1 vccd1 _18248_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2381 _14613_/X vssd1 vssd1 vccd1 vccd1 _18100_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14821_ hold2058/X _14828_/B _14820_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _14821_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2392 _18000_/Q vssd1 vssd1 vccd1 vccd1 hold2392/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1680 _15739_/Q vssd1 vssd1 vccd1 vccd1 hold1680/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17540_ _18380_/CLK _17540_/D vssd1 vssd1 vccd1 vccd1 _17540_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ _15145_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14752_/X sky130_fd_sc_hd__or2_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1691 _09169_/X vssd1 vssd1 vccd1 vccd1 _16197_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _12255_/A _11964_/B vssd1 vssd1 vccd1 vccd1 _11964_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ hold2420/X hold3952/X _13817_/C vssd1 vssd1 vccd1 vccd1 _13704_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_196_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10915_ hold5201/X _11171_/B _10914_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _10915_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17471_ _17471_/CLK _17471_/D vssd1 vssd1 vccd1 vccd1 _17471_/Q sky130_fd_sc_hd__dfxtp_1
X_14683_ hold2113/X _14718_/B _14682_/X _14853_/C1 vssd1 vssd1 vccd1 vccd1 _14683_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11895_ _13749_/A _11895_/B vssd1 vssd1 vccd1 vccd1 _11895_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16422_ _18377_/CLK _16422_/D vssd1 vssd1 vccd1 vccd1 _16422_/Q sky130_fd_sc_hd__dfxtp_1
X_13634_ hold2499/X hold4731/X _13862_/C vssd1 vssd1 vccd1 vccd1 _13635_/B sky130_fd_sc_hd__mux2_1
X_10846_ hold5364/X _11744_/B _10845_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _10846_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16353_ _18298_/CLK _16353_/D vssd1 vssd1 vccd1 vccd1 _16353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13565_ hold940/X _17642_/Q _13874_/C vssd1 vssd1 vccd1 vccd1 _13566_/B sky130_fd_sc_hd__mux2_1
X_10777_ hold4837/X _11162_/B _10776_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _10777_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15304_ _15344_/A _15304_/B vssd1 vssd1 vccd1 vccd1 _18406_/D sky130_fd_sc_hd__and2_1
X_12516_ _15284_/A _12516_/B vssd1 vssd1 vccd1 vccd1 _17348_/D sky130_fd_sc_hd__and2_1
XFILLER_0_70_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16284_ _18411_/CLK _16284_/D vssd1 vssd1 vccd1 vccd1 _16284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13496_ hold1632/X hold5418/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13497_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15235_ hold870/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15235_/X sky130_fd_sc_hd__or2_1
X_18023_ _18023_/CLK _18023_/D vssd1 vssd1 vccd1 vccd1 _18023_/Q sky130_fd_sc_hd__dfxtp_1
X_12447_ hold226/X _12445_/A _12445_/B _12446_/X _15374_/A vssd1 vssd1 vccd1 vccd1
+ hold27/A sky130_fd_sc_hd__o311a_1
XFILLER_0_48_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15166_ hold2550/X _15165_/B _15165_/Y _15042_/A vssd1 vssd1 vccd1 vccd1 _15166_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12378_ hold4320/X _13407_/A _12377_/X vssd1 vssd1 vccd1 vccd1 _12378_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_205_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_1318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14117_ hold3049/X _14142_/B _14116_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14117_/X
+ sky130_fd_sc_hd__o211a_1
X_11329_ hold5591/X _12305_/B _11328_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _11329_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_239_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15097_ _15205_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15097_/X sky130_fd_sc_hd__or2_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_238_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14048_ _15229_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14048_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17807_ _17871_/CLK _17807_/D vssd1 vssd1 vccd1 vccd1 _17807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15999_ _16082_/CLK _15999_/D vssd1 vssd1 vccd1 vccd1 hold412/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08540_ hold71/X hold324/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08541_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_206_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17738_ _17738_/CLK _17738_/D vssd1 vssd1 vccd1 vccd1 _17738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08471_ hold1430/X _08486_/B _08470_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _08471_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17669_ _17733_/CLK _17669_/D vssd1 vssd1 vccd1 vccd1 _17669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09023_ _12426_/A hold434/X vssd1 vssd1 vccd1 vccd1 _16128_/D sky130_fd_sc_hd__and2_1
XFILLER_0_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5902 output72/X vssd1 vssd1 vccd1 vccd1 data_out[0] sky130_fd_sc_hd__buf_12
Xhold5913 _18415_/Q vssd1 vssd1 vccd1 vccd1 hold5913/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5924 _18406_/Q vssd1 vssd1 vccd1 vccd1 hold5924/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold210 input6/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5935 hold5935/A vssd1 vssd1 vccd1 vccd1 hold5935/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_206_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold221 hold221/A vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5946 hold5946/A vssd1 vssd1 vccd1 vccd1 hold5946/X sky130_fd_sc_hd__clkbuf_4
Xhold232 la_data_in[19] vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5957 hold5957/A vssd1 vssd1 vccd1 vccd1 hold5957/X sky130_fd_sc_hd__clkbuf_4
Xhold243 hold61/X vssd1 vssd1 vccd1 vccd1 input14/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5968 hold6099/X vssd1 vssd1 vccd1 vccd1 hold5968/X sky130_fd_sc_hd__clkbuf_4
Xhold254 hold50/X vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_229_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5979 _07797_/X vssd1 vssd1 vccd1 vccd1 _18459_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 hold265/A vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold276 hold67/X vssd1 vssd1 vccd1 vccd1 input29/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 hold287/A vssd1 vssd1 vccd1 vccd1 input53/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout701 fanout739/X vssd1 vssd1 vccd1 vccd1 _08851_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout712 _15491_/A vssd1 vssd1 vccd1 vccd1 _15364_/A sky130_fd_sc_hd__clkbuf_4
X_09925_ _10019_/A _10046_/B _09924_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09925_/X
+ sky130_fd_sc_hd__o211a_1
Xhold298 hold298/A vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout723 _15404_/A vssd1 vssd1 vccd1 vccd1 _15234_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_141_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_382_wb_clk_i clkbuf_6_33_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17266_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout734 _08954_/A vssd1 vssd1 vccd1 vccd1 _15042_/A sky130_fd_sc_hd__buf_4
Xfanout745 _08111_/A vssd1 vssd1 vccd1 vccd1 _08143_/A sky130_fd_sc_hd__buf_4
Xfanout756 _14380_/A vssd1 vssd1 vccd1 vccd1 _13903_/A sky130_fd_sc_hd__buf_4
X_09856_ hold3543/X _10046_/B _09855_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09856_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout767 fanout791/X vssd1 vssd1 vccd1 vccd1 _08347_/A sky130_fd_sc_hd__buf_4
XFILLER_0_176_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout778 _13917_/A vssd1 vssd1 vccd1 vccd1 _13925_/A sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_311_wb_clk_i clkbuf_6_45_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18005_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout789 fanout791/X vssd1 vssd1 vccd1 vccd1 _14346_/A sky130_fd_sc_hd__buf_4
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08807_ _12410_/A hold795/X vssd1 vssd1 vccd1 vccd1 _16022_/D sky130_fd_sc_hd__and2_1
XFILLER_0_77_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ hold3736/X _10049_/B _09786_/X _15212_/C1 vssd1 vssd1 vccd1 vccd1 _09787_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _12426_/A hold824/X vssd1 vssd1 vccd1 vccd1 _15989_/D sky130_fd_sc_hd__and2_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 _15056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_116 hold915/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _15173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ hold131/X hold189/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold190/A sky130_fd_sc_hd__mux2_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10700_ hold2952/X hold4350/X _11660_/S vssd1 vssd1 vccd1 vccd1 _10701_/B sky130_fd_sc_hd__mux2_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ hold5291/X _11771_/B _11679_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _11680_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10631_ _16701_/Q _10631_/B _10637_/C vssd1 vssd1 vccd1 vccd1 _10631_/X sky130_fd_sc_hd__and3_1
XFILLER_0_181_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13350_ _13734_/A _13350_/B vssd1 vssd1 vccd1 vccd1 _13350_/X sky130_fd_sc_hd__or2_1
X_10562_ hold1283/X hold3848/X _10634_/C vssd1 vssd1 vccd1 vccd1 _10563_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12301_ _12301_/A _12301_/B vssd1 vssd1 vccd1 vccd1 _17257_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_133_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13281_ _13281_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13281_/X sky130_fd_sc_hd__and2_1
XFILLER_0_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10493_ hold2051/X hold3337/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10494_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_228_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15020_ hold113/X _15182_/B vssd1 vssd1 vccd1 vccd1 _15020_/X sky130_fd_sc_hd__or2_4
XFILLER_0_32_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12232_ hold4871/X _12356_/B _12231_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _12232_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12163_ hold4885/X _12353_/B _12162_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _12163_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11114_ hold2314/X _16862_/Q _11753_/C vssd1 vssd1 vccd1 vccd1 _11115_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_236_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12094_ hold5571/X _12305_/B _12093_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _12094_/X
+ sky130_fd_sc_hd__o211a_1
X_16971_ _17883_/CLK _16971_/D vssd1 vssd1 vccd1 vccd1 _16971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15922_ _18417_/CLK _15922_/D vssd1 vssd1 vccd1 vccd1 hold722/A sky130_fd_sc_hd__dfxtp_1
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11045_ hold1867/X hold3836/X _11144_/C vssd1 vssd1 vccd1 vccd1 _11046_/B sky130_fd_sc_hd__mux2_1
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15853_ _17742_/CLK _15853_/D vssd1 vssd1 vccd1 vccd1 _15853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14804_ _15197_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14804_/X sky130_fd_sc_hd__or2_1
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ _15244_/A _12996_/B vssd1 vssd1 vccd1 vccd1 _17508_/D sky130_fd_sc_hd__and2_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15784_ _17716_/CLK _15784_/D vssd1 vssd1 vccd1 vccd1 _15784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17523_ _17523_/CLK hold906/X vssd1 vssd1 vccd1 vccd1 _17523_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14735_ _14735_/A _15182_/B vssd1 vssd1 vccd1 vccd1 _14780_/B sky130_fd_sc_hd__or2_4
XFILLER_0_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11947_ hold5695/X _12329_/B _11946_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _11947_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _15221_/A _14666_/B vssd1 vssd1 vccd1 vccd1 _14666_/Y sky130_fd_sc_hd__nand2_1
X_17454_ _17456_/CLK _17454_/D vssd1 vssd1 vccd1 vccd1 _17454_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11878_ hold5117/X _12356_/B _11877_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _11878_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16405_ _18324_/CLK _16405_/D vssd1 vssd1 vccd1 vccd1 _16405_/Q sky130_fd_sc_hd__dfxtp_1
X_13617_ _13722_/A _13617_/B vssd1 vssd1 vccd1 vccd1 _13617_/X sky130_fd_sc_hd__or2_1
XFILLER_0_95_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10829_ hold2008/X hold5372/X _11213_/C vssd1 vssd1 vccd1 vccd1 _10830_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_172_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14597_ hold1271/X _14612_/B _14596_/X _14895_/C1 vssd1 vssd1 vccd1 vccd1 _14597_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17385_ _18438_/CLK _17385_/D vssd1 vssd1 vccd1 vccd1 _17385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16336_ _18379_/CLK _16336_/D vssd1 vssd1 vccd1 vccd1 _16336_/Q sky130_fd_sc_hd__dfxtp_1
X_13548_ _13773_/A _13548_/B vssd1 vssd1 vccd1 vccd1 _13548_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16267_ _17978_/CLK _16267_/D vssd1 vssd1 vccd1 vccd1 _16267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13479_ _13737_/A _13479_/B vssd1 vssd1 vccd1 vccd1 _13479_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5209 _16857_/Q vssd1 vssd1 vccd1 vccd1 hold5209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15218_ hold1177/X _15221_/B _15217_/Y _15218_/C1 vssd1 vssd1 vccd1 vccd1 _15218_/X
+ sky130_fd_sc_hd__o211a_1
X_18006_ _18061_/CLK _18006_/D vssd1 vssd1 vccd1 vccd1 _18006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16198_ _17481_/CLK _16198_/D vssd1 vssd1 vccd1 vccd1 _16198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4508 _11803_/Y vssd1 vssd1 vccd1 vccd1 _17091_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4519 _17354_/Q vssd1 vssd1 vccd1 vccd1 hold4519/X sky130_fd_sc_hd__dlygate4sd3_1
X_15149_ _15203_/A _15157_/B vssd1 vssd1 vccd1 vccd1 _15149_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3807 _17417_/Q vssd1 vssd1 vccd1 vccd1 hold3807/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3818 _17168_/Q vssd1 vssd1 vccd1 vccd1 hold3818/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3829 _10666_/X vssd1 vssd1 vccd1 vccd1 _16712_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07971_ hold1752/X _07978_/B _07970_/X _08363_/A vssd1 vssd1 vccd1 vccd1 _07971_/X
+ sky130_fd_sc_hd__o211a_1
X_09710_ hold1423/X hold4604/X _11162_/C vssd1 vssd1 vccd1 vccd1 _09711_/B sky130_fd_sc_hd__mux2_1
X_09641_ hold1827/X hold3560/X _10025_/C vssd1 vssd1 vccd1 vccd1 _09642_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_93_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09572_ hold996/X _13254_/A _10040_/C vssd1 vssd1 vccd1 vccd1 _09573_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08523_ _08730_/A _13046_/C vssd1 vssd1 vccd1 vccd1 _08528_/S sky130_fd_sc_hd__or2_2
XFILLER_0_89_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08454_ _15513_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08454_/X sky130_fd_sc_hd__or2_1
XFILLER_0_77_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08385_ _08385_/A _08385_/B vssd1 vssd1 vccd1 vccd1 _15824_/D sky130_fd_sc_hd__and2_1
XFILLER_0_11_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09006_ hold684/X hold835/X _09056_/S vssd1 vssd1 vccd1 vccd1 hold836/A sky130_fd_sc_hd__mux2_1
Xhold5710 _12361_/Y vssd1 vssd1 vccd1 vccd1 _17277_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5721 _13806_/Y vssd1 vssd1 vccd1 vccd1 _13807_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5732 _11944_/X vssd1 vssd1 vccd1 vccd1 _17138_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5743 _17204_/Q vssd1 vssd1 vccd1 vccd1 hold5743/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5754 _10023_/Y vssd1 vssd1 vccd1 vccd1 _10024_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5765 _17177_/Q vssd1 vssd1 vccd1 vccd1 hold5765/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5776 _12064_/X vssd1 vssd1 vccd1 vccd1 _17178_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5787 _17657_/Q vssd1 vssd1 vccd1 vccd1 hold5787/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5798 _13612_/X vssd1 vssd1 vccd1 vccd1 _17657_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout520 _10619_/C vssd1 vssd1 vccd1 vccd1 _10637_/C sky130_fd_sc_hd__clkbuf_8
Xfanout531 _09178_/Y vssd1 vssd1 vccd1 vccd1 _09218_/B sky130_fd_sc_hd__buf_4
XFILLER_0_217_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout542 _08498_/B vssd1 vssd1 vccd1 vccd1 _08500_/B sky130_fd_sc_hd__clkbuf_8
X_09908_ hold1475/X _16460_/Q _10028_/C vssd1 vssd1 vccd1 vccd1 _09909_/B sky130_fd_sc_hd__mux2_1
Xfanout553 _08260_/B vssd1 vssd1 vccd1 vccd1 _08280_/B sky130_fd_sc_hd__buf_8
Xfanout564 _08043_/B vssd1 vssd1 vccd1 vccd1 _08045_/B sky130_fd_sc_hd__buf_8
Xfanout575 _07829_/Y vssd1 vssd1 vccd1 vccd1 _07869_/B sky130_fd_sc_hd__clkbuf_8
Xfanout586 _13310_/B vssd1 vssd1 vccd1 vccd1 _13294_/B sky130_fd_sc_hd__buf_8
X_09839_ hold2037/X _16437_/Q _10031_/C vssd1 vssd1 vccd1 vccd1 _09840_/B sky130_fd_sc_hd__mux2_1
Xfanout597 _12871_/S vssd1 vssd1 vccd1 vccd1 _12922_/S sky130_fd_sc_hd__buf_6
XFILLER_0_225_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12850_ hold1246/X _17461_/Q _12850_/S vssd1 vssd1 vccd1 vccd1 _12850_/X sky130_fd_sc_hd__mux2_1
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11801_ _17091_/Q _12335_/B _12335_/C vssd1 vssd1 vccd1 vccd1 _11801_/X sky130_fd_sc_hd__and3_1
XFILLER_0_186_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12781_ hold2289/X hold3619/X _12838_/S vssd1 vssd1 vccd1 vccd1 _12781_/X sky130_fd_sc_hd__mux2_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ hold3093/X _14541_/B _14519_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _14520_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _17068_/Q _11732_/B _11732_/C vssd1 vssd1 vccd1 vccd1 _11732_/X sky130_fd_sc_hd__and3_1
XFILLER_0_166_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14451_ hold915/X _14499_/B vssd1 vssd1 vccd1 vccd1 _14451_/X sky130_fd_sc_hd__or2_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11663_ hold2248/X hold5239/X _11765_/C vssd1 vssd1 vccd1 vccd1 _11664_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_166_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ hold5418/X _13883_/B _13401_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13402_/X
+ sky130_fd_sc_hd__o211a_1
X_10614_ hold3206/X _10542_/A _10613_/X vssd1 vssd1 vccd1 vccd1 _10614_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17170_ _17202_/CLK _17170_/D vssd1 vssd1 vccd1 vccd1 _17170_/Q sky130_fd_sc_hd__dfxtp_1
X_14382_ _15060_/A _14382_/B vssd1 vssd1 vccd1 vccd1 _17990_/D sky130_fd_sc_hd__and2_1
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11594_ _17870_/Q _17022_/Q _12329_/C vssd1 vssd1 vccd1 vccd1 _11595_/B sky130_fd_sc_hd__mux2_1
X_16121_ _17336_/CLK _16121_/D vssd1 vssd1 vccd1 vccd1 hold280/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13333_ hold4697/X _13811_/B _13332_/X _08363_/A vssd1 vssd1 vccd1 vccd1 _13333_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10545_ _10551_/A _10545_/B vssd1 vssd1 vccd1 vccd1 _10545_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16052_ _17338_/CLK _16052_/D vssd1 vssd1 vccd1 vccd1 hold697/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13264_ _13257_/X _13263_/X _13296_/B1 vssd1 vssd1 vccd1 vccd1 _17551_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_122_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10476_ _10476_/A _10476_/B vssd1 vssd1 vccd1 vccd1 _10476_/X sky130_fd_sc_hd__or2_1
X_15003_ hold2009/X hold447/X _15002_/Y _15068_/A vssd1 vssd1 vccd1 vccd1 _15003_/X
+ sky130_fd_sc_hd__o211a_1
X_12215_ hold1887/X _17229_/Q _12227_/S vssd1 vssd1 vccd1 vccd1 _12216_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13195_ _13194_/X _16917_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13195_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_233_wb_clk_i clkbuf_6_62_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18224_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12146_ hold2697/X hold5050/X _12242_/S vssd1 vssd1 vccd1 vccd1 _12147_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_102_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12077_ hold2910/X _17183_/Q _12173_/S vssd1 vssd1 vccd1 vccd1 _12078_/B sky130_fd_sc_hd__mux2_1
X_16954_ _17834_/CLK _16954_/D vssd1 vssd1 vccd1 vccd1 _16954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15905_ _17321_/CLK _15905_/D vssd1 vssd1 vccd1 vccd1 hold542/A sky130_fd_sc_hd__dfxtp_1
X_11028_ _11124_/A _11028_/B vssd1 vssd1 vccd1 vccd1 _11028_/X sky130_fd_sc_hd__or2_1
XFILLER_0_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16885_ _18056_/CLK _16885_/D vssd1 vssd1 vccd1 vccd1 _16885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15836_ _17709_/CLK _15836_/D vssd1 vssd1 vccd1 vccd1 _15836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12979_ hold2447/X _17504_/Q _12985_/S vssd1 vssd1 vccd1 vccd1 _12979_/X sky130_fd_sc_hd__mux2_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15767_ _17686_/CLK _15767_/D vssd1 vssd1 vccd1 vccd1 _15767_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17506_ _17506_/CLK _17506_/D vssd1 vssd1 vccd1 vccd1 _17506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14718_ _15165_/A _14718_/B vssd1 vssd1 vccd1 vccd1 _14718_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_86_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15698_ _17209_/CLK _15698_/D vssd1 vssd1 vccd1 vccd1 hold941/A sky130_fd_sc_hd__dfxtp_1
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17437_ _17437_/CLK _17437_/D vssd1 vssd1 vccd1 vccd1 _17437_/Q sky130_fd_sc_hd__dfxtp_1
X_14649_ hold2681/X _14664_/B _14648_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14649_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_16 _13132_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_27 _13180_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 _13260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08170_ _15521_/A hold2645/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08171_/B sky130_fd_sc_hd__mux2_1
X_17368_ _17978_/CLK _17368_/D vssd1 vssd1 vccd1 vccd1 _17368_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_49 _15555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16319_ _16319_/CLK _16319_/D vssd1 vssd1 vccd1 vccd1 _16319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17299_ _17299_/CLK _17299_/D vssd1 vssd1 vccd1 vccd1 hold770/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5006 _17560_/Q vssd1 vssd1 vccd1 vccd1 hold5006/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5017 _11704_/X vssd1 vssd1 vccd1 vccd1 _17058_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5028 _17159_/Q vssd1 vssd1 vccd1 vccd1 hold5028/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput101 _13113_/A vssd1 vssd1 vccd1 vccd1 hold5886/A sky130_fd_sc_hd__buf_6
XFILLER_0_141_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5039 _11077_/X vssd1 vssd1 vccd1 vccd1 _16849_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4305 _13846_/Y vssd1 vssd1 vccd1 vccd1 _17735_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput112 hold5933/X vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_12
Xoutput123 hold5959/X vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_12
Xhold4316 _12318_/Y vssd1 vssd1 vccd1 vccd1 _12319_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4327 _11205_/Y vssd1 vssd1 vccd1 vccd1 _11206_/B sky130_fd_sc_hd__dlygate4sd3_1
Xoutput134 hold5935/X vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_12
Xoutput145 hold5938/X vssd1 vssd1 vccd1 vccd1 hold5939/A sky130_fd_sc_hd__buf_6
XFILLER_0_100_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4338 _11766_/Y vssd1 vssd1 vccd1 vccd1 _11767_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3604 _16447_/Q vssd1 vssd1 vccd1 vccd1 hold3604/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4349 _11215_/Y vssd1 vssd1 vccd1 vccd1 _16895_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3615 _09760_/X vssd1 vssd1 vccd1 vccd1 _16410_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3626 _16628_/Q vssd1 vssd1 vccd1 vccd1 hold3626/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3637 _12566_/X vssd1 vssd1 vccd1 vccd1 _12567_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3648 _16359_/Q vssd1 vssd1 vccd1 vccd1 hold3648/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2903 _17757_/Q vssd1 vssd1 vccd1 vccd1 hold2903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3659 _09895_/X vssd1 vssd1 vccd1 vccd1 _16455_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2914 _16155_/Q vssd1 vssd1 vccd1 vccd1 hold2914/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2925 _09131_/X vssd1 vssd1 vccd1 vccd1 _16178_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2936 _18208_/Q vssd1 vssd1 vccd1 vccd1 hold2936/X sky130_fd_sc_hd__dlygate4sd3_1
X_07954_ _14517_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07954_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2947 _08243_/X vssd1 vssd1 vccd1 vccd1 _15756_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2958 _18223_/Q vssd1 vssd1 vccd1 vccd1 hold2958/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2969 _17954_/Q vssd1 vssd1 vccd1 vccd1 hold2969/X sky130_fd_sc_hd__dlygate4sd3_1
X_07885_ hold355/X _14789_/A vssd1 vssd1 vccd1 vccd1 _07916_/B sky130_fd_sc_hd__or2_4
XFILLER_0_177_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09624_ _09948_/A _09624_/B vssd1 vssd1 vccd1 vccd1 _09624_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_29_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_29_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_210_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09555_ _09957_/A _09555_/B vssd1 vssd1 vccd1 vccd1 _09555_/X sky130_fd_sc_hd__or2_1
XFILLER_0_167_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_37_wb_clk_i clkbuf_6_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18429_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_214_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08506_ hold2041/X _08503_/Y _08505_/X _13417_/C1 vssd1 vssd1 vccd1 vccd1 _08506_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09486_ hold1418/X hold5981/X _09485_/Y vssd1 vssd1 vccd1 vccd1 _16323_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08437_ _14330_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08437_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08368_ _15537_/A hold1081/X hold115/X vssd1 vssd1 vccd1 vccd1 _08369_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08299_ _14517_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08299_/X sky130_fd_sc_hd__or2_1
XFILLER_0_6_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10330_ hold4054/X _10616_/B _10329_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10330_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5540 _11356_/X vssd1 vssd1 vccd1 vccd1 _16942_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10261_ hold4573/X _10646_/B _10260_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10261_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5551 _16760_/Q vssd1 vssd1 vccd1 vccd1 hold5551/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5562 _11305_/X vssd1 vssd1 vccd1 vccd1 _16925_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5573 _17746_/Q vssd1 vssd1 vccd1 vccd1 hold5573/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12000_ _13797_/A _12000_/B vssd1 vssd1 vccd1 vccd1 _12000_/X sky130_fd_sc_hd__or2_1
Xhold5584 _11641_/X vssd1 vssd1 vccd1 vccd1 _17037_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4850 _09832_/X vssd1 vssd1 vccd1 vccd1 _16434_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5595 _17651_/Q vssd1 vssd1 vccd1 vccd1 hold5595/X sky130_fd_sc_hd__dlygate4sd3_1
X_10192_ hold4013/X _11186_/B _10191_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10192_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4861 _16869_/Q vssd1 vssd1 vccd1 vccd1 hold4861/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4872 _12232_/X vssd1 vssd1 vccd1 vccd1 _17234_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4883 _16982_/Q vssd1 vssd1 vccd1 vccd1 hold4883/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4894 _12130_/X vssd1 vssd1 vccd1 vccd1 _17200_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout350 _08930_/S vssd1 vssd1 vccd1 vccd1 _08932_/S sky130_fd_sc_hd__buf_8
XFILLER_0_219_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout361 _15560_/A2 vssd1 vssd1 vccd1 vccd1 _15547_/B sky130_fd_sc_hd__buf_4
XFILLER_0_205_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout372 _15020_/X vssd1 vssd1 vccd1 vccd1 _15071_/S sky130_fd_sc_hd__clkbuf_16
Xfanout383 _14830_/B vssd1 vssd1 vccd1 vccd1 _14840_/B sky130_fd_sc_hd__buf_8
X_13951_ hold1628/X _13995_/A2 _13950_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _13951_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout394 _14626_/Y vssd1 vssd1 vccd1 vccd1 _14666_/B sky130_fd_sc_hd__buf_8
XFILLER_0_57_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12902_ hold3305/X _12901_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12903_/B sky130_fd_sc_hd__mux2_1
X_16670_ _18164_/CLK _16670_/D vssd1 vssd1 vccd1 vccd1 _16670_/Q sky130_fd_sc_hd__dfxtp_1
X_13882_ _13888_/A _13882_/B vssd1 vssd1 vccd1 vccd1 _13882_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_202_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12833_ hold3965/X _12832_/X _12839_/S vssd1 vssd1 vccd1 vccd1 _12833_/X sky130_fd_sc_hd__mux2_1
X_15621_ _17154_/CLK _15621_/D vssd1 vssd1 vccd1 vccd1 _15621_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _18374_/CLK _18340_/D vssd1 vssd1 vccd1 vccd1 _18340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12764_ hold3769/X _12763_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12764_/X sky130_fd_sc_hd__mux2_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ hold2006/X _15560_/A2 _15551_/X _12849_/A vssd1 vssd1 vccd1 vccd1 _15552_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14503_ hold927/X _14553_/B vssd1 vssd1 vccd1 vccd1 _14503_/X sky130_fd_sc_hd__or2_1
X_11715_ _12093_/A _11715_/B vssd1 vssd1 vccd1 vccd1 _11715_/X sky130_fd_sc_hd__or2_1
X_15483_ hold764/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15483_/X sky130_fd_sc_hd__or2_1
X_18271_ _18271_/CLK _18271_/D vssd1 vssd1 vccd1 vccd1 _18271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ hold4074/X _12694_/X _12839_/S vssd1 vssd1 vccd1 vccd1 _12696_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_83_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17222_ _17222_/CLK _17222_/D vssd1 vssd1 vccd1 vccd1 _17222_/Q sky130_fd_sc_hd__dfxtp_1
X_14434_ hold2613/X _14433_/B _14433_/Y _14368_/A vssd1 vssd1 vccd1 vccd1 _14434_/X
+ sky130_fd_sc_hd__o211a_1
X_11646_ _12219_/A _11646_/B vssd1 vssd1 vccd1 vccd1 _11646_/X sky130_fd_sc_hd__or2_1
XFILLER_0_154_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput14 input14/A vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_1
XFILLER_0_126_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput25 hold85/X vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__buf_6
XFILLER_0_154_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14365_ _15099_/A hold2804/X _14381_/S vssd1 vssd1 vccd1 vccd1 _14366_/B sky130_fd_sc_hd__mux2_1
X_17153_ _17153_/CLK _17153_/D vssd1 vssd1 vccd1 vccd1 _17153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput36 input36/A vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11577_ _11694_/A _11577_/B vssd1 vssd1 vccd1 vccd1 _11577_/X sky130_fd_sc_hd__or2_1
XFILLER_0_108_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_414_wb_clk_i clkbuf_6_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18428_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xinput47 input47/A vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__buf_6
XFILLER_0_220_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16104_ _17331_/CLK _16104_/D vssd1 vssd1 vccd1 vccd1 _16104_/Q sky130_fd_sc_hd__dfxtp_1
Xinput58 input58/A vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__buf_6
X_13316_ hold1637/X hold4743/X _13796_/S vssd1 vssd1 vccd1 vccd1 _13317_/B sky130_fd_sc_hd__mux2_1
Xinput69 input69/A vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_1
X_10528_ hold3710/X _10649_/B _10527_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10528_/X
+ sky130_fd_sc_hd__o211a_1
X_17084_ _17900_/CLK _17084_/D vssd1 vssd1 vccd1 vccd1 _17084_/Q sky130_fd_sc_hd__dfxtp_1
Xhold809 hold809/A vssd1 vssd1 vccd1 vccd1 hold809/X sky130_fd_sc_hd__dlygate4sd3_1
X_14296_ hold945/X _14338_/B vssd1 vssd1 vccd1 vccd1 _14296_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13247_ _13311_/A1 _13245_/X _13246_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13247_/X
+ sky130_fd_sc_hd__o211a_1
X_16035_ _17314_/CLK _16035_/D vssd1 vssd1 vccd1 vccd1 hold890/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10459_ hold3895/X _10649_/B _10458_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10459_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13178_ _17573_/Q _17107_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13178_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12129_ _13314_/A _12129_/B vssd1 vssd1 vccd1 vccd1 _12129_/X sky130_fd_sc_hd__or2_1
XFILLER_0_100_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17986_ _18019_/CLK _17986_/D vssd1 vssd1 vccd1 vccd1 hold783/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1509 _18323_/Q vssd1 vssd1 vccd1 vccd1 hold1509/X sky130_fd_sc_hd__dlygate4sd3_1
X_16937_ _18432_/CLK _16937_/D vssd1 vssd1 vccd1 vccd1 _16937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16868_ _18073_/CLK _16868_/D vssd1 vssd1 vccd1 vccd1 _16868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15819_ _17726_/CLK _15819_/D vssd1 vssd1 vccd1 vccd1 hold613/A sky130_fd_sc_hd__dfxtp_1
X_16799_ _18194_/CLK _16799_/D vssd1 vssd1 vccd1 vccd1 _16799_/Q sky130_fd_sc_hd__dfxtp_1
X_09340_ _18460_/Q _07802_/B _15481_/A1 vssd1 vssd1 vccd1 vccd1 _09340_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09271_ hold235/X _16247_/Q hold271/X vssd1 vssd1 vccd1 vccd1 hold272/A sky130_fd_sc_hd__mux2_1
X_08222_ hold1291/X _08209_/B _08221_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _08222_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08153_ _08153_/A _08153_/B vssd1 vssd1 vccd1 vccd1 _15715_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_155_wb_clk_i clkbuf_6_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16098_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08084_ _15163_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08084_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_114_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4102 _11398_/X vssd1 vssd1 vccd1 vccd1 _16956_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4113 _16889_/Q vssd1 vssd1 vccd1 vccd1 hold4113/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_1384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4124 _13399_/X vssd1 vssd1 vccd1 vccd1 _17586_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4135 _16761_/Q vssd1 vssd1 vccd1 vccd1 hold4135/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4146 _09628_/X vssd1 vssd1 vccd1 vccd1 _16366_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3401 _12725_/X vssd1 vssd1 vccd1 vccd1 _12726_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3412 _10002_/Y vssd1 vssd1 vccd1 vccd1 _10003_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4157 _11389_/X vssd1 vssd1 vccd1 vccd1 _16953_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3423 _16523_/Q vssd1 vssd1 vccd1 vccd1 hold3423/X sky130_fd_sc_hd__clkbuf_2
Xhold4168 _10882_/X vssd1 vssd1 vccd1 vccd1 _16784_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3434 _10060_/Y vssd1 vssd1 vccd1 vccd1 _16510_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4179 _17032_/Q vssd1 vssd1 vccd1 vccd1 hold4179/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2700 _15013_/X vssd1 vssd1 vccd1 vccd1 _18292_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3445 _16329_/Q vssd1 vssd1 vccd1 vccd1 _13102_/A sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_5618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3456 _16332_/Q vssd1 vssd1 vccd1 vccd1 _13126_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2711 _17810_/Q vssd1 vssd1 vccd1 vccd1 hold2711/X sky130_fd_sc_hd__dlygate4sd3_1
X_08986_ _15491_/A _08986_/B vssd1 vssd1 vccd1 vccd1 _16110_/D sky130_fd_sc_hd__and2_1
XFILLER_0_228_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2722 _14641_/X vssd1 vssd1 vccd1 vccd1 _18113_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3467 _11776_/Y vssd1 vssd1 vccd1 vccd1 _17082_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2733 _15727_/Q vssd1 vssd1 vccd1 vccd1 hold2733/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3478 _11221_/Y vssd1 vssd1 vccd1 vccd1 _16897_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3489 _10608_/Y vssd1 vssd1 vccd1 vccd1 _10609_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2744 _14757_/X vssd1 vssd1 vccd1 vccd1 _18169_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2755 _09215_/X vssd1 vssd1 vccd1 vccd1 _16219_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07937_ hold1459/X _07924_/B _07936_/X _08167_/A vssd1 vssd1 vccd1 vccd1 _07937_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2766 _14635_/X vssd1 vssd1 vccd1 vccd1 _18110_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2777 _17941_/Q vssd1 vssd1 vccd1 vccd1 hold2777/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2788 _17787_/Q vssd1 vssd1 vccd1 vccd1 hold2788/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2799 _13981_/X vssd1 vssd1 vccd1 vccd1 _17797_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07868_ hold2439/X _07869_/B _07867_/Y _08131_/A vssd1 vssd1 vccd1 vccd1 _07868_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09607_ hold3911/X _10004_/B _09606_/X _15482_/A vssd1 vssd1 vccd1 vccd1 _09607_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07799_ _11158_/A _07799_/B vssd1 vssd1 vccd1 vccd1 _18460_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_6_1406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09538_ hold5837/X _10022_/B _09537_/X _15202_/C1 vssd1 vssd1 vccd1 vccd1 _09538_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09469_ hold739/X _09472_/C _09472_/D vssd1 vssd1 vccd1 vccd1 _09471_/B sky130_fd_sc_hd__and3_1
XFILLER_0_66_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11500_ hold5410/X _11786_/B _11499_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11500_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12480_ _17333_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12480_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11431_ hold5669/X _12299_/B _11430_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _11431_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14150_ _15549_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14150_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11362_ hold5235/X _11741_/B _11361_/X _14211_/C1 vssd1 vssd1 vccd1 vccd1 _11362_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13101_ _13100_/X hold3475/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13101_/X sky130_fd_sc_hd__mux2_1
Xhold6060 _18335_/Q vssd1 vssd1 vccd1 vccd1 hold6060/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10313_ hold1994/X _16595_/Q _10595_/C vssd1 vssd1 vccd1 vccd1 _10314_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_225_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6071 _18358_/Q vssd1 vssd1 vccd1 vccd1 hold6071/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6082 _18360_/Q vssd1 vssd1 vccd1 vccd1 hold6082/X sky130_fd_sc_hd__dlygate4sd3_1
X_14081_ hold2771/X _14094_/B _14080_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _14081_/X
+ sky130_fd_sc_hd__o211a_1
Xhold6093 _18419_/Q vssd1 vssd1 vccd1 vccd1 hold6093/X sky130_fd_sc_hd__dlygate4sd3_1
X_11293_ hold5693/X _11771_/B _11292_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _11293_/X
+ sky130_fd_sc_hd__o211a_1
X_13032_ _13056_/C hold896/X hold905/A vssd1 vssd1 vccd1 vccd1 _13032_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5370 _16977_/Q vssd1 vssd1 vccd1 vccd1 hold5370/X sky130_fd_sc_hd__dlygate4sd3_1
X_10244_ hold2643/X _16572_/Q _10628_/C vssd1 vssd1 vccd1 vccd1 _10245_/B sky130_fd_sc_hd__mux2_1
Xhold5381 _11839_/X vssd1 vssd1 vccd1 vccd1 _17103_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5392 _17086_/Q vssd1 vssd1 vccd1 vccd1 hold5392/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4680 _09610_/X vssd1 vssd1 vccd1 vccd1 _16360_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17840_ _17840_/CLK _17840_/D vssd1 vssd1 vccd1 vccd1 _17840_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4691 _16397_/Q vssd1 vssd1 vccd1 vccd1 hold4691/X sky130_fd_sc_hd__dlygate4sd3_1
X_10175_ hold1905/X _16549_/Q _10601_/C vssd1 vssd1 vccd1 vccd1 _10176_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_218_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3990 _13582_/X vssd1 vssd1 vccd1 vccd1 _17647_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17771_ _17771_/CLK _17771_/D vssd1 vssd1 vccd1 vccd1 _17771_/Q sky130_fd_sc_hd__dfxtp_1
X_14983_ hold1072/X hold447/X _14982_/X _15048_/A vssd1 vssd1 vccd1 vccd1 _14983_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout180 fanout210/X vssd1 vssd1 vccd1 vccd1 _11741_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_234_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout191 _13877_/B vssd1 vssd1 vccd1 vccd1 _13883_/B sky130_fd_sc_hd__clkbuf_8
X_16722_ _18020_/CLK _16722_/D vssd1 vssd1 vccd1 vccd1 _16722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13934_ _14543_/A hold1097/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13935_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16653_ _18211_/CLK _16653_/D vssd1 vssd1 vccd1 vccd1 _16653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13865_ _17742_/Q _13871_/B _13865_/C vssd1 vssd1 vccd1 vccd1 _13865_/X sky130_fd_sc_hd__and3_1
XFILLER_0_57_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15604_ _17910_/CLK _15604_/D vssd1 vssd1 vccd1 vccd1 _15604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12816_ _12837_/A _12816_/B vssd1 vssd1 vccd1 vccd1 _17448_/D sky130_fd_sc_hd__and2_1
XFILLER_0_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16584_ _18206_/CLK _16584_/D vssd1 vssd1 vccd1 vccd1 _16584_/Q sky130_fd_sc_hd__dfxtp_1
X_13796_ hold1672/X _17719_/Q _13796_/S vssd1 vssd1 vccd1 vccd1 _13797_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18323_ _18323_/CLK _18323_/D vssd1 vssd1 vccd1 vccd1 _18323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15535_ _15535_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15535_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12750_/A _12747_/B vssd1 vssd1 vccd1 vccd1 _17425_/D sky130_fd_sc_hd__and2_1
XFILLER_0_173_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ _18356_/CLK _18254_/D vssd1 vssd1 vccd1 vccd1 _18254_/Q sky130_fd_sc_hd__dfxtp_1
X_15466_ hold323/X _09386_/A _15484_/B1 hold610/X vssd1 vssd1 vccd1 vccd1 _15471_/B
+ sky130_fd_sc_hd__a22o_1
X_12678_ _12837_/A _12678_/B vssd1 vssd1 vccd1 vccd1 _17402_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17205_ _17269_/CLK _17205_/D vssd1 vssd1 vccd1 vccd1 _17205_/Q sky130_fd_sc_hd__dfxtp_1
X_11629_ hold5406/X _11726_/B _11628_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _11629_/X
+ sky130_fd_sc_hd__o211a_1
X_14417_ _14596_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14417_/X sky130_fd_sc_hd__or2_1
X_18185_ _18223_/CLK _18185_/D vssd1 vssd1 vccd1 vccd1 _18185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15397_ hold387/X _09357_/A _15484_/B1 _15897_/Q _15396_/X vssd1 vssd1 vccd1 vccd1
+ _15402_/B sky130_fd_sc_hd__a221o_2
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17136_ _17229_/CLK _17136_/D vssd1 vssd1 vccd1 vccd1 _17136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14348_ _14348_/A _14348_/B vssd1 vssd1 vccd1 vccd1 _17973_/D sky130_fd_sc_hd__and2_1
Xhold606 input10/X vssd1 vssd1 vccd1 vccd1 hold606/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold617 input16/X vssd1 vssd1 vccd1 vccd1 hold617/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap336 wire337/X vssd1 vssd1 vccd1 vccd1 fanout335/A sky130_fd_sc_hd__buf_2
Xhold628 hold628/A vssd1 vssd1 vccd1 vccd1 input42/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 hold639/A vssd1 vssd1 vccd1 vccd1 hold639/X sky130_fd_sc_hd__dlygate4sd3_1
X_17067_ _17883_/CLK _17067_/D vssd1 vssd1 vccd1 vccd1 _17067_/Q sky130_fd_sc_hd__dfxtp_1
X_14279_ hold2729/X _14272_/B _14278_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _14279_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16018_ _16125_/CLK _16018_/D vssd1 vssd1 vccd1 vccd1 hold747/A sky130_fd_sc_hd__dfxtp_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ hold245/X hold500/X _08866_/S vssd1 vssd1 vccd1 vccd1 _08841_/B sky130_fd_sc_hd__mux2_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2007 _15552_/X vssd1 vssd1 vccd1 vccd1 _18454_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2018 _08202_/X vssd1 vssd1 vccd1 vccd1 _15737_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2029 _17869_/Q vssd1 vssd1 vccd1 vccd1 hold2029/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1306 _08106_/X vssd1 vssd1 vccd1 vccd1 _08107_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08771_ hold5/X _16006_/Q _08779_/S vssd1 vssd1 vccd1 vccd1 hold123/A sky130_fd_sc_hd__mux2_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1317 _15676_/Q vssd1 vssd1 vccd1 vccd1 hold1317/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1328 _08273_/X vssd1 vssd1 vccd1 vccd1 _15771_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17969_ _18028_/CLK _17969_/D vssd1 vssd1 vccd1 vccd1 _17969_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1339 _09145_/X vssd1 vssd1 vccd1 vccd1 _16185_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09323_ _15545_/A _09323_/B vssd1 vssd1 vccd1 vccd1 _09323_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_165_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_336_wb_clk_i clkbuf_6_43_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17153_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ _12753_/A _09254_/B vssd1 vssd1 vccd1 vccd1 _16238_/D sky130_fd_sc_hd__and2_1
XFILLER_0_29_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08205_ _14194_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08205_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09185_ hold2625/X _09218_/B _09184_/X _12786_/A vssd1 vssd1 vccd1 vccd1 _09185_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08136_ hold384/X hold535/X hold108/X vssd1 vssd1 vccd1 vccd1 hold536/A sky130_fd_sc_hd__mux2_1
XFILLER_0_44_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08067_ hold2832/X _08097_/A2 _08066_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _08067_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3220 _17367_/Q vssd1 vssd1 vccd1 vccd1 hold3220/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3231 _12809_/X vssd1 vssd1 vccd1 vccd1 _12810_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3242 _17499_/Q vssd1 vssd1 vccd1 vccd1 hold3242/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3253 _16679_/Q vssd1 vssd1 vccd1 vccd1 _10565_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3264 _12608_/X vssd1 vssd1 vccd1 vccd1 _12609_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2530 _17864_/Q vssd1 vssd1 vccd1 vccd1 hold2530/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3275 _10093_/X vssd1 vssd1 vccd1 vccd1 _16521_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2541 _15812_/Q vssd1 vssd1 vccd1 vccd1 hold2541/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3286 _17377_/Q vssd1 vssd1 vccd1 vccd1 hold3286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3297 _10429_/X vssd1 vssd1 vccd1 vccd1 _16633_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_wb_clk_i clkbuf_6_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18051_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2552 _16238_/Q vssd1 vssd1 vccd1 vccd1 hold2552/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08969_ hold254/X _16102_/Q _08997_/S vssd1 vssd1 vccd1 vccd1 hold255/A sky130_fd_sc_hd__mux2_1
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2563 _09161_/X vssd1 vssd1 vccd1 vccd1 _16193_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2574 _14488_/X vssd1 vssd1 vccd1 vccd1 _18041_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1840 _14749_/X vssd1 vssd1 vccd1 vccd1 _18165_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2585 _18103_/Q vssd1 vssd1 vccd1 vccd1 hold2585/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2596 _18302_/Q vssd1 vssd1 vccd1 vccd1 hold2596/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1851 _17955_/Q vssd1 vssd1 vccd1 vccd1 hold1851/X sky130_fd_sc_hd__dlygate4sd3_1
X_11980_ hold5785/X _12362_/B _11979_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _11980_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1862 _15001_/X vssd1 vssd1 vccd1 vccd1 _18286_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1873 _17843_/Q vssd1 vssd1 vccd1 vccd1 hold1873/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1884 _08158_/X vssd1 vssd1 vccd1 vccd1 _08159_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1895 _16312_/Q vssd1 vssd1 vccd1 vccd1 _09456_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10931_ hold3091/X hold3820/X _11765_/C vssd1 vssd1 vccd1 vccd1 _10932_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_233_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13650_ _13752_/A _13650_/B vssd1 vssd1 vccd1 vccd1 _13650_/X sky130_fd_sc_hd__or2_1
X_10862_ hold1777/X hold4127/X _11723_/C vssd1 vssd1 vccd1 vccd1 _10863_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_196_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12601_ _16276_/Q hold3265/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12601_/X sky130_fd_sc_hd__mux2_1
X_13581_ _13581_/A _13581_/B vssd1 vssd1 vccd1 vccd1 _13581_/X sky130_fd_sc_hd__or2_1
XFILLER_0_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ hold1875/X hold4853/X _11171_/C vssd1 vssd1 vccd1 vccd1 _10794_/B sky130_fd_sc_hd__mux2_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15320_ hold498/X _15448_/A2 _15446_/B1 hold806/X vssd1 vssd1 vccd1 vccd1 _15320_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12532_ hold2378/X _17355_/Q _12925_/S vssd1 vssd1 vccd1 vccd1 _12532_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12463_ hold452/X _12445_/A _12445_/B _12462_/X _15491_/A vssd1 vssd1 vccd1 vccd1
+ hold204/A sky130_fd_sc_hd__o311a_1
X_15251_ _16289_/Q _15477_/A2 _15487_/B1 hold675/X _15250_/X vssd1 vssd1 vccd1 vccd1
+ _15252_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_192_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11414_ hold2711/X _16962_/Q _12173_/S vssd1 vssd1 vccd1 vccd1 _11415_/B sky130_fd_sc_hd__mux2_1
X_14202_ _15221_/A _14202_/B vssd1 vssd1 vccd1 vccd1 _14202_/Y sky130_fd_sc_hd__nand2_1
X_15182_ _15182_/A _15182_/B vssd1 vssd1 vccd1 vccd1 _15227_/B sky130_fd_sc_hd__or2_4
XFILLER_0_227_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12394_ _12394_/A _12394_/B vssd1 vssd1 vccd1 vccd1 _17290_/D sky130_fd_sc_hd__and2_1
XFILLER_0_2_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14133_ hold6051/X _14148_/B hold521/X _13933_/A vssd1 vssd1 vccd1 vccd1 hold522/A
+ sky130_fd_sc_hd__o211a_1
X_11345_ hold2788/X hold4901/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11346_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_162_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14064_ _14457_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14064_/X sky130_fd_sc_hd__or2_1
X_11276_ hold2930/X hold4549/X _12242_/S vssd1 vssd1 vccd1 vccd1 _11277_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13015_ _15519_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13015_/X sky130_fd_sc_hd__or2_1
X_10227_ _10413_/A _10227_/B vssd1 vssd1 vccd1 vccd1 _10227_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_234_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17823_ _17823_/CLK _17823_/D vssd1 vssd1 vccd1 vccd1 _17823_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10158_ _10524_/A _10158_/B vssd1 vssd1 vccd1 vccd1 _10158_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17754_ _17754_/CLK _17754_/D vssd1 vssd1 vccd1 vccd1 _17754_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_5993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10089_ _10476_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10089_/X sky130_fd_sc_hd__or2_1
X_14966_ hold445/X _15182_/B vssd1 vssd1 vccd1 vccd1 hold446/A sky130_fd_sc_hd__nor2_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16705_ _18232_/CLK _16705_/D vssd1 vssd1 vccd1 vccd1 _16705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13917_ _13917_/A _13917_/B vssd1 vssd1 vccd1 vccd1 _17766_/D sky130_fd_sc_hd__and2_1
X_17685_ _17746_/CLK _17685_/D vssd1 vssd1 vccd1 vccd1 _17685_/Q sky130_fd_sc_hd__dfxtp_1
X_14897_ _14897_/A _15182_/B vssd1 vssd1 vccd1 vccd1 _14910_/B sky130_fd_sc_hd__or2_2
XFILLER_0_162_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16636_ _18226_/CLK _16636_/D vssd1 vssd1 vccd1 vccd1 _16636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13848_ hold3527/X _13581_/A _13847_/X vssd1 vssd1 vccd1 vccd1 _13848_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16567_ _18125_/CLK _16567_/D vssd1 vssd1 vccd1 vccd1 _16567_/Q sky130_fd_sc_hd__dfxtp_1
X_13779_ _13788_/A _13779_/B vssd1 vssd1 vccd1 vccd1 _13779_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18306_ _18368_/CLK _18306_/D vssd1 vssd1 vccd1 vccd1 _18306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15518_ hold2331/X _15560_/A2 _15517_/X _12864_/A vssd1 vssd1 vccd1 vccd1 _15518_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16498_ _18379_/CLK _16498_/D vssd1 vssd1 vccd1 vccd1 _16498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18237_ _18271_/CLK _18237_/D vssd1 vssd1 vccd1 vccd1 _18237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15449_ _15958_/Q _15484_/A2 _15447_/X vssd1 vssd1 vccd1 vccd1 _15452_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_170_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18168_ _18168_/CLK _18168_/D vssd1 vssd1 vccd1 vccd1 _18168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold403 hold403/A vssd1 vssd1 vccd1 vccd1 input56/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold414 hold414/A vssd1 vssd1 vccd1 vccd1 hold414/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17119_ _17247_/CLK _17119_/D vssd1 vssd1 vccd1 vccd1 _17119_/Q sky130_fd_sc_hd__dfxtp_1
Xhold425 hold425/A vssd1 vssd1 vccd1 vccd1 hold425/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 hold40/X vssd1 vssd1 vccd1 vccd1 input22/A sky130_fd_sc_hd__dlygate4sd3_1
X_18099_ _18099_/CLK _18099_/D vssd1 vssd1 vccd1 vccd1 _18099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold447 hold447/A vssd1 vssd1 vccd1 vccd1 hold447/X sky130_fd_sc_hd__buf_8
Xhold458 hold458/A vssd1 vssd1 vccd1 vccd1 hold458/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09941_ hold1199/X _16471_/Q _10049_/C vssd1 vssd1 vccd1 vccd1 _09942_/B sky130_fd_sc_hd__mux2_1
Xhold469 hold469/A vssd1 vssd1 vccd1 vccd1 hold469/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout905 hold579/X vssd1 vssd1 vccd1 vccd1 _14732_/A sky130_fd_sc_hd__buf_12
Xfanout916 hold1137/X vssd1 vssd1 vccd1 vccd1 hold1138/A sky130_fd_sc_hd__buf_6
Xfanout927 hold1253/X vssd1 vssd1 vccd1 vccd1 _15539_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_239_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09872_ hold2157/X hold3744/X _10067_/C vssd1 vssd1 vccd1 vccd1 _09873_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_141_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout938 hold1075/X vssd1 vssd1 vccd1 vccd1 hold1076/A sky130_fd_sc_hd__buf_6
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08823_ _15414_/A hold831/X vssd1 vssd1 vccd1 vccd1 _16030_/D sky130_fd_sc_hd__and2_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 _15638_/Q vssd1 vssd1 vccd1 vccd1 hold1103/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1114 _14751_/X vssd1 vssd1 vccd1 vccd1 _18166_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1125 _15833_/Q vssd1 vssd1 vccd1 vccd1 hold1125/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 hold1222/X vssd1 vssd1 vccd1 vccd1 hold1223/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08754_ _15284_/A hold480/X vssd1 vssd1 vccd1 vccd1 _15997_/D sky130_fd_sc_hd__and2_1
Xhold1147 input40/X vssd1 vssd1 vccd1 vccd1 hold1147/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1158 _14993_/X vssd1 vssd1 vccd1 vccd1 _18282_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1169 _17994_/Q vssd1 vssd1 vccd1 vccd1 hold1169/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_240_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ hold23/X hold513/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08686_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_240_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_170_wb_clk_i clkbuf_6_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18049_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_222_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09306_ hold1990/X _09323_/B _09305_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _09306_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09237_ _15513_/A hold2564/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09238_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09168_ hold992/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09168_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08119_ _08119_/A hold942/X vssd1 vssd1 vccd1 vccd1 _15698_/D sky130_fd_sc_hd__and2_1
XFILLER_0_47_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09099_ hold1931/X _09102_/B _09098_/X _12978_/A vssd1 vssd1 vccd1 vccd1 _09099_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11130_ _11670_/A _11130_/B vssd1 vssd1 vccd1 vccd1 _11130_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold970 hold970/A vssd1 vssd1 vccd1 vccd1 hold970/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 hold981/A vssd1 vssd1 vccd1 vccd1 hold981/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11061_ _11061_/A _11061_/B vssd1 vssd1 vccd1 vccd1 _11061_/X sky130_fd_sc_hd__or2_1
Xhold992 hold992/A vssd1 vssd1 vccd1 vccd1 hold992/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3050 _14117_/X vssd1 vssd1 vccd1 vccd1 _17862_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10012_ _11158_/A _10012_/B vssd1 vssd1 vccd1 vccd1 _16494_/D sky130_fd_sc_hd__nor2_1
Xhold3061 _17891_/Q vssd1 vssd1 vccd1 vccd1 hold3061/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3072 _18279_/Q vssd1 vssd1 vccd1 vccd1 hold3072/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3083 _14699_/X vssd1 vssd1 vccd1 vccd1 _18141_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3094 _14520_/X vssd1 vssd1 vccd1 vccd1 _18056_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2360 _08089_/X vssd1 vssd1 vccd1 vccd1 _15684_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ _15213_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14820_/X sky130_fd_sc_hd__or2_1
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2371 _16180_/Q vssd1 vssd1 vccd1 vccd1 hold2371/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2382 _16153_/Q vssd1 vssd1 vccd1 vccd1 hold2382/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2393 _14404_/X vssd1 vssd1 vccd1 vccd1 _18000_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1670 _17929_/Q vssd1 vssd1 vccd1 vccd1 hold1670/X sky130_fd_sc_hd__dlygate4sd3_1
X_14751_ hold1113/X _14774_/B _14750_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14751_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1681 _08206_/X vssd1 vssd1 vccd1 vccd1 _15739_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1692 _18184_/Q vssd1 vssd1 vccd1 vccd1 hold1692/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11963_ hold1513/X hold5741/X _13463_/S vssd1 vssd1 vccd1 vccd1 _11964_/B sky130_fd_sc_hd__mux2_1
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_258_wb_clk_i clkbuf_6_58_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18067_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ hold5169/X _13814_/B _13701_/X _13801_/C1 vssd1 vssd1 vccd1 vccd1 _13702_/X
+ sky130_fd_sc_hd__o211a_1
X_10914_ _11010_/A _10914_/B vssd1 vssd1 vccd1 vccd1 _10914_/X sky130_fd_sc_hd__or2_1
X_17470_ _17471_/CLK _17470_/D vssd1 vssd1 vccd1 vccd1 _17470_/Q sky130_fd_sc_hd__dfxtp_1
X_14682_ hold927/X _14732_/B vssd1 vssd1 vccd1 vccd1 _14682_/X sky130_fd_sc_hd__or2_1
XFILLER_0_169_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11894_ hold1079/X hold4387/X _13748_/S vssd1 vssd1 vccd1 vccd1 _11895_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16421_ _18334_/CLK _16421_/D vssd1 vssd1 vccd1 vccd1 _16421_/Q sky130_fd_sc_hd__dfxtp_1
X_10845_ _11649_/A _10845_/B vssd1 vssd1 vccd1 vccd1 _10845_/X sky130_fd_sc_hd__or2_1
X_13633_ hold4779/X _13862_/B _13632_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _13633_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16352_ _16480_/CLK _16352_/D vssd1 vssd1 vccd1 vccd1 _16352_/Q sky130_fd_sc_hd__dfxtp_1
X_10776_ _11067_/A _10776_/B vssd1 vssd1 vccd1 vccd1 _10776_/X sky130_fd_sc_hd__or2_1
X_13564_ hold5557/X _13880_/B _13563_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13564_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15303_ _15490_/A1 _15295_/X _15302_/X _15490_/B1 hold5925/A vssd1 vssd1 vccd1 vccd1
+ _15303_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_87_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12515_ _07826_/A _12514_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12516_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16283_ _17750_/CLK _16283_/D vssd1 vssd1 vccd1 vccd1 _16283_/Q sky130_fd_sc_hd__dfxtp_4
X_13495_ hold4125/X _13880_/B _13494_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _13495_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18022_ _18054_/CLK _18022_/D vssd1 vssd1 vccd1 vccd1 _18022_/Q sky130_fd_sc_hd__dfxtp_1
X_12446_ _17316_/Q _12506_/B vssd1 vssd1 vccd1 vccd1 _12446_/X sky130_fd_sc_hd__or2_1
X_15234_ hold1803/X _15221_/B _15233_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _15234_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15165_ _15165_/A _15165_/B vssd1 vssd1 vccd1 vccd1 _15165_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_140_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12377_ _17283_/Q _13886_/B _13886_/C vssd1 vssd1 vccd1 vccd1 _12377_/X sky130_fd_sc_hd__and3_1
XFILLER_0_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_239_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ _12093_/A _11328_/B vssd1 vssd1 vccd1 vccd1 _11328_/X sky130_fd_sc_hd__or2_1
X_14116_ _15189_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14116_/X sky130_fd_sc_hd__or2_1
XFILLER_0_240_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15096_ hold1213/X hold340/X _15095_/X _15212_/C1 vssd1 vssd1 vccd1 vccd1 _15096_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_240_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14047_ hold2967/X _14040_/B _14046_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _14047_/X
+ sky130_fd_sc_hd__o211a_1
X_11259_ _11649_/A _11259_/B vssd1 vssd1 vccd1 vccd1 _11259_/X sky130_fd_sc_hd__or2_1
XFILLER_0_240_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17806_ _17838_/CLK _17806_/D vssd1 vssd1 vccd1 vccd1 _17806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15998_ _16058_/CLK _15998_/D vssd1 vssd1 vccd1 vccd1 hold766/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17737_ _17737_/CLK _17737_/D vssd1 vssd1 vccd1 vccd1 _17737_/Q sky130_fd_sc_hd__dfxtp_1
X_14949_ hold996/X _14952_/B _14948_/Y _15226_/C1 vssd1 vssd1 vccd1 vccd1 hold997/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08470_ _15203_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08470_/X sky130_fd_sc_hd__or2_1
X_17668_ _17732_/CLK _17668_/D vssd1 vssd1 vccd1 vccd1 _17668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16619_ _18217_/CLK _16619_/D vssd1 vssd1 vccd1 vccd1 _16619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17599_ _17599_/CLK _17599_/D vssd1 vssd1 vccd1 vccd1 _17599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09022_ hold163/X hold433/X _09060_/S vssd1 vssd1 vccd1 vccd1 hold434/A sky130_fd_sc_hd__mux2_1
XFILLER_0_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5903 hold6033/X vssd1 vssd1 vccd1 vccd1 _13073_/A sky130_fd_sc_hd__buf_1
Xhold5914 hold5914/A vssd1 vssd1 vccd1 vccd1 hold5914/X sky130_fd_sc_hd__buf_2
Xhold200 hold200/A vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold211 hold211/A vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5925 hold5925/A vssd1 vssd1 vccd1 vccd1 hold5925/X sky130_fd_sc_hd__buf_2
Xhold5936 _16282_/Q vssd1 vssd1 vccd1 vccd1 hold5936/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold222 hold222/A vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5947 hold6091/X vssd1 vssd1 vccd1 vccd1 hold5947/X sky130_fd_sc_hd__clkbuf_4
Xhold5958 _18424_/Q vssd1 vssd1 vccd1 vccd1 hold5958/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 hold96/X vssd1 vssd1 vccd1 vccd1 input47/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 input14/X vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__buf_1
Xhold255 hold255/A vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5969 hold5969/A vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_12
Xhold266 hold350/X vssd1 vssd1 vccd1 vccd1 hold351/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 input29/X vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold288 input53/X vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__clkbuf_2
Xfanout702 _09047_/A vssd1 vssd1 vccd1 vccd1 _12416_/A sky130_fd_sc_hd__clkbuf_4
X_09924_ _10560_/A _09924_/B vssd1 vssd1 vccd1 vccd1 _09924_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold299 hold299/A vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout713 _15491_/A vssd1 vssd1 vccd1 vccd1 _12440_/A sky130_fd_sc_hd__buf_2
XFILLER_0_102_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout724 _15176_/C1 vssd1 vssd1 vccd1 vccd1 _15404_/A sky130_fd_sc_hd__buf_2
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout735 _09907_/C1 vssd1 vssd1 vccd1 vccd1 _08954_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_238_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout746 fanout843/X vssd1 vssd1 vccd1 vccd1 _08111_/A sky130_fd_sc_hd__clkbuf_4
X_09855_ _09978_/A _09855_/B vssd1 vssd1 vccd1 vccd1 _09855_/X sky130_fd_sc_hd__or2_1
Xfanout757 _14380_/A vssd1 vssd1 vccd1 vccd1 _13909_/A sky130_fd_sc_hd__buf_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout768 fanout791/X vssd1 vssd1 vccd1 vccd1 _13684_/C1 sky130_fd_sc_hd__buf_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout779 _13917_/A vssd1 vssd1 vccd1 vccd1 _13941_/A sky130_fd_sc_hd__buf_4
XFILLER_0_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ hold618/X hold794/X _08866_/S vssd1 vssd1 vccd1 vccd1 hold795/A sky130_fd_sc_hd__mux2_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09786_ _09954_/A _09786_/B vssd1 vssd1 vccd1 vccd1 _09786_/X sky130_fd_sc_hd__or2_1
XFILLER_0_213_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08737_ hold684/X hold823/X _08793_/S vssd1 vssd1 vccd1 vccd1 hold824/A sky130_fd_sc_hd__mux2_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_106 _11203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_351_wb_clk_i clkbuf_6_40_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17716_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 hold915/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_128 _15173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08668_ _12426_/A hold792/X vssd1 vssd1 vccd1 vccd1 _15955_/D sky130_fd_sc_hd__and2_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_233_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ hold226/X hold722/X _08657_/S vssd1 vssd1 vccd1 vccd1 hold723/A sky130_fd_sc_hd__mux2_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10630_ _11206_/A _10630_/B vssd1 vssd1 vccd1 vccd1 _16700_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_14_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10561_ hold3930/X _10568_/B _10560_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _16677_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_1231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12300_ hold4762/X _12210_/A _12299_/X vssd1 vssd1 vccd1 vccd1 _12300_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13280_ _13273_/X _13279_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17553_/D sky130_fd_sc_hd__o21a_1
X_10492_ hold3940/X _10625_/B _10491_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10492_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12231_ _13482_/A _12231_/B vssd1 vssd1 vccd1 vccd1 _12231_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12162_ _13314_/A _12162_/B vssd1 vssd1 vccd1 vccd1 _12162_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11113_ _11207_/A _11222_/B _11112_/X _14526_/C1 vssd1 vssd1 vccd1 vccd1 _11113_/X
+ sky130_fd_sc_hd__o211a_1
X_12093_ _12093_/A _12093_/B vssd1 vssd1 vccd1 vccd1 _12093_/X sky130_fd_sc_hd__or2_1
X_16970_ _17850_/CLK _16970_/D vssd1 vssd1 vccd1 vccd1 _16970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15921_ _17320_/CLK _15921_/D vssd1 vssd1 vccd1 vccd1 hold490/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11044_ hold5273/X _11732_/B _11043_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _11044_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_217_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_439_wb_clk_i clkbuf_6_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17624_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15852_ _17672_/CLK _15852_/D vssd1 vssd1 vccd1 vccd1 _15852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2190 _14085_/X vssd1 vssd1 vccd1 vccd1 _17847_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14803_ hold1978/X _14826_/B _14802_/X _14853_/C1 vssd1 vssd1 vccd1 vccd1 _14803_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _17747_/CLK _15783_/D vssd1 vssd1 vccd1 vccd1 _15783_/Q sky130_fd_sc_hd__dfxtp_1
X_12995_ hold4747/X _12994_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12995_/X sky130_fd_sc_hd__mux2_1
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ _17523_/CLK _17522_/D vssd1 vssd1 vccd1 vccd1 _17522_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14734_ _14735_/A _14843_/B vssd1 vssd1 vccd1 vccd1 _14734_/Y sky130_fd_sc_hd__nor2_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11946_ _12234_/A _11946_/B vssd1 vssd1 vccd1 vccd1 _11946_/X sky130_fd_sc_hd__or2_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17453_ _17456_/CLK _17453_/D vssd1 vssd1 vccd1 vccd1 _17453_/Q sky130_fd_sc_hd__dfxtp_1
X_14665_ hold2689/X _14666_/B _14664_/Y _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14665_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _13482_/A _11877_/B vssd1 vssd1 vccd1 vccd1 _11877_/X sky130_fd_sc_hd__or2_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16404_ _18381_/CLK _16404_/D vssd1 vssd1 vccd1 vccd1 _16404_/Q sky130_fd_sc_hd__dfxtp_1
X_13616_ hold2669/X _17659_/Q _13817_/C vssd1 vssd1 vccd1 vccd1 _13617_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10828_ hold4081/X _11210_/B _10827_/X _14528_/C1 vssd1 vssd1 vccd1 vccd1 _10828_/X
+ sky130_fd_sc_hd__o211a_1
X_17384_ _18437_/CLK _17384_/D vssd1 vssd1 vccd1 vccd1 _17384_/Q sky130_fd_sc_hd__dfxtp_1
X_14596_ _14596_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14596_/X sky130_fd_sc_hd__or2_1
XFILLER_0_184_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16335_ _18250_/CLK _16335_/D vssd1 vssd1 vccd1 vccd1 _16335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13547_ _15821_/Q hold5046/X _13871_/C vssd1 vssd1 vccd1 vccd1 _13548_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_171_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10759_ hold3842/X _11144_/B _10758_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _10759_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16266_ _17978_/CLK _16266_/D vssd1 vssd1 vccd1 vccd1 _16266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13478_ hold2542/X _17613_/Q _13766_/S vssd1 vssd1 vccd1 vccd1 _13479_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_207_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18005_ _18005_/CLK _18005_/D vssd1 vssd1 vccd1 vccd1 _18005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15217_ _15217_/A _15221_/B vssd1 vssd1 vccd1 vccd1 _15217_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12429_ hold143/X hold653/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12430_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_113_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16197_ _17477_/CLK _16197_/D vssd1 vssd1 vccd1 vccd1 _16197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4509 _16428_/Q vssd1 vssd1 vccd1 vccd1 hold4509/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15148_ hold3080/X _15167_/B _15147_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _15148_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3808 _16851_/Q vssd1 vssd1 vccd1 vccd1 hold3808/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3819 _11938_/X vssd1 vssd1 vccd1 vccd1 _17136_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07970_ _15539_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07970_/X sky130_fd_sc_hd__or2_1
X_15079_ _15187_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15079_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09640_ hold4974/X _11171_/B _09639_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _09640_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_109_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17297_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09571_ hold3237/X _10046_/B _09570_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09571_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_6_19_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_19_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08522_ hold937/X _17519_/Q vssd1 vssd1 vccd1 vccd1 _13046_/C sky130_fd_sc_hd__nand2b_1
XFILLER_0_222_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08453_ hold1395/X _08488_/B _08452_/X _13795_/C1 vssd1 vssd1 vccd1 vccd1 _08453_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08384_ _14726_/A hold2661/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08385_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_45_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09005_ _15434_/A hold176/X vssd1 vssd1 vccd1 vccd1 _16119_/D sky130_fd_sc_hd__and2_1
XFILLER_0_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5700 _11851_/X vssd1 vssd1 vccd1 vccd1 _17107_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5711 _17110_/Q vssd1 vssd1 vccd1 vccd1 hold5711/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5722 _13807_/Y vssd1 vssd1 vccd1 vccd1 _17722_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5733 _17640_/Q vssd1 vssd1 vccd1 vccd1 hold5733/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5744 _12046_/X vssd1 vssd1 vccd1 vccd1 _17172_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5755 _17241_/Q vssd1 vssd1 vccd1 vccd1 hold5755/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5766 _11965_/X vssd1 vssd1 vccd1 vccd1 _17145_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5777 _17693_/Q vssd1 vssd1 vccd1 vccd1 hold5777/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5788 _13516_/X vssd1 vssd1 vccd1 vccd1 _17625_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5799 _17146_/Q vssd1 vssd1 vccd1 vccd1 hold5799/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout510 _10475_/S vssd1 vssd1 vccd1 vccd1 _10067_/C sky130_fd_sc_hd__clkbuf_8
Xclkbuf_6_58_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_58_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout521 _09499_/Y vssd1 vssd1 vccd1 vccd1 _10619_/C sky130_fd_sc_hd__clkbuf_8
X_09907_ hold3525/X _10025_/B _09906_/X _09907_/C1 vssd1 vssd1 vccd1 vccd1 _09907_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout532 _09156_/B vssd1 vssd1 vccd1 vccd1 _09176_/B sky130_fd_sc_hd__buf_4
Xfanout543 _08448_/Y vssd1 vssd1 vccd1 vccd1 _08488_/B sky130_fd_sc_hd__clkbuf_8
Xfanout554 _08228_/Y vssd1 vssd1 vccd1 vccd1 _08268_/B sky130_fd_sc_hd__buf_8
Xfanout565 _07993_/Y vssd1 vssd1 vccd1 vccd1 _08029_/B sky130_fd_sc_hd__buf_8
Xfanout576 _14622_/B vssd1 vssd1 vccd1 vccd1 _14624_/B sky130_fd_sc_hd__clkbuf_8
Xfanout587 _13305_/B vssd1 vssd1 vccd1 vccd1 _13185_/B sky130_fd_sc_hd__buf_4
X_09838_ hold4547/X _10028_/B _09837_/X _15048_/A vssd1 vssd1 vccd1 vccd1 _09838_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout598 _12985_/S vssd1 vssd1 vccd1 vccd1 _12925_/S sky130_fd_sc_hd__buf_6
XFILLER_0_38_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_1260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09769_ hold3612/X _10049_/B _09768_/X _15212_/C1 vssd1 vssd1 vccd1 vccd1 _09769_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _12337_/A _11800_/B vssd1 vssd1 vccd1 vccd1 _11800_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_213_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12780_ _12786_/A _12780_/B vssd1 vssd1 vccd1 vccd1 _17436_/D sky130_fd_sc_hd__and2_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_213_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _12301_/A _11731_/B vssd1 vssd1 vccd1 vccd1 _17067_/D sky130_fd_sc_hd__nor2_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14450_ hold2171/X _14487_/B _14449_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _14450_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11662_ hold5408/X _11195_/B _11661_/X _14462_/C1 vssd1 vssd1 vccd1 vccd1 _11662_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13401_ _13791_/A _13401_/B vssd1 vssd1 vccd1 vccd1 _13401_/X sky130_fd_sc_hd__or2_1
X_10613_ _16695_/Q _10637_/B _10619_/C vssd1 vssd1 vccd1 vccd1 _10613_/X sky130_fd_sc_hd__and3_1
X_14381_ _15169_/A hold1406/X _14381_/S vssd1 vssd1 vccd1 vccd1 _14382_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11593_ hold5677/X _11786_/B _11592_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _11593_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16120_ _16120_/CLK _16120_/D vssd1 vssd1 vccd1 vccd1 hold835/A sky130_fd_sc_hd__dfxtp_1
X_10544_ hold1060/X hold3610/X _10646_/C vssd1 vssd1 vccd1 vccd1 _10545_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_135_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13332_ _13716_/A _13332_/B vssd1 vssd1 vccd1 vccd1 _13332_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16051_ _18308_/CLK _16051_/D vssd1 vssd1 vccd1 vccd1 hold401/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13263_ _13311_/A1 _13261_/X _13262_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13263_/X
+ sky130_fd_sc_hd__o211a_1
X_10475_ hold2865/X _16649_/Q _10475_/S vssd1 vssd1 vccd1 vccd1 _10476_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15002_ _15217_/A hold447/X vssd1 vssd1 vccd1 vccd1 _15002_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_150_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12214_ hold4561/X _12308_/B _12213_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _12214_/X
+ sky130_fd_sc_hd__o211a_1
X_13194_ _17575_/Q _17109_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13194_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_206_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_7_wb_clk_i clkbuf_6_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17450_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12145_ hold5468/X _12335_/B _12144_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _12145_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12076_ hold5789/X _12362_/B _12075_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _12076_/X
+ sky130_fd_sc_hd__o211a_1
X_16953_ _17894_/CLK _16953_/D vssd1 vssd1 vccd1 vccd1 _16953_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_273_wb_clk_i clkbuf_6_51_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18214_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_237_1319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15904_ _17322_/CLK _15904_/D vssd1 vssd1 vccd1 vccd1 hold610/A sky130_fd_sc_hd__dfxtp_1
X_11027_ hold1407/X _16833_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _11028_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16884_ _18063_/CLK _16884_/D vssd1 vssd1 vccd1 vccd1 _16884_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_202_wb_clk_i clkbuf_6_55_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18388_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_194_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15835_ _17718_/CLK _15835_/D vssd1 vssd1 vccd1 vccd1 _15835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_235_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15766_ _17653_/CLK _15766_/D vssd1 vssd1 vccd1 vccd1 _15766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12978_ _12978_/A _12978_/B vssd1 vssd1 vccd1 vccd1 _17502_/D sky130_fd_sc_hd__and2_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _17506_/CLK _17505_/D vssd1 vssd1 vccd1 vccd1 _17505_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14717_ hold2302/X _14720_/B _14716_/Y _14895_/C1 vssd1 vssd1 vccd1 vccd1 _14717_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_234_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11929_ hold4026/X _12356_/B _11928_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _11929_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_185_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15697_ _17900_/CLK _15697_/D vssd1 vssd1 vccd1 vccd1 _15697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17436_ _17437_/CLK _17436_/D vssd1 vssd1 vccd1 vccd1 _17436_/Q sky130_fd_sc_hd__dfxtp_1
X_14648_ _14988_/A _14672_/B vssd1 vssd1 vccd1 vccd1 _14648_/X sky130_fd_sc_hd__or2_1
XFILLER_0_172_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_17 _13132_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_28 _13180_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 _13260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ _17514_/CLK _17367_/D vssd1 vssd1 vccd1 vccd1 _17367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14579_ hold1728/X _14610_/B _14578_/X _14893_/C1 vssd1 vssd1 vccd1 vccd1 _14579_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16318_ _16319_/CLK _16318_/D vssd1 vssd1 vccd1 vccd1 hold733/A sky130_fd_sc_hd__dfxtp_1
X_17298_ _17319_/CLK _17298_/D vssd1 vssd1 vccd1 vccd1 hold781/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5007 _13801_/X vssd1 vssd1 vccd1 vccd1 _17720_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16249_ _17445_/CLK _16249_/D vssd1 vssd1 vccd1 vccd1 _16249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5018 _16771_/Q vssd1 vssd1 vccd1 vccd1 hold5018/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5029 _11911_/X vssd1 vssd1 vccd1 vccd1 _17127_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput102 _13121_/A vssd1 vssd1 vccd1 vccd1 hold5888/A sky130_fd_sc_hd__buf_6
XFILLER_0_141_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput113 hold5914/X vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_12
Xhold4306 _17111_/Q vssd1 vssd1 vccd1 vccd1 hold4306/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput124 hold5974/X vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_12
Xhold4317 _12319_/Y vssd1 vssd1 vccd1 vccd1 _17263_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4328 _16713_/Q vssd1 vssd1 vccd1 vccd1 hold4328/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput135 hold5925/X vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_12
Xoutput146 _18463_/X vssd1 vssd1 vccd1 vccd1 slv_enable sky130_fd_sc_hd__buf_12
Xhold4339 _11767_/Y vssd1 vssd1 vccd1 vccd1 _17079_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3605 _09775_/X vssd1 vssd1 vccd1 vccd1 _16415_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_227_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3616 _16552_/Q vssd1 vssd1 vccd1 vccd1 hold3616/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3627 _10318_/X vssd1 vssd1 vccd1 vccd1 _16596_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3638 _17352_/Q vssd1 vssd1 vccd1 vccd1 hold3638/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2904 _18443_/Q vssd1 vssd1 vccd1 vccd1 hold2904/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3649 _09511_/X vssd1 vssd1 vccd1 vccd1 _16327_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2915 _09081_/X vssd1 vssd1 vccd1 vccd1 _16155_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2926 _16257_/Q vssd1 vssd1 vccd1 vccd1 hold2926/X sky130_fd_sc_hd__dlygate4sd3_1
X_07953_ hold2910/X _07991_/A2 _07952_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _07953_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2937 _14837_/X vssd1 vssd1 vccd1 vccd1 _18208_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2948 _18379_/Q vssd1 vssd1 vccd1 vccd1 hold2948/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2959 _14869_/X vssd1 vssd1 vccd1 vccd1 _18223_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07884_ hold355/X _14789_/A vssd1 vssd1 vccd1 vccd1 _07884_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_39_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09623_ hold3102/X hold4591/X _10031_/C vssd1 vssd1 vccd1 vccd1 _09624_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_207_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09554_ hold1315/X _13206_/A _10040_/C vssd1 vssd1 vccd1 vccd1 _09555_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_214_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08505_ _14164_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08505_/X sky130_fd_sc_hd__or2_1
X_09485_ hold1418/X hold5981/X _09478_/B vssd1 vssd1 vccd1 vccd1 _09485_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_92_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08436_ hold1227/X _08433_/B _08435_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08436_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_77_wb_clk_i clkbuf_6_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17513_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08367_ _08367_/A _08367_/B vssd1 vssd1 vccd1 vccd1 _15815_/D sky130_fd_sc_hd__and2_1
XFILLER_0_0_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08298_ hold2956/X _08336_/A2 _08297_/X _13684_/C1 vssd1 vssd1 vccd1 vccd1 _08298_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5530 _11494_/X vssd1 vssd1 vccd1 vccd1 _16988_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10260_ _10551_/A _10260_/B vssd1 vssd1 vccd1 vccd1 _10260_/X sky130_fd_sc_hd__or2_1
Xhold5541 _16742_/Q vssd1 vssd1 vccd1 vccd1 hold5541/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5552 _10714_/X vssd1 vssd1 vccd1 vccd1 _16728_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5563 _17644_/Q vssd1 vssd1 vccd1 vccd1 hold5563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5574 _13783_/X vssd1 vssd1 vccd1 vccd1 _17714_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4840 _09736_/X vssd1 vssd1 vccd1 vccd1 _16402_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5585 _16961_/Q vssd1 vssd1 vccd1 vccd1 hold5585/X sky130_fd_sc_hd__dlygate4sd3_1
X_10191_ _11091_/A _10191_/B vssd1 vssd1 vccd1 vccd1 _10191_/X sky130_fd_sc_hd__or2_1
Xhold5596 _13498_/X vssd1 vssd1 vccd1 vccd1 _17619_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4851 _17192_/Q vssd1 vssd1 vccd1 vccd1 hold4851/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4862 _11041_/X vssd1 vssd1 vccd1 vccd1 _16837_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4873 _17158_/Q vssd1 vssd1 vccd1 vccd1 hold4873/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4884 _11380_/X vssd1 vssd1 vccd1 vccd1 _16950_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4895 _17026_/Q vssd1 vssd1 vccd1 vccd1 hold4895/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout340 _12441_/S vssd1 vssd1 vccd1 vccd1 _12443_/S sky130_fd_sc_hd__buf_8
XFILLER_0_79_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout351 _08910_/S vssd1 vssd1 vccd1 vccd1 _08930_/S sky130_fd_sc_hd__buf_8
XFILLER_0_121_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout362 _15507_/Y vssd1 vssd1 vccd1 vccd1 _15560_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout373 _15020_/X vssd1 vssd1 vccd1 vccd1 _15069_/S sky130_fd_sc_hd__clkbuf_8
X_13950_ _14166_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13950_/X sky130_fd_sc_hd__or2_1
XFILLER_0_219_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout384 _14788_/Y vssd1 vssd1 vccd1 vccd1 _14828_/B sky130_fd_sc_hd__buf_8
XFILLER_0_156_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout395 _14543_/B vssd1 vssd1 vccd1 vccd1 _14553_/B sky130_fd_sc_hd__buf_8
X_12901_ hold2479/X hold3141/X _12916_/S vssd1 vssd1 vccd1 vccd1 _12901_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_236_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13881_ hold4514/X _13791_/A _13880_/X vssd1 vssd1 vccd1 vccd1 _13881_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15620_ _17153_/CLK _15620_/D vssd1 vssd1 vccd1 vccd1 _15620_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12832_ hold1929/X _17455_/Q _12838_/S vssd1 vssd1 vccd1 vccd1 _12832_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ hold992/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15551_/X sky130_fd_sc_hd__or2_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12763_ hold973/X _17432_/Q _12766_/S vssd1 vssd1 vccd1 vccd1 _12763_/X sky130_fd_sc_hd__mux2_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _15182_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14543_/B sky130_fd_sc_hd__or2_4
X_18270_ _18423_/CLK _18270_/D vssd1 vssd1 vccd1 vccd1 _18270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11714_ hold1525/X _17062_/Q _12305_/C vssd1 vssd1 vccd1 vccd1 _11715_/B sky130_fd_sc_hd__mux2_1
X_15482_ _15482_/A _15482_/B vssd1 vssd1 vccd1 vccd1 _18424_/D sky130_fd_sc_hd__and2_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ hold1269/X hold3964/X _12838_/S vssd1 vssd1 vccd1 vccd1 _12694_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17221_ _17221_/CLK _17221_/D vssd1 vssd1 vccd1 vccd1 _17221_/Q sky130_fd_sc_hd__dfxtp_1
X_14433_ _15547_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _14433_/Y sky130_fd_sc_hd__nand2_1
X_11645_ hold1962/X hold4087/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11646_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_182_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17152_ _17280_/CLK _17152_/D vssd1 vssd1 vccd1 vccd1 _17152_/Q sky130_fd_sc_hd__dfxtp_1
Xinput15 input15/A vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14364_ _14364_/A _14364_/B vssd1 vssd1 vccd1 vccd1 _17981_/D sky130_fd_sc_hd__and2_1
Xinput26 input26/A vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_6
X_11576_ hold2530/X hold4875/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11577_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_13_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput37 input37/A vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__buf_1
XFILLER_0_107_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16103_ _17325_/CLK _16103_/D vssd1 vssd1 vccd1 vccd1 _16103_/Q sky130_fd_sc_hd__dfxtp_1
Xinput48 input48/A vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput59 input59/A vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__buf_6
X_13315_ hold4681/X _12353_/B _13314_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _13315_/X
+ sky130_fd_sc_hd__o211a_1
X_10527_ _10554_/A _10527_/B vssd1 vssd1 vccd1 vccd1 _10527_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17083_ _17771_/CLK _17083_/D vssd1 vssd1 vccd1 vccd1 _17083_/Q sky130_fd_sc_hd__dfxtp_1
X_14295_ hold2175/X _14333_/A2 _14294_/X _14364_/A vssd1 vssd1 vccd1 vccd1 _14295_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16034_ _17309_/CLK _16034_/D vssd1 vssd1 vccd1 vccd1 hold379/A sky130_fd_sc_hd__dfxtp_1
X_13246_ _13246_/A _13294_/B vssd1 vssd1 vccd1 vccd1 _13246_/X sky130_fd_sc_hd__or2_1
X_10458_ _10554_/A _10458_/B vssd1 vssd1 vccd1 vccd1 _10458_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_454_wb_clk_i clkbuf_6_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17661_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_209_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13177_ _13177_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13177_/X sky130_fd_sc_hd__and2_1
XFILLER_0_202_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10389_ _10530_/A _10389_/B vssd1 vssd1 vccd1 vccd1 _10389_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_236_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12128_ hold1604/X hold4791/X _13409_/S vssd1 vssd1 vccd1 vccd1 _12129_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17985_ _17985_/CLK _17985_/D vssd1 vssd1 vccd1 vccd1 _17985_/Q sky130_fd_sc_hd__dfxtp_1
X_12059_ hold1336/X _17177_/Q _13463_/S vssd1 vssd1 vccd1 vccd1 _12060_/B sky130_fd_sc_hd__mux2_1
X_16936_ _18429_/CLK _16936_/D vssd1 vssd1 vccd1 vccd1 _16936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_236_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16867_ _18070_/CLK _16867_/D vssd1 vssd1 vccd1 vccd1 _16867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15818_ _17729_/CLK hold231/X vssd1 vssd1 vccd1 vccd1 _15818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16798_ _18053_/CLK _16798_/D vssd1 vssd1 vccd1 vccd1 _16798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15749_ _17718_/CLK _15749_/D vssd1 vssd1 vccd1 vccd1 _15749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09270_ _09272_/A hold365/X vssd1 vssd1 vccd1 vccd1 _16246_/D sky130_fd_sc_hd__and2_1
XFILLER_0_111_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08221_ _15555_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08221_/X sky130_fd_sc_hd__or2_1
X_17419_ _17427_/CLK _17419_/D vssd1 vssd1 vccd1 vccd1 _17419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18399_ _18399_/CLK _18399_/D vssd1 vssd1 vccd1 vccd1 _18399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08152_ _15557_/A hold1112/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08153_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08083_ hold3047/X _08088_/B _08082_/Y _13943_/A vssd1 vssd1 vccd1 vccd1 _08083_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4103 _16893_/Q vssd1 vssd1 vccd1 vccd1 _11207_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4114 _11101_/X vssd1 vssd1 vccd1 vccd1 _16857_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_195_wb_clk_i clkbuf_6_53_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18324_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4125 _17650_/Q vssd1 vssd1 vccd1 vccd1 hold4125/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4136 _10717_/X vssd1 vssd1 vccd1 vccd1 _16729_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3402 hold5949/X vssd1 vssd1 vccd1 vccd1 hold5950/A sky130_fd_sc_hd__buf_6
XFILLER_0_144_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4147 _16830_/Q vssd1 vssd1 vccd1 vccd1 hold4147/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3413 _10003_/Y vssd1 vssd1 vccd1 vccd1 _16491_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_124_wb_clk_i clkbuf_6_22_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17337_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4158 _16476_/Q vssd1 vssd1 vccd1 vccd1 hold4158/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3424 _10578_/Y vssd1 vssd1 vccd1 vccd1 _10579_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4169 _16438_/Q vssd1 vssd1 vccd1 vccd1 hold4169/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3435 _16524_/Q vssd1 vssd1 vccd1 vccd1 hold3435/X sky130_fd_sc_hd__buf_2
XFILLER_0_227_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3446 _09997_/Y vssd1 vssd1 vccd1 vccd1 _16489_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2701 _17956_/Q vssd1 vssd1 vccd1 vccd1 hold2701/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3457 _10005_/Y vssd1 vssd1 vccd1 vccd1 _10006_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2712 _14009_/X vssd1 vssd1 vccd1 vccd1 _17810_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08985_ hold438/X hold569/X _08991_/S vssd1 vssd1 vccd1 vccd1 _08986_/B sky130_fd_sc_hd__mux2_1
Xhold2723 _18116_/Q vssd1 vssd1 vccd1 vccd1 hold2723/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3468 _16528_/Q vssd1 vssd1 vccd1 vccd1 hold3468/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_139_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3479 _16716_/Q vssd1 vssd1 vccd1 vccd1 hold3479/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2734 _08182_/X vssd1 vssd1 vccd1 vccd1 _15727_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2745 _18445_/Q vssd1 vssd1 vccd1 vccd1 hold2745/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07936_ _15559_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07936_/X sky130_fd_sc_hd__or2_1
Xhold2756 _18455_/Q vssd1 vssd1 vccd1 vccd1 hold2756/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2767 _16264_/Q vssd1 vssd1 vccd1 vccd1 hold2767/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2778 _14281_/X vssd1 vssd1 vccd1 vccd1 _17941_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2789 _13961_/X vssd1 vssd1 vccd1 vccd1 _17787_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07867_ _15545_/A _07869_/B vssd1 vssd1 vccd1 vccd1 _07867_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09606_ _09984_/A _09606_/B vssd1 vssd1 vccd1 vccd1 _09606_/X sky130_fd_sc_hd__or2_1
XFILLER_0_195_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07798_ _07804_/A _09342_/A _09339_/B hold3129/X vssd1 vssd1 vccd1 vccd1 _07798_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09537_ _09981_/A _09537_/B vssd1 vssd1 vccd1 vccd1 _09537_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09468_ _09472_/C _09472_/D hold739/X vssd1 vssd1 vccd1 vccd1 _09468_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_94_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08419_ _15207_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08419_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09399_ _15559_/A _14555_/C _09399_/C _09398_/X vssd1 vssd1 vccd1 vccd1 _09400_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_0_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11430_ _12210_/A _11430_/B vssd1 vssd1 vccd1 vccd1 _11430_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11361_ _11553_/A _11361_/B vssd1 vssd1 vccd1 vccd1 _11361_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6050 _16202_/Q vssd1 vssd1 vccd1 vccd1 hold6050/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6061 _18346_/Q vssd1 vssd1 vccd1 vccd1 hold6061/X sky130_fd_sc_hd__dlygate4sd3_1
X_10312_ hold4501/X _10628_/B _10311_/X _14895_/C1 vssd1 vssd1 vccd1 vccd1 _10312_/X
+ sky130_fd_sc_hd__o211a_1
X_13100_ hold4328/X _13099_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13100_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_15_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11292_ _12243_/A _11292_/B vssd1 vssd1 vccd1 vccd1 _11292_/X sky130_fd_sc_hd__or2_1
X_14080_ _15533_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14080_/X sky130_fd_sc_hd__or2_1
Xhold6072 _17884_/Q vssd1 vssd1 vccd1 vccd1 hold6072/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6083 data_in[0] vssd1 vssd1 vccd1 vccd1 hold223/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6094 la_data_in[21] vssd1 vssd1 vccd1 vccd1 hold988/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5360 _11341_/X vssd1 vssd1 vccd1 vccd1 _16937_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13031_ hold896/X hold905/X hold936/X vssd1 vssd1 vccd1 vccd1 _17520_/D sky130_fd_sc_hd__and3b_1
X_10243_ hold3712/X _10625_/B _10242_/X _14893_/C1 vssd1 vssd1 vccd1 vccd1 _10243_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5371 _11365_/X vssd1 vssd1 vccd1 vccd1 _16945_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5382 _17070_/Q vssd1 vssd1 vccd1 vccd1 hold5382/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5393 _11692_/X vssd1 vssd1 vccd1 vccd1 _17054_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4670 _17125_/Q vssd1 vssd1 vccd1 vccd1 hold4670/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10174_ hold3654/X _11186_/B _10173_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10174_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4681 _17590_/Q vssd1 vssd1 vccd1 vccd1 hold4681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4692 _09625_/X vssd1 vssd1 vccd1 vccd1 _16365_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3980 _16853_/Q vssd1 vssd1 vccd1 vccd1 hold3980/X sky130_fd_sc_hd__dlygate4sd3_1
X_17770_ _17832_/CLK _17770_/D vssd1 vssd1 vccd1 vccd1 _17770_/Q sky130_fd_sc_hd__dfxtp_1
X_14982_ hold933/X hold510/A vssd1 vssd1 vccd1 vccd1 _14982_/X sky130_fd_sc_hd__or2_1
Xhold3991 _16876_/Q vssd1 vssd1 vccd1 vccd1 hold3991/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout170 _12217_/A2 vssd1 vssd1 vccd1 vccd1 _12356_/B sky130_fd_sc_hd__buf_4
Xfanout181 _11071_/A2 vssd1 vssd1 vccd1 vccd1 _11744_/B sky130_fd_sc_hd__buf_4
X_16721_ _18052_/CLK _16721_/D vssd1 vssd1 vccd1 vccd1 _16721_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout192 _13877_/B vssd1 vssd1 vccd1 vccd1 _13874_/B sky130_fd_sc_hd__clkbuf_4
X_13933_ _13933_/A hold298/X vssd1 vssd1 vccd1 vccd1 hold299/A sky130_fd_sc_hd__and2_1
XFILLER_0_199_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16652_ _18146_/CLK _16652_/D vssd1 vssd1 vccd1 vccd1 _16652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13864_ _13864_/A _13864_/B vssd1 vssd1 vccd1 vccd1 _13864_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_187_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15603_ _17280_/CLK _15603_/D vssd1 vssd1 vccd1 vccd1 _15603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12815_ hold3937/X _12814_/X _12839_/S vssd1 vssd1 vccd1 vccd1 _12816_/B sky130_fd_sc_hd__mux2_1
X_16583_ _18115_/CLK _16583_/D vssd1 vssd1 vccd1 vccd1 _16583_/Q sky130_fd_sc_hd__dfxtp_1
X_13795_ hold4676/X _13795_/A2 _13794_/X _13795_/C1 vssd1 vssd1 vccd1 vccd1 _17718_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18322_ _18342_/CLK _18322_/D vssd1 vssd1 vccd1 vccd1 _18322_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ hold2745/X _15547_/B _15533_/X _12822_/A vssd1 vssd1 vccd1 vccd1 _15534_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12746_ hold3178/X _12745_/X _12749_/S vssd1 vssd1 vccd1 vccd1 _12746_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18253_ _18357_/CLK _18253_/D vssd1 vssd1 vccd1 vccd1 _18253_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15465_ _15465_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15465_/X sky130_fd_sc_hd__or2_1
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12677_ hold3154/X _12676_/X _12851_/S vssd1 vssd1 vccd1 vccd1 _12677_/X sky130_fd_sc_hd__mux2_1
X_17204_ _17204_/CLK _17204_/D vssd1 vssd1 vccd1 vccd1 _17204_/Q sky130_fd_sc_hd__dfxtp_1
X_14416_ hold2805/X _14446_/A2 _14415_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _14416_/X
+ sky130_fd_sc_hd__o211a_1
X_18184_ _18226_/CLK _18184_/D vssd1 vssd1 vccd1 vccd1 _18184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11628_ _11631_/A _11628_/B vssd1 vssd1 vccd1 vccd1 _11628_/X sky130_fd_sc_hd__or2_1
X_15396_ _17343_/Q _15486_/B1 _15485_/B1 hold835/X vssd1 vssd1 vccd1 vccd1 _15396_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17135_ _17771_/CLK _17135_/D vssd1 vssd1 vccd1 vccd1 _17135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14347_ _15189_/A hold3191/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14348_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_53_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11559_ _11658_/A _11559_/B vssd1 vssd1 vccd1 vccd1 _11559_/X sky130_fd_sc_hd__or2_1
Xhold607 hold607/A vssd1 vssd1 vccd1 vccd1 hold607/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 hold618/A vssd1 vssd1 vccd1 vccd1 hold618/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold629 input42/X vssd1 vssd1 vccd1 vccd1 hold629/X sky130_fd_sc_hd__clkbuf_2
X_17066_ _17850_/CLK _17066_/D vssd1 vssd1 vccd1 vccd1 _17066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14278_ _14726_/A _14282_/B vssd1 vssd1 vccd1 vccd1 _14278_/X sky130_fd_sc_hd__or2_1
XFILLER_0_111_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16017_ _18240_/CLK _16017_/D vssd1 vssd1 vccd1 vccd1 hold602/A sky130_fd_sc_hd__dfxtp_1
X_13229_ _13228_/X hold3200/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13229_/X sky130_fd_sc_hd__mux2_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2008 _17970_/Q vssd1 vssd1 vccd1 vccd1 hold2008/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2019 _18122_/Q vssd1 vssd1 vccd1 vccd1 hold2019/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1307 _15735_/Q vssd1 vssd1 vccd1 vccd1 hold1307/X sky130_fd_sc_hd__dlygate4sd3_1
X_08770_ _15364_/A _08770_/B vssd1 vssd1 vccd1 vccd1 _16005_/D sky130_fd_sc_hd__and2_1
Xhold1318 _08073_/X vssd1 vssd1 vccd1 vccd1 _15676_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17968_ _17968_/CLK _17968_/D vssd1 vssd1 vccd1 vccd1 _17968_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1329 _15711_/Q vssd1 vssd1 vccd1 vccd1 hold1329/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16919_ _18069_/CLK _16919_/D vssd1 vssd1 vccd1 vccd1 _16919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17899_ _17899_/CLK _17899_/D vssd1 vssd1 vccd1 vccd1 _17899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09322_ hold2944/X _09323_/B _09321_/Y _12588_/A vssd1 vssd1 vccd1 vccd1 _09322_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09253_ _15529_/A hold2552/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09254_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08204_ hold1397/X _08209_/B _08203_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _08204_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09184_ _15513_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09184_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_376_wb_clk_i clkbuf_6_32_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17678_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08135_ _08135_/A _08135_/B vssd1 vssd1 vccd1 vccd1 _15706_/D sky130_fd_sc_hd__and2_1
XFILLER_0_181_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_305_wb_clk_i clkbuf_6_44_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17874_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08066_ _15525_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08066_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3210 _17445_/Q vssd1 vssd1 vccd1 vccd1 hold3210/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3221 _12572_/X vssd1 vssd1 vccd1 vccd1 _12573_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3232 _17497_/Q vssd1 vssd1 vccd1 vccd1 hold3232/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3243 _16677_/Q vssd1 vssd1 vccd1 vccd1 hold3243/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3254 _10471_/X vssd1 vssd1 vccd1 vccd1 _16647_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2520 _17851_/Q vssd1 vssd1 vccd1 vccd1 hold2520/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3265 _17378_/Q vssd1 vssd1 vccd1 vccd1 hold3265/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3276 _16439_/Q vssd1 vssd1 vccd1 vccd1 hold3276/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2531 _14121_/X vssd1 vssd1 vccd1 vccd1 _17864_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2542 _15850_/Q vssd1 vssd1 vccd1 vccd1 hold2542/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3287 _12602_/X vssd1 vssd1 vccd1 vccd1 _12603_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08968_ _15491_/A hold738/X vssd1 vssd1 vccd1 vccd1 _16101_/D sky130_fd_sc_hd__and2_1
XFILLER_0_216_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3298 _16663_/Q vssd1 vssd1 vccd1 vccd1 hold3298/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2553 _17877_/Q vssd1 vssd1 vccd1 vccd1 hold2553/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2564 _16230_/Q vssd1 vssd1 vccd1 vccd1 hold2564/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1830 _14893_/X vssd1 vssd1 vccd1 vccd1 _18235_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2575 _15876_/Q vssd1 vssd1 vccd1 vccd1 hold2575/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2586 _14619_/X vssd1 vssd1 vccd1 vccd1 _18103_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1841 _15789_/Q vssd1 vssd1 vccd1 vccd1 hold1841/X sky130_fd_sc_hd__dlygate4sd3_1
X_07919_ hold2792/X _07918_/B _07918_/Y _08153_/A vssd1 vssd1 vccd1 vccd1 _07919_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1852 _14311_/X vssd1 vssd1 vccd1 vccd1 _17955_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2597 _17811_/Q vssd1 vssd1 vccd1 vccd1 hold2597/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1863 _18227_/Q vssd1 vssd1 vccd1 vccd1 hold1863/X sky130_fd_sc_hd__dlygate4sd3_1
X_08899_ _12418_/A _08899_/B vssd1 vssd1 vccd1 vccd1 _16067_/D sky130_fd_sc_hd__and2_1
XFILLER_0_230_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_230_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1874 _14077_/X vssd1 vssd1 vccd1 vccd1 _17843_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1885 _18062_/Q vssd1 vssd1 vccd1 vccd1 hold1885/X sky130_fd_sc_hd__dlygate4sd3_1
X_10930_ hold5064/X _11225_/B _10929_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _10930_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_1322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1896 _09417_/X vssd1 vssd1 vccd1 vccd1 _16294_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_92_wb_clk_i clkbuf_6_17_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16315_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10861_ hold4053/X _11144_/B _10860_/X _14354_/A vssd1 vssd1 vccd1 vccd1 _16777_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_21_wb_clk_i clkbuf_6_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17477_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_190_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _12612_/A _12600_/B vssd1 vssd1 vccd1 vccd1 _17376_/D sky130_fd_sc_hd__and2_1
XFILLER_0_183_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13580_ hold2341/X _17647_/Q _13868_/C vssd1 vssd1 vccd1 vccd1 _13581_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10792_ hold4059/X _11210_/B _10791_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _10792_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _12984_/A _12531_/B vssd1 vssd1 vccd1 vccd1 _17353_/D sky130_fd_sc_hd__and2_1
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ hold639/X _15448_/A2 _15446_/B1 hold797/X vssd1 vssd1 vccd1 vccd1 _15250_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12462_ _17324_/Q _12506_/B vssd1 vssd1 vccd1 vccd1 _12462_/X sky130_fd_sc_hd__or2_1
XFILLER_0_152_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14201_ hold2609/X _14202_/B _14200_/Y _14348_/A vssd1 vssd1 vccd1 vccd1 _14201_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11413_ hold4089/X _11792_/B _11412_/X _14143_/C1 vssd1 vssd1 vccd1 vccd1 _11413_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15181_ _15182_/A _15182_/B vssd1 vssd1 vccd1 vccd1 _15181_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12393_ hold29/X hold274/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12394_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14132_ hold520/X _14160_/B vssd1 vssd1 vccd1 vccd1 hold521/A sky130_fd_sc_hd__or2_1
XFILLER_0_105_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11344_ hold5517/X _11726_/B _11343_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _11344_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14063_ hold2884/X _14094_/B _14062_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _14063_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11275_ hold5645/X _11753_/B _11274_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11275_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5190 _11575_/X vssd1 vssd1 vccd1 vccd1 _17015_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13014_ hold6058/X _13003_/Y hold946/X _12984_/A vssd1 vssd1 vccd1 vccd1 hold947/A
+ sky130_fd_sc_hd__o211a_1
X_10226_ hold2295/X hold4436/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10227_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_219_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10157_ hold1764/X _16543_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10158_/B sky130_fd_sc_hd__mux2_1
X_17822_ _17825_/CLK _17822_/D vssd1 vssd1 vccd1 vccd1 _17822_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_234_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_234_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10088_ hold2231/X hold3428/X _10571_/C vssd1 vssd1 vccd1 vccd1 _10089_/B sky130_fd_sc_hd__mux2_1
X_14965_ hold2075/X _14952_/B _14964_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _14965_/X
+ sky130_fd_sc_hd__o211a_1
X_17753_ _17753_/CLK input71/X vssd1 vssd1 vccd1 vccd1 _17753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_238_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16704_ _18224_/CLK _16704_/D vssd1 vssd1 vccd1 vccd1 _16704_/Q sky130_fd_sc_hd__dfxtp_1
X_13916_ _14596_/A hold1196/X hold297/X vssd1 vssd1 vccd1 vccd1 _13916_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_96_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17684_ _17716_/CLK _17684_/D vssd1 vssd1 vccd1 vccd1 _17684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14896_ _14897_/A _15182_/B vssd1 vssd1 vccd1 vccd1 _14896_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16635_ _18225_/CLK _16635_/D vssd1 vssd1 vccd1 vccd1 _16635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13847_ _17736_/Q _13847_/B _13868_/C vssd1 vssd1 vccd1 vccd1 _13847_/X sky130_fd_sc_hd__and3_1
XFILLER_0_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16566_ _18156_/CLK _16566_/D vssd1 vssd1 vccd1 vccd1 _16566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13778_ hold1425/X _17713_/Q _13874_/C vssd1 vssd1 vccd1 vccd1 _13779_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_146_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18305_ _18416_/CLK _18305_/D vssd1 vssd1 vccd1 vccd1 _18305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15517_ _15517_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15517_/X sky130_fd_sc_hd__or2_1
XFILLER_0_139_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12729_ _12753_/A _12729_/B vssd1 vssd1 vccd1 vccd1 _17419_/D sky130_fd_sc_hd__and2_1
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16497_ _18378_/CLK _16497_/D vssd1 vssd1 vccd1 vccd1 _16497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18236_ _18236_/CLK _18236_/D vssd1 vssd1 vccd1 vccd1 _18236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15448_ _15930_/Q _15448_/A2 _15486_/B1 hold310/X vssd1 vssd1 vccd1 vccd1 _15448_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_217_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18167_ _18232_/CLK _18167_/D vssd1 vssd1 vccd1 vccd1 _18167_/Q sky130_fd_sc_hd__dfxtp_1
X_15379_ hold812/X _09365_/B _15488_/A2 hold633/X _15378_/X vssd1 vssd1 vccd1 vccd1
+ _15382_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_68_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold404 input56/X vssd1 vssd1 vccd1 vccd1 hold404/X sky130_fd_sc_hd__dlygate4sd3_1
X_17118_ _17278_/CLK _17118_/D vssd1 vssd1 vccd1 vccd1 _17118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold415 hold415/A vssd1 vssd1 vccd1 vccd1 hold415/X sky130_fd_sc_hd__dlygate4sd3_1
X_18098_ _18162_/CLK _18098_/D vssd1 vssd1 vccd1 vccd1 _18098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold426 hold426/A vssd1 vssd1 vccd1 vccd1 hold426/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 input22/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__buf_1
Xhold448 hold448/A vssd1 vssd1 vccd1 vccd1 hold448/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 hold459/A vssd1 vssd1 vccd1 vccd1 hold459/X sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ hold5833/X _10022_/B _09939_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09940_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17049_ _17865_/CLK _17049_/D vssd1 vssd1 vccd1 vccd1 _17049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout906 hold579/X vssd1 vssd1 vccd1 vccd1 _15233_/A sky130_fd_sc_hd__buf_4
XFILLER_0_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09871_ hold3628/X _10049_/B _09870_/X _15212_/C1 vssd1 vssd1 vccd1 vccd1 _09871_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout917 hold991/X vssd1 vssd1 vccd1 vccd1 hold992/A sky130_fd_sc_hd__clkbuf_16
Xfanout928 hold1253/X vssd1 vssd1 vccd1 vccd1 _14604_/A sky130_fd_sc_hd__buf_8
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout939 hold1007/X vssd1 vssd1 vccd1 vccd1 hold1008/A sky130_fd_sc_hd__buf_4
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08822_ hold673/X hold830/X _08860_/S vssd1 vssd1 vccd1 vccd1 hold831/A sky130_fd_sc_hd__mux2_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 _07991_/X vssd1 vssd1 vccd1 vccd1 _15638_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1115 _15757_/Q vssd1 vssd1 vccd1 vccd1 hold1115/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 _08406_/X vssd1 vssd1 vccd1 vccd1 _15833_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 hold1224/X vssd1 vssd1 vccd1 vccd1 hold1137/X sky130_fd_sc_hd__buf_1
X_08753_ hold163/X hold479/X _08779_/S vssd1 vssd1 vccd1 vccd1 hold480/A sky130_fd_sc_hd__mux2_1
Xhold1148 _15154_/X vssd1 vssd1 vccd1 vccd1 _18360_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 _17969_/Q vssd1 vssd1 vccd1 vccd1 hold1159/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ _12418_/A hold857/X vssd1 vssd1 vccd1 vccd1 _15963_/D sky130_fd_sc_hd__and2_1
XFILLER_0_205_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09305_ hold951/X _09315_/B vssd1 vssd1 vccd1 vccd1 _09305_/X sky130_fd_sc_hd__or2_1
XFILLER_0_118_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09236_ _12843_/A _09236_/B vssd1 vssd1 vccd1 vccd1 _16229_/D sky130_fd_sc_hd__and2_1
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09167_ hold1641/X _09177_/A2 _09166_/X _12906_/A vssd1 vssd1 vccd1 vccd1 _09167_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08118_ _14517_/A hold941/X _08152_/S vssd1 vssd1 vccd1 vccd1 hold942/A sky130_fd_sc_hd__mux2_1
XFILLER_0_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09098_ _15539_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _09098_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08049_ hold355/X _14627_/A vssd1 vssd1 vccd1 vccd1 _08100_/B sky130_fd_sc_hd__or2_4
Xhold960 hold960/A vssd1 vssd1 vccd1 vccd1 hold960/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 hold971/A vssd1 vssd1 vccd1 vccd1 hold971/X sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ hold636/X hold3310/X _11144_/C vssd1 vssd1 vccd1 vccd1 _11061_/B sky130_fd_sc_hd__mux2_1
Xhold982 hold982/A vssd1 vssd1 vccd1 vccd1 hold982/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 hold993/A vssd1 vssd1 vccd1 vccd1 hold993/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3040 _14143_/X vssd1 vssd1 vccd1 vccd1 _17875_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10011_ _13142_/A _09981_/A _10010_/X vssd1 vssd1 vccd1 vccd1 _10011_/Y sky130_fd_sc_hd__a21oi_1
Xhold3051 _18293_/Q vssd1 vssd1 vccd1 vccd1 hold3051/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3062 _14177_/X vssd1 vssd1 vccd1 vccd1 _17891_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3073 _14987_/X vssd1 vssd1 vccd1 vccd1 _18279_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3084 hold5895/X vssd1 vssd1 vccd1 vccd1 _09339_/A sky130_fd_sc_hd__clkbuf_4
XTAP_5246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2350 _15192_/X vssd1 vssd1 vccd1 vccd1 _18378_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3095 _15621_/Q vssd1 vssd1 vccd1 vccd1 hold3095/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2361 _16258_/Q vssd1 vssd1 vccd1 vccd1 hold2361/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2372 _09135_/X vssd1 vssd1 vccd1 vccd1 _16180_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2383 _09077_/X vssd1 vssd1 vccd1 vccd1 _16153_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2394 _15873_/Q vssd1 vssd1 vccd1 vccd1 hold2394/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1660 _17828_/Q vssd1 vssd1 vccd1 vccd1 hold1660/X sky130_fd_sc_hd__dlygate4sd3_1
X_14750_ _15197_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14750_/X sky130_fd_sc_hd__or2_1
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1671 _14257_/X vssd1 vssd1 vccd1 vccd1 _17929_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1682 _17946_/Q vssd1 vssd1 vccd1 vccd1 hold1682/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11962_ hold5179/X _12374_/B _11961_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _11962_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1693 _14787_/X vssd1 vssd1 vccd1 vccd1 _18184_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _13800_/A _13701_/B vssd1 vssd1 vccd1 vccd1 _13701_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10913_ hold2013/X hold5072/X _11171_/C vssd1 vssd1 vccd1 vccd1 _10914_/B sky130_fd_sc_hd__mux2_1
X_14681_ _14681_/A _14843_/B vssd1 vssd1 vccd1 vccd1 _14730_/B sky130_fd_sc_hd__or2_4
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ hold4072/X _13886_/B _11892_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _11893_/X
+ sky130_fd_sc_hd__o211a_1
X_16420_ _18379_/CLK _16420_/D vssd1 vssd1 vccd1 vccd1 _16420_/Q sky130_fd_sc_hd__dfxtp_1
X_13632_ _13737_/A _13632_/B vssd1 vssd1 vccd1 vccd1 _13632_/X sky130_fd_sc_hd__or2_1
X_10844_ _17975_/Q hold4085/X _11738_/C vssd1 vssd1 vccd1 vccd1 _10845_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_184_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_298_wb_clk_i clkbuf_6_39_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17892_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16351_ _18296_/CLK _16351_/D vssd1 vssd1 vccd1 vccd1 _16351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13563_ _13791_/A _13563_/B vssd1 vssd1 vccd1 vccd1 _13563_/X sky130_fd_sc_hd__or2_1
X_10775_ hold3112/X hold4668/X _11162_/C vssd1 vssd1 vccd1 vccd1 _10776_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_227_wb_clk_i clkbuf_6_63_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18221_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15302_ _15489_/A _15302_/B _15302_/C _15302_/D vssd1 vssd1 vccd1 vccd1 _15302_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_66_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12514_ hold1528/X hold4477/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12514_/X sky130_fd_sc_hd__mux2_1
X_16282_ _17750_/CLK _16282_/D vssd1 vssd1 vccd1 vccd1 _16282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13494_ _13599_/A _13494_/B vssd1 vssd1 vccd1 vccd1 _13494_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18021_ _18021_/CLK _18021_/D vssd1 vssd1 vccd1 vccd1 _18021_/Q sky130_fd_sc_hd__dfxtp_1
X_15233_ _15233_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15233_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12445_ _12445_/A _12445_/B vssd1 vssd1 vccd1 vccd1 _12508_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_23_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15164_ hold2422/X _15167_/B _15163_/Y _15202_/C1 vssd1 vssd1 vccd1 vccd1 _15164_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12376_ _13888_/A _12376_/B vssd1 vssd1 vccd1 vccd1 _12376_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_105_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_238_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14115_ hold1849/X _14142_/B _14114_/X _14346_/A vssd1 vssd1 vccd1 vccd1 _14115_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11327_ hold2039/X hold4091/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11328_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_239_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15095_ _15203_/A _15119_/B vssd1 vssd1 vccd1 vccd1 _15095_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14046_ _14726_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14046_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11258_ hold2890/X hold4417/X _11738_/C vssd1 vssd1 vccd1 vccd1 _11259_/B sky130_fd_sc_hd__mux2_1
X_10209_ _10563_/A _10209_/B vssd1 vssd1 vccd1 vccd1 _10209_/X sky130_fd_sc_hd__or2_1
XFILLER_0_101_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11189_ _16887_/Q _11225_/B _11216_/C vssd1 vssd1 vccd1 vccd1 _11189_/X sky130_fd_sc_hd__and3_1
XFILLER_0_101_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17805_ _17891_/CLK _17805_/D vssd1 vssd1 vccd1 vccd1 _17805_/Q sky130_fd_sc_hd__dfxtp_1
X_15997_ _16093_/CLK _15997_/D vssd1 vssd1 vccd1 vccd1 hold479/A sky130_fd_sc_hd__dfxtp_1
XTAP_5780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14948_ _15217_/A _14952_/B vssd1 vssd1 vccd1 vccd1 _14948_/Y sky130_fd_sc_hd__nand2_1
X_17736_ _17740_/CLK _17736_/D vssd1 vssd1 vccd1 vccd1 _17736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14879_ hold1095/X hold332/X _14878_/Y _14895_/C1 vssd1 vssd1 vccd1 vccd1 _14879_/X
+ sky130_fd_sc_hd__o211a_1
X_17667_ _17697_/CLK _17667_/D vssd1 vssd1 vccd1 vccd1 _17667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_212_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16618_ _18208_/CLK _16618_/D vssd1 vssd1 vccd1 vccd1 _16618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17598_ _17630_/CLK _17598_/D vssd1 vssd1 vccd1 vccd1 _17598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16549_ _18262_/CLK _16549_/D vssd1 vssd1 vccd1 vccd1 _16549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09021_ _15434_/A _09021_/B vssd1 vssd1 vccd1 vccd1 _16127_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18219_ _18227_/CLK _18219_/D vssd1 vssd1 vccd1 vccd1 _18219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5904 output94/X vssd1 vssd1 vccd1 vccd1 data_out[2] sky130_fd_sc_hd__buf_12
XFILLER_0_5_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5915 _18401_/Q vssd1 vssd1 vccd1 vccd1 hold5915/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold201 hold201/A vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5926 _18403_/Q vssd1 vssd1 vccd1 vccd1 hold5926/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 hold212/A vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5937 hold5937/A vssd1 vssd1 vccd1 vccd1 hold5937/X sky130_fd_sc_hd__clkbuf_4
Xhold223 hold223/A vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5948 hold5948/A vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_12
XFILLER_0_223_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold234 input47/X vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold5959 hold5959/A vssd1 vssd1 vccd1 vccd1 hold5959/X sky130_fd_sc_hd__clkbuf_4
Xhold245 hold62/X vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__buf_4
XFILLER_0_106_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold256 hold256/A vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold267 hold352/X vssd1 vssd1 vccd1 vccd1 hold353/A sky130_fd_sc_hd__buf_4
Xhold278 hold68/X vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__clkbuf_8
Xclkbuf_6_48_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_48_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_09923_ hold2349/X _16465_/Q _10475_/S vssd1 vssd1 vccd1 vccd1 _09924_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_229_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout703 _09047_/A vssd1 vssd1 vccd1 vccd1 _15254_/A sky130_fd_sc_hd__buf_2
Xhold289 hold289/A vssd1 vssd1 vccd1 vccd1 hold289/X sky130_fd_sc_hd__buf_12
Xfanout714 fanout739/X vssd1 vssd1 vccd1 vccd1 _15491_/A sky130_fd_sc_hd__buf_4
XFILLER_0_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout725 _09907_/C1 vssd1 vssd1 vccd1 vccd1 _15176_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_238_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout736 _15473_/A vssd1 vssd1 vccd1 vccd1 _15062_/A sky130_fd_sc_hd__buf_4
XFILLER_0_141_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09854_ hold984/X _16442_/Q _10067_/C vssd1 vssd1 vccd1 vccd1 _09855_/B sky130_fd_sc_hd__mux2_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout747 _13777_/C1 vssd1 vssd1 vccd1 vccd1 _08381_/A sky130_fd_sc_hd__buf_4
XFILLER_0_42_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout758 _14131_/C1 vssd1 vssd1 vccd1 vccd1 _14380_/A sky130_fd_sc_hd__buf_4
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout769 _08131_/A vssd1 vssd1 vccd1 vccd1 _08135_/A sky130_fd_sc_hd__buf_4
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _15374_/A hold311/X vssd1 vssd1 vccd1 vccd1 _16021_/D sky130_fd_sc_hd__and2_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ hold1213/X hold3584/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09786_/B sky130_fd_sc_hd__mux2_1
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ _15434_/A hold132/X vssd1 vssd1 vccd1 vccd1 _15988_/D sky130_fd_sc_hd__and2_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 _11203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 hold915/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ hold618/X hold791/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold792/A sky130_fd_sc_hd__mux2_1
XANTENNA_129 _15173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_240_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08598_ _12380_/A _12445_/A vssd1 vssd1 vccd1 vccd1 _08623_/S sky130_fd_sc_hd__or2_2
XFILLER_0_7_1365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_391_wb_clk_i clkbuf_6_38_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17901_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_37_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_320_wb_clk_i clkbuf_6_47_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17831_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_64_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10560_ _10560_/A _10560_/B vssd1 vssd1 vccd1 vccd1 _10560_/X sky130_fd_sc_hd__or2_1
XFILLER_0_119_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09219_ hold2557/X _09218_/B _09218_/Y _12837_/A vssd1 vssd1 vccd1 vccd1 _09219_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10491_ _10554_/A _10491_/B vssd1 vssd1 vccd1 vccd1 _10491_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12230_ hold1025/X _17234_/Q _13481_/S vssd1 vssd1 vccd1 vccd1 _12231_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_224_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12161_ hold3074/X hold4815/X _13409_/S vssd1 vssd1 vccd1 vccd1 _12162_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_31_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11112_ _11127_/A _11112_/B vssd1 vssd1 vccd1 vccd1 _11112_/X sky130_fd_sc_hd__or2_1
X_12092_ hold1382/X _17188_/Q _12305_/C vssd1 vssd1 vccd1 vccd1 _12093_/B sky130_fd_sc_hd__mux2_1
Xhold790 hold790/A vssd1 vssd1 vccd1 vccd1 hold790/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15920_ _17299_/CLK _15920_/D vssd1 vssd1 vccd1 vccd1 hold872/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11043_ _11043_/A _11043_/B vssd1 vssd1 vccd1 vccd1 _11043_/X sky130_fd_sc_hd__or2_1
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15851_ _17614_/CLK _15851_/D vssd1 vssd1 vccd1 vccd1 _15851_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2180 _15538_/X vssd1 vssd1 vccd1 vccd1 _18447_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14802_ _15195_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14802_/X sky130_fd_sc_hd__or2_1
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2191 _18333_/Q vssd1 vssd1 vccd1 vccd1 hold2191/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15782_ _17745_/CLK _15782_/D vssd1 vssd1 vccd1 vccd1 _15782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12994_ hold2031/X _17509_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12994_/X sky130_fd_sc_hd__mux2_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1490 _08218_/X vssd1 vssd1 vccd1 vccd1 _15745_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17521_ _17523_/CLK hold897/X vssd1 vssd1 vccd1 vccd1 _17521_/Q sky130_fd_sc_hd__dfxtp_1
X_14733_ hold1220/X _14720_/B _14732_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14733_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11945_ hold2197/X _17139_/Q _12329_/C vssd1 vssd1 vccd1 vccd1 _11946_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_87_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_408_wb_clk_i clkbuf_6_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17823_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _17452_/CLK _17452_/D vssd1 vssd1 vccd1 vccd1 _17452_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _15165_/A _14664_/B vssd1 vssd1 vccd1 vccd1 _14664_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_170_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11876_ hold622/X hold4370/X _13481_/S vssd1 vssd1 vccd1 vccd1 _11877_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ _18342_/CLK _16403_/D vssd1 vssd1 vccd1 vccd1 _16403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13615_ hold5781/X _13808_/B _13614_/X _12738_/A vssd1 vssd1 vccd1 vccd1 _13615_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10827_ _11100_/A _10827_/B vssd1 vssd1 vccd1 vccd1 _10827_/X sky130_fd_sc_hd__or2_1
X_17383_ _18437_/CLK _17383_/D vssd1 vssd1 vccd1 vccd1 _17383_/Q sky130_fd_sc_hd__dfxtp_1
X_14595_ hold2886/X _14610_/B _14594_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _14595_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16334_ _18375_/CLK _16334_/D vssd1 vssd1 vccd1 vccd1 _16334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13546_ hold4771/X _13862_/B _13545_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _13546_/X
+ sky130_fd_sc_hd__o211a_1
X_10758_ _11049_/A _10758_/B vssd1 vssd1 vccd1 vccd1 _10758_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16265_ _17514_/CLK _16265_/D vssd1 vssd1 vccd1 vccd1 _16265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13477_ hold5563/X _13847_/B _13476_/X _13765_/C1 vssd1 vssd1 vccd1 vccd1 _13477_/X
+ sky130_fd_sc_hd__o211a_1
X_10689_ _11655_/A _10689_/B vssd1 vssd1 vccd1 vccd1 _10689_/X sky130_fd_sc_hd__or2_1
XFILLER_0_113_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15216_ hold2852/X _15219_/B _15215_/Y _15030_/A vssd1 vssd1 vccd1 vccd1 _15216_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18004_ _18069_/CLK _18004_/D vssd1 vssd1 vccd1 vccd1 _18004_/Q sky130_fd_sc_hd__dfxtp_1
X_12428_ _12438_/A hold127/X vssd1 vssd1 vccd1 vccd1 _17307_/D sky130_fd_sc_hd__and2_1
X_16196_ _17481_/CLK _16196_/D vssd1 vssd1 vccd1 vccd1 _16196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15147_ _15201_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15147_/X sky130_fd_sc_hd__or2_1
XFILLER_0_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12359_ _17277_/Q _12362_/B _12362_/C vssd1 vssd1 vccd1 vccd1 _12359_/X sky130_fd_sc_hd__and3_1
XFILLER_0_61_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3809 _10987_/X vssd1 vssd1 vccd1 vccd1 _16819_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15078_ hold1509/X hold341/X _15077_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _15078_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14029_ hold2062/X _14038_/B _14028_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _14029_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09570_ _10560_/A _09570_/B vssd1 vssd1 vccd1 vccd1 _09570_/X sky130_fd_sc_hd__or2_1
XFILLER_0_214_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08521_ _08868_/B _13056_/C _17520_/Q vssd1 vssd1 vccd1 vccd1 _08730_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_171_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17719_ _17719_/CLK _17719_/D vssd1 vssd1 vccd1 vccd1 _17719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_149_wb_clk_i clkbuf_6_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18370_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_175_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08452_ _15511_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08452_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08383_ _08387_/A _08383_/B vssd1 vssd1 vccd1 vccd1 _15823_/D sky130_fd_sc_hd__and2_1
XFILLER_0_46_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09004_ hold131/X hold175/X _09056_/S vssd1 vssd1 vccd1 vccd1 hold176/A sky130_fd_sc_hd__mux2_1
XFILLER_0_144_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5701 _17081_/Q vssd1 vssd1 vccd1 vccd1 hold5701/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5712 _12339_/Y vssd1 vssd1 vccd1 vccd1 _12340_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5723 _17563_/Q vssd1 vssd1 vccd1 vccd1 hold5723/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5734 _13465_/X vssd1 vssd1 vccd1 vccd1 _17608_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5745 _17209_/Q vssd1 vssd1 vccd1 vccd1 hold5745/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5756 _12157_/X vssd1 vssd1 vccd1 vccd1 _17209_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5767 _17661_/Q vssd1 vssd1 vccd1 vccd1 hold5767/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5778 _13624_/X vssd1 vssd1 vccd1 vccd1 _17661_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5789 _17214_/Q vssd1 vssd1 vccd1 vccd1 hold5789/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout500 _10538_/S vssd1 vssd1 vccd1 vccd1 _10985_/S sky130_fd_sc_hd__buf_4
XFILLER_0_228_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout511 _10475_/S vssd1 vssd1 vccd1 vccd1 _10571_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09906_ _09912_/A _09906_/B vssd1 vssd1 vccd1 vccd1 _09906_/X sky130_fd_sc_hd__or2_1
Xfanout522 _09340_/X vssd1 vssd1 vccd1 vccd1 _15490_/B1 sky130_fd_sc_hd__buf_8
XFILLER_0_158_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout533 _09124_/Y vssd1 vssd1 vccd1 vccd1 _09177_/A2 sky130_fd_sc_hd__buf_4
Xfanout544 _08448_/Y vssd1 vssd1 vccd1 vccd1 _08486_/B sky130_fd_sc_hd__clkbuf_8
Xfanout555 _08228_/Y vssd1 vssd1 vccd1 vccd1 _08262_/B sky130_fd_sc_hd__buf_6
Xfanout566 _07993_/Y vssd1 vssd1 vccd1 vccd1 _08033_/B sky130_fd_sc_hd__clkbuf_8
X_09837_ _09933_/A _09837_/B vssd1 vssd1 vccd1 vccd1 _09837_/X sky130_fd_sc_hd__or2_1
Xfanout577 _14572_/X vssd1 vssd1 vccd1 vccd1 _14612_/B sky130_fd_sc_hd__buf_6
Xfanout588 _13225_/B vssd1 vssd1 vccd1 vccd1 _13305_/B sky130_fd_sc_hd__buf_4
XFILLER_0_232_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout599 _12985_/S vssd1 vssd1 vccd1 vccd1 _13000_/S sky130_fd_sc_hd__buf_6
XFILLER_0_38_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09768_ _09954_/A _09768_/B vssd1 vssd1 vccd1 vccd1 _09768_/X sky130_fd_sc_hd__or2_1
XFILLER_0_214_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08719_ hold82/X hold634/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold635/A sky130_fd_sc_hd__mux2_1
XFILLER_0_69_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09699_ _09987_/A _09699_/B vssd1 vssd1 vccd1 vccd1 _09699_/X sky130_fd_sc_hd__or2_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11730_ hold4345/X _11637_/A _11729_/X vssd1 vssd1 vccd1 vccd1 _11730_/Y sky130_fd_sc_hd__a21oi_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11661_ _11661_/A _11661_/B vssd1 vssd1 vccd1 vccd1 _11661_/X sky130_fd_sc_hd__or2_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13400_ hold2575/X hold4514/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13401_/B sky130_fd_sc_hd__mux2_1
X_10612_ _11206_/A _10612_/B vssd1 vssd1 vccd1 vccd1 _16694_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_36_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14380_ _14380_/A hold98/X vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__and2_1
X_11592_ _12234_/A _11592_/B vssd1 vssd1 vccd1 vccd1 _11592_/X sky130_fd_sc_hd__or2_1
XFILLER_0_187_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13331_ hold2355/X hold4270/X _13811_/C vssd1 vssd1 vccd1 vccd1 _13332_/B sky130_fd_sc_hd__mux2_1
X_10543_ hold3905/X _10637_/B _10542_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10543_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16050_ _18424_/CLK _16050_/D vssd1 vssd1 vccd1 vccd1 hold556/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13262_ _13262_/A _13294_/B vssd1 vssd1 vccd1 vccd1 _13262_/X sky130_fd_sc_hd__or2_1
XFILLER_0_165_1363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10474_ hold3672/X _10568_/B _10473_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _10474_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15001_ hold1861/X _15004_/B _15000_/Y _15146_/C1 vssd1 vssd1 vccd1 vccd1 _15001_/X
+ sky130_fd_sc_hd__o211a_1
X_12213_ _13797_/A _12213_/B vssd1 vssd1 vccd1 vccd1 _12213_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13193_ _13193_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13193_/X sky130_fd_sc_hd__and2_1
XFILLER_0_20_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12144_ _12240_/A _12144_/B vssd1 vssd1 vccd1 vccd1 _12144_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12075_ _12267_/A _12075_/B vssd1 vssd1 vccd1 vccd1 _12075_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16952_ _17874_/CLK _16952_/D vssd1 vssd1 vccd1 vccd1 _16952_/Q sky130_fd_sc_hd__dfxtp_1
X_15903_ _17321_/CLK _15903_/D vssd1 vssd1 vccd1 vccd1 hold504/A sky130_fd_sc_hd__dfxtp_1
X_11026_ hold5074/X _11225_/B _11025_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _11026_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16883_ _18054_/CLK _16883_/D vssd1 vssd1 vccd1 vccd1 _16883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15834_ _17722_/CLK _15834_/D vssd1 vssd1 vccd1 vccd1 _15834_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12977_ hold3787/X _12976_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12978_/B sky130_fd_sc_hd__mux2_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15765_ _17748_/CLK _15765_/D vssd1 vssd1 vccd1 vccd1 _15765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_242_wb_clk_i clkbuf_6_57_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18236_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _17512_/CLK _17504_/D vssd1 vssd1 vccd1 vccd1 _17504_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14716_ _15163_/A _14720_/B vssd1 vssd1 vccd1 vccd1 _14716_/Y sky130_fd_sc_hd__nand2_1
X_11928_ _12216_/A _11928_/B vssd1 vssd1 vccd1 vccd1 _11928_/X sky130_fd_sc_hd__or2_1
X_15696_ _17264_/CLK _15696_/D vssd1 vssd1 vccd1 vccd1 _15696_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14647_ hold2723/X _14666_/B _14646_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _14647_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17435_ _17435_/CLK _17435_/D vssd1 vssd1 vccd1 vccd1 _17435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11859_ _12255_/A _11859_/B vssd1 vssd1 vccd1 vccd1 _11859_/X sky130_fd_sc_hd__or2_1
XFILLER_0_200_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_18 _13164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_29 _13180_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14578_ hold911/X _14622_/B vssd1 vssd1 vccd1 vccd1 _14578_/X sky130_fd_sc_hd__or2_1
X_17366_ _17514_/CLK _17366_/D vssd1 vssd1 vccd1 vccd1 _17366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16317_ _16319_/CLK _16317_/D vssd1 vssd1 vccd1 vccd1 _16317_/Q sky130_fd_sc_hd__dfxtp_1
X_13529_ hold1198/X hold3646/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13530_/B sky130_fd_sc_hd__mux2_1
X_17297_ _17297_/CLK _17297_/D vssd1 vssd1 vccd1 vccd1 _17297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16248_ _17427_/CLK _16248_/D vssd1 vssd1 vccd1 vccd1 _16248_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5008 _16486_/Q vssd1 vssd1 vccd1 vccd1 hold5008/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5019 _10747_/X vssd1 vssd1 vccd1 vccd1 _16739_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput103 _13129_/A vssd1 vssd1 vccd1 vccd1 hold5868/A sky130_fd_sc_hd__buf_6
XFILLER_0_141_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput114 hold5923/X vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_12
Xhold4307 _12342_/Y vssd1 vssd1 vccd1 vccd1 _12343_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16179_ _17464_/CLK _16179_/D vssd1 vssd1 vccd1 vccd1 _16179_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4318 _16726_/Q vssd1 vssd1 vccd1 vccd1 hold4318/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput125 hold5931/X vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_12
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4329 _11148_/Y vssd1 vssd1 vccd1 vccd1 _11149_/B sky130_fd_sc_hd__dlygate4sd3_1
Xoutput136 hold4199/X vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_12
XFILLER_0_220_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3606 _16382_/Q vssd1 vssd1 vccd1 vccd1 hold3606/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3617 _16413_/Q vssd1 vssd1 vccd1 vccd1 hold3617/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3628 _16479_/Q vssd1 vssd1 vccd1 vccd1 hold3628/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3639 _12527_/X vssd1 vssd1 vccd1 vccd1 _12528_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2905 _15530_/X vssd1 vssd1 vccd1 vccd1 _18443_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2916 _16152_/Q vssd1 vssd1 vccd1 vccd1 hold2916/X sky130_fd_sc_hd__dlygate4sd3_1
X_07952_ _14461_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07952_/X sky130_fd_sc_hd__or2_1
Xhold2927 _09294_/X vssd1 vssd1 vccd1 vccd1 _16257_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2938 _15667_/Q vssd1 vssd1 vccd1 vccd1 hold2938/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2949 _15194_/X vssd1 vssd1 vccd1 vccd1 _18379_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07883_ hold405/X hold337/X hold509/X hold444/X vssd1 vssd1 vccd1 vccd1 _14789_/A
+ sky130_fd_sc_hd__or4bb_4
XFILLER_0_177_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09622_ hold4463/X _10028_/B _09621_/X _15048_/A vssd1 vssd1 vccd1 vccd1 _09622_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09553_ hold3946/X _10049_/B _09552_/X _15146_/C1 vssd1 vssd1 vccd1 vccd1 _09553_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08504_ _08504_/A _14897_/A vssd1 vssd1 vccd1 vccd1 _08517_/B sky130_fd_sc_hd__or2_2
XFILLER_0_37_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09484_ hold5981/X _09484_/B _09484_/C vssd1 vssd1 vccd1 vccd1 _16322_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_77_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08435_ _14543_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08435_/X sky130_fd_sc_hd__or2_1
XFILLER_0_77_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08366_ _09313_/A hold1198/X hold115/X vssd1 vssd1 vccd1 vccd1 _08367_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08297_ _14461_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08297_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_wb_clk_i clkbuf_6_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18041_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5520 _13378_/X vssd1 vssd1 vccd1 vccd1 _17579_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5531 _16980_/Q vssd1 vssd1 vccd1 vccd1 hold5531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5542 _10660_/X vssd1 vssd1 vccd1 vccd1 _16710_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5553 _17734_/Q vssd1 vssd1 vccd1 vccd1 hold5553/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5564 _13477_/X vssd1 vssd1 vccd1 vccd1 _17612_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4830 _09745_/X vssd1 vssd1 vccd1 vccd1 _16405_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5575 _17173_/Q vssd1 vssd1 vccd1 vccd1 hold5575/X sky130_fd_sc_hd__dlygate4sd3_1
X_10190_ hold2739/X _16554_/Q _10985_/S vssd1 vssd1 vccd1 vccd1 _10191_/B sky130_fd_sc_hd__mux2_1
Xhold4841 _17724_/Q vssd1 vssd1 vccd1 vccd1 hold4841/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5586 _11317_/X vssd1 vssd1 vccd1 vccd1 _16929_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5597 _17638_/Q vssd1 vssd1 vccd1 vccd1 hold5597/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4852 _12010_/X vssd1 vssd1 vccd1 vccd1 _17160_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4863 _17174_/Q vssd1 vssd1 vccd1 vccd1 hold4863/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4874 _11908_/X vssd1 vssd1 vccd1 vccd1 _17126_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4885 _17243_/Q vssd1 vssd1 vccd1 vccd1 hold4885/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout330 _10470_/A vssd1 vssd1 vccd1 vccd1 _10530_/A sky130_fd_sc_hd__buf_4
XFILLER_0_22_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4896 _11512_/X vssd1 vssd1 vccd1 vccd1 _16994_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout341 _12405_/S vssd1 vssd1 vccd1 vccd1 _12441_/S sky130_fd_sc_hd__buf_8
Xfanout352 _08779_/S vssd1 vssd1 vccd1 vccd1 _08793_/S sky130_fd_sc_hd__buf_8
XFILLER_0_195_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout363 _15227_/B vssd1 vssd1 vccd1 vccd1 _15233_/B sky130_fd_sc_hd__buf_6
Xfanout374 hold510/X vssd1 vssd1 vccd1 vccd1 _15018_/B sky130_fd_sc_hd__buf_6
XFILLER_0_22_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout385 _14788_/Y vssd1 vssd1 vccd1 vccd1 _14826_/B sky130_fd_sc_hd__buf_6
XFILLER_0_226_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12900_ _12906_/A _12900_/B vssd1 vssd1 vccd1 vccd1 _17476_/D sky130_fd_sc_hd__and2_1
Xfanout396 _14501_/Y vssd1 vssd1 vccd1 vccd1 _14537_/B sky130_fd_sc_hd__buf_8
XFILLER_0_214_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13880_ _17747_/Q _13880_/B _13880_/C vssd1 vssd1 vccd1 vccd1 _13880_/X sky130_fd_sc_hd__and3_1
XFILLER_0_202_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12831_ _12837_/A _12831_/B vssd1 vssd1 vccd1 vccd1 _17453_/D sky130_fd_sc_hd__and2_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_232_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_232_1228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ hold2000/X _15547_/B _15549_/X _12837_/A vssd1 vssd1 vccd1 vccd1 _15550_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12762_ _12810_/A _12762_/B vssd1 vssd1 vccd1 vccd1 _17430_/D sky130_fd_sc_hd__and2_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14501_ _15182_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14501_/Y sky130_fd_sc_hd__nor2_2
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ hold5653/X _11717_/B _11712_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _11713_/X
+ sky130_fd_sc_hd__o211a_1
X_15481_ _15481_/A1 _15474_/X _15480_/X _15481_/B1 hold5959/A vssd1 vssd1 vccd1 vccd1
+ _15481_/X sky130_fd_sc_hd__a32o_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12843_/A _12693_/B vssd1 vssd1 vccd1 vccd1 _17407_/D sky130_fd_sc_hd__and2_1
XFILLER_0_210_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ hold2629/X _14433_/B _14431_/Y _14354_/A vssd1 vssd1 vccd1 vccd1 _14432_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _17908_/CLK _17220_/D vssd1 vssd1 vccd1 vccd1 _17220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11644_ hold5382/X _11744_/B _11643_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _11644_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17151_ _17247_/CLK _17151_/D vssd1 vssd1 vccd1 vccd1 _17151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14363_ _14596_/A hold1777/X _14381_/S vssd1 vssd1 vccd1 vccd1 _14363_/X sky130_fd_sc_hd__mux2_1
Xinput16 input16/A vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_1
X_11575_ hold5189/X _11765_/B _11574_/X _14346_/A vssd1 vssd1 vccd1 vccd1 _11575_/X
+ sky130_fd_sc_hd__o211a_1
Xinput27 input27/A vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_1
X_16102_ _17325_/CLK _16102_/D vssd1 vssd1 vccd1 vccd1 _16102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput38 input38/A vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_1
X_13314_ _13314_/A _13314_/B vssd1 vssd1 vccd1 vccd1 _13314_/X sky130_fd_sc_hd__or2_1
X_10526_ hold2153/X _16666_/Q _10640_/C vssd1 vssd1 vccd1 vccd1 _10527_/B sky130_fd_sc_hd__mux2_1
Xinput49 input49/A vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_6
X_17082_ _17834_/CLK _17082_/D vssd1 vssd1 vccd1 vccd1 _17082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14294_ _14974_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14294_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16033_ _18413_/CLK _16033_/D vssd1 vssd1 vccd1 vccd1 hold292/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13245_ _13244_/X hold3420/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13245_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_165_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10457_ hold1754/X hold3795/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10458_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_110_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13176_ _13169_/X _13175_/X _13296_/B1 vssd1 vssd1 vccd1 vccd1 _17540_/D sky130_fd_sc_hd__o21a_1
X_10388_ hold1033/X _16620_/Q _10625_/C vssd1 vssd1 vccd1 vccd1 _10389_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12127_ hold4968/X _12317_/B _12126_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _12127_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_237_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17984_ _18016_/CLK _17984_/D vssd1 vssd1 vccd1 vccd1 _17984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_236_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12058_ hold4915/X _12374_/B _12057_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _12058_/X
+ sky130_fd_sc_hd__o211a_1
X_16935_ _18429_/CLK _16935_/D vssd1 vssd1 vccd1 vccd1 _16935_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_423_wb_clk_i clkbuf_6_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17229_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_174_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11009_ hold3110/X hold5201/X _11171_/C vssd1 vssd1 vccd1 vccd1 _11010_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_74_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16866_ _18069_/CLK _16866_/D vssd1 vssd1 vccd1 vccd1 _16866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_215_1404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15817_ _17697_/CLK _15817_/D vssd1 vssd1 vccd1 vccd1 _15817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16797_ _18059_/CLK _16797_/D vssd1 vssd1 vccd1 vccd1 _16797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15748_ _17221_/CLK _15748_/D vssd1 vssd1 vccd1 vccd1 _15748_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15679_ _17107_/CLK _15679_/D vssd1 vssd1 vccd1 vccd1 _15679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08220_ hold2671/X _08213_/B _08219_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _08220_/X
+ sky130_fd_sc_hd__o211a_1
X_17418_ _17427_/CLK _17418_/D vssd1 vssd1 vccd1 vccd1 _17418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18398_ _18398_/CLK _18398_/D vssd1 vssd1 vccd1 vccd1 _18398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08151_ _08151_/A _08151_/B vssd1 vssd1 vccd1 vccd1 _15714_/D sky130_fd_sc_hd__and2_1
X_17349_ _17512_/CLK _17349_/D vssd1 vssd1 vccd1 vccd1 _17349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08082_ _15215_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08082_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_28_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4104 _11113_/X vssd1 vssd1 vccd1 vccd1 _16861_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4115 _17027_/Q vssd1 vssd1 vccd1 vccd1 hold4115/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4126 _13495_/X vssd1 vssd1 vccd1 vccd1 _17618_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4137 _17501_/Q vssd1 vssd1 vccd1 vccd1 hold4137/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3403 _09397_/X vssd1 vssd1 vccd1 vccd1 _16285_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4148 _10924_/X vssd1 vssd1 vccd1 vccd1 _16798_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3414 _16333_/Q vssd1 vssd1 vccd1 vccd1 _13134_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4159 _17078_/Q vssd1 vssd1 vccd1 vccd1 _11762_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3425 _16339_/Q vssd1 vssd1 vccd1 vccd1 _13182_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3436 _10581_/Y vssd1 vssd1 vccd1 vccd1 _10582_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08984_ _12438_/A _08984_/B vssd1 vssd1 vccd1 vccd1 _16109_/D sky130_fd_sc_hd__and2_1
XTAP_5609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3447 _16327_/Q vssd1 vssd1 vccd1 vccd1 _13086_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2702 _14313_/X vssd1 vssd1 vccd1 vccd1 _17956_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3458 _10006_/Y vssd1 vssd1 vccd1 vccd1 _16492_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2713 _17993_/Q vssd1 vssd1 vccd1 vccd1 hold2713/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2724 _14647_/X vssd1 vssd1 vccd1 vccd1 _18116_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3469 _10593_/Y vssd1 vssd1 vccd1 vccd1 _10594_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2735 _18220_/Q vssd1 vssd1 vccd1 vccd1 hold2735/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2746 _15534_/X vssd1 vssd1 vccd1 vccd1 _18445_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07935_ hold1831/X _07924_/B _07934_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _07935_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2757 _15554_/X vssd1 vssd1 vccd1 vccd1 _18455_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_164_wb_clk_i clkbuf_6_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18369_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2768 _09308_/X vssd1 vssd1 vccd1 vccd1 _16264_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2779 _17823_/Q vssd1 vssd1 vccd1 vccd1 hold2779/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07866_ hold2318/X _07865_/B _07865_/Y _08143_/A vssd1 vssd1 vccd1 vccd1 _07866_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09605_ hold1609/X hold3648/X _10004_/C vssd1 vssd1 vccd1 vccd1 _09606_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_155_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07797_ hold5978/X _07788_/Y _07809_/B hold3129/X _11158_/A vssd1 vssd1 vccd1 vccd1
+ _07797_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09536_ hold2977/X _13158_/A _10022_/C vssd1 vssd1 vccd1 vccd1 _09537_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09467_ _09472_/C _09465_/A _09466_/Y vssd1 vssd1 vccd1 vccd1 _09467_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_210_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_231_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08418_ hold1045/X _08442_/A2 _08417_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _08418_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09398_ hold337/X hold509/A hold353/A vssd1 vssd1 vccd1 vccd1 _09398_/X sky130_fd_sc_hd__and3_1
XFILLER_0_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08349_ _08385_/A _08349_/B vssd1 vssd1 vccd1 vccd1 _15806_/D sky130_fd_sc_hd__and2_1
XFILLER_0_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11360_ hold1239/X hold4018/X _12317_/C vssd1 vssd1 vccd1 vccd1 _11361_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_6_7_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6040 data_in[19] vssd1 vssd1 vccd1 vccd1 hold212/A sky130_fd_sc_hd__dlygate4sd3_1
X_10311_ _10515_/A _10311_/B vssd1 vssd1 vccd1 vccd1 _10311_/X sky130_fd_sc_hd__or2_1
Xhold6051 _17870_/Q vssd1 vssd1 vccd1 vccd1 hold6051/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6062 _18071_/Q vssd1 vssd1 vccd1 vccd1 hold6062/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6073 _18328_/Q vssd1 vssd1 vccd1 vccd1 hold6073/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11291_ hold2070/X hold4717/X _12242_/S vssd1 vssd1 vccd1 vccd1 _11292_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_225_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6084 _18294_/Q vssd1 vssd1 vccd1 vccd1 hold6084/X sky130_fd_sc_hd__dlygate4sd3_1
X_13030_ _17520_/Q _13034_/D hold904/A vssd1 vssd1 vccd1 vccd1 hold896/A sky130_fd_sc_hd__and3_1
Xhold6095 la_data_in[24] vssd1 vssd1 vccd1 vccd1 hold286/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5350 _11395_/X vssd1 vssd1 vccd1 vccd1 _16955_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10242_ _10470_/A _10242_/B vssd1 vssd1 vccd1 vccd1 _10242_/X sky130_fd_sc_hd__or2_1
Xhold5361 hold6134/X vssd1 vssd1 vccd1 vccd1 _07826_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_104_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5372 _16767_/Q vssd1 vssd1 vccd1 vccd1 hold5372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5383 _11644_/X vssd1 vssd1 vccd1 vccd1 _17038_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5394 _17649_/Q vssd1 vssd1 vccd1 vccd1 hold5394/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4660 _17691_/Q vssd1 vssd1 vccd1 vccd1 hold4660/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10173_ _10563_/A _10173_/B vssd1 vssd1 vccd1 vccd1 _10173_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4671 _11809_/X vssd1 vssd1 vccd1 vccd1 _17093_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4682 _13315_/X vssd1 vssd1 vccd1 vccd1 _17558_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4693 _16426_/Q vssd1 vssd1 vccd1 vccd1 hold4693/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3970 _16653_/Q vssd1 vssd1 vccd1 vccd1 hold3970/X sky130_fd_sc_hd__dlygate4sd3_1
X_14981_ hold2842/X _15004_/B _14980_/X _15473_/A vssd1 vssd1 vccd1 vccd1 _14981_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3981 _10993_/X vssd1 vssd1 vccd1 vccd1 _16821_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout160 _13814_/B vssd1 vssd1 vccd1 vccd1 _13808_/B sky130_fd_sc_hd__clkbuf_8
Xhold3992 _11062_/X vssd1 vssd1 vccd1 vccd1 _16844_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout171 fanout210/X vssd1 vssd1 vccd1 vccd1 _12217_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_233_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16720_ _18051_/CLK _16720_/D vssd1 vssd1 vccd1 vccd1 _16720_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout182 _11071_/A2 vssd1 vssd1 vccd1 vccd1 _11165_/B sky130_fd_sc_hd__clkbuf_8
Xfanout193 _13877_/B vssd1 vssd1 vccd1 vccd1 _13880_/B sky130_fd_sc_hd__clkbuf_8
X_13932_ hold235/X _17774_/Q hold297/X vssd1 vssd1 vccd1 vccd1 hold298/A sky130_fd_sc_hd__mux2_1
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_214_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16651_ _18217_/CLK _16651_/D vssd1 vssd1 vccd1 vccd1 _16651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13863_ hold4293/X _13737_/A _13862_/X vssd1 vssd1 vccd1 vccd1 _13864_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12814_ hold1823/X hold3380/X _12838_/S vssd1 vssd1 vccd1 vccd1 _12814_/X sky130_fd_sc_hd__mux2_1
X_15602_ _17250_/CLK _15602_/D vssd1 vssd1 vccd1 vccd1 _15602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16582_ _18236_/CLK _16582_/D vssd1 vssd1 vccd1 vccd1 _16582_/Q sky130_fd_sc_hd__dfxtp_1
X_13794_ _13794_/A _13794_/B vssd1 vssd1 vccd1 vccd1 _13794_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18321_ _18321_/CLK _18321_/D vssd1 vssd1 vccd1 vccd1 _18321_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _16246_/Q hold3175/X _12811_/S vssd1 vssd1 vccd1 vccd1 _12745_/X sky130_fd_sc_hd__mux2_1
X_15533_ _15533_/A _15549_/B vssd1 vssd1 vccd1 vccd1 _15533_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18252_ _18342_/CLK _18252_/D vssd1 vssd1 vccd1 vccd1 _18252_/Q sky130_fd_sc_hd__dfxtp_1
X_15464_ _15482_/A _15464_/B vssd1 vssd1 vccd1 vccd1 _18422_/D sky130_fd_sc_hd__and2_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12676_ hold2006/X _17403_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12676_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_210_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14415_ _14988_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14415_/X sky130_fd_sc_hd__or2_1
X_17203_ _17897_/CLK _17203_/D vssd1 vssd1 vccd1 vccd1 _17203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11627_ hold2844/X hold5374/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11628_/B sky130_fd_sc_hd__mux2_1
X_18183_ _18197_/CLK _18183_/D vssd1 vssd1 vccd1 vccd1 _18183_/Q sky130_fd_sc_hd__dfxtp_1
X_15395_ hold611/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15395_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17134_ _17262_/CLK _17134_/D vssd1 vssd1 vccd1 vccd1 _17134_/Q sky130_fd_sc_hd__dfxtp_1
X_14346_ _14346_/A _14346_/B vssd1 vssd1 vccd1 vccd1 _17972_/D sky130_fd_sc_hd__and2_1
XFILLER_0_181_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11558_ hold1010/X hold5111/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11559_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_53_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold608 hold608/A vssd1 vssd1 vccd1 vccd1 hold608/X sky130_fd_sc_hd__dlygate4sd3_1
X_10509_ _10551_/A _10509_/B vssd1 vssd1 vccd1 vccd1 _10509_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17065_ _17981_/CLK _17065_/D vssd1 vssd1 vccd1 vccd1 _17065_/Q sky130_fd_sc_hd__dfxtp_1
Xhold619 hold619/A vssd1 vssd1 vccd1 vccd1 hold619/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14277_ hold1402/X _14272_/B _14276_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14277_/X
+ sky130_fd_sc_hd__o211a_1
X_11489_ hold2989/X _16987_/Q _12317_/C vssd1 vssd1 vccd1 vccd1 _11490_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16016_ _18423_/CLK _16016_/D vssd1 vssd1 vccd1 vccd1 _16016_/Q sky130_fd_sc_hd__dfxtp_1
X_13228_ hold3590/X _13227_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13228_/X sky130_fd_sc_hd__mux2_4
XFILLER_0_111_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13159_ _13199_/A1 _13157_/X _13158_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13159_/X
+ sky130_fd_sc_hd__o211a_2
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2009 _18287_/Q vssd1 vssd1 vccd1 vccd1 hold2009/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17967_ _17967_/CLK _17967_/D vssd1 vssd1 vccd1 vccd1 _17967_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1308 _08198_/X vssd1 vssd1 vccd1 vccd1 _15735_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1319 _16201_/Q vssd1 vssd1 vccd1 vccd1 hold1319/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16918_ _17936_/CLK _16918_/D vssd1 vssd1 vccd1 vccd1 _16918_/Q sky130_fd_sc_hd__dfxtp_1
X_17898_ _17898_/CLK _17898_/D vssd1 vssd1 vccd1 vccd1 _17898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16849_ _18052_/CLK _16849_/D vssd1 vssd1 vccd1 vccd1 _16849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09321_ _15543_/A _09323_/B vssd1 vssd1 vccd1 vccd1 _09321_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_165_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _12810_/A hold952/X vssd1 vssd1 vccd1 vccd1 hold953/A sky130_fd_sc_hd__and2_1
XFILLER_0_146_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08203_ _15537_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08203_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09183_ hold6069/X _09218_/B _09182_/X _12777_/A vssd1 vssd1 vccd1 vccd1 _09183_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08134_ _14604_/A _15706_/Q _08152_/S vssd1 vssd1 vccd1 vccd1 _08134_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08065_ hold1293/X _08097_/A2 _08064_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _08065_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_226_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3200 _16537_/Q vssd1 vssd1 vccd1 vccd1 hold3200/X sky130_fd_sc_hd__buf_1
XTAP_6107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_345_wb_clk_i clkbuf_6_42_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17705_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3211 _12806_/X vssd1 vssd1 vccd1 vccd1 _12807_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3222 _17500_/Q vssd1 vssd1 vccd1 vccd1 hold3222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3233 _16497_/Q vssd1 vssd1 vccd1 vccd1 _10019_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3244 _10465_/X vssd1 vssd1 vccd1 vccd1 _16645_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3255 _16702_/Q vssd1 vssd1 vccd1 vccd1 _10634_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2510 _08032_/X vssd1 vssd1 vccd1 vccd1 _15657_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3266 _16481_/Q vssd1 vssd1 vccd1 vccd1 hold3266/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2521 _14093_/X vssd1 vssd1 vccd1 vccd1 _17851_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3277 _09751_/X vssd1 vssd1 vccd1 vccd1 _16407_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08967_ hold185/X hold737/X _08991_/S vssd1 vssd1 vccd1 vccd1 hold738/A sky130_fd_sc_hd__mux2_1
XTAP_5439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2532 _17791_/Q vssd1 vssd1 vccd1 vccd1 hold2532/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2543 _08440_/X vssd1 vssd1 vccd1 vccd1 _15850_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3288 _17465_/Q vssd1 vssd1 vccd1 vccd1 hold3288/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3299 _10423_/X vssd1 vssd1 vccd1 vccd1 _16631_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2554 _14147_/X vssd1 vssd1 vccd1 vccd1 _17877_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1820 _08477_/X vssd1 vssd1 vccd1 vccd1 _15867_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2565 _18450_/Q vssd1 vssd1 vccd1 vccd1 hold2565/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07918_ _15215_/A _07918_/B vssd1 vssd1 vccd1 vccd1 _07918_/Y sky130_fd_sc_hd__nand2_1
Xhold1831 _15611_/Q vssd1 vssd1 vccd1 vccd1 hold1831/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2576 _08495_/X vssd1 vssd1 vccd1 vccd1 _15876_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2587 _18151_/Q vssd1 vssd1 vccd1 vccd1 hold2587/X sky130_fd_sc_hd__dlygate4sd3_1
X_08898_ hold172/X hold802/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08899_/B sky130_fd_sc_hd__mux2_1
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1842 _08312_/X vssd1 vssd1 vccd1 vccd1 _15789_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1853 _18246_/Q vssd1 vssd1 vccd1 vccd1 hold1853/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2598 _14011_/X vssd1 vssd1 vccd1 vccd1 _17811_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1864 _14877_/X vssd1 vssd1 vccd1 vccd1 _18227_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1875 _17958_/Q vssd1 vssd1 vccd1 vccd1 hold1875/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1886 _14532_/X vssd1 vssd1 vccd1 vccd1 _18062_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07849_ _14413_/A _07871_/B vssd1 vssd1 vccd1 vccd1 _07849_/X sky130_fd_sc_hd__or2_1
XFILLER_0_230_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1897 _18007_/Q vssd1 vssd1 vccd1 vccd1 hold1897/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_233_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10860_ _11049_/A _10860_/B vssd1 vssd1 vccd1 vccd1 _10860_/X sky130_fd_sc_hd__or2_1
XFILLER_0_195_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09519_ _09987_/A _09519_/B vssd1 vssd1 vccd1 vccd1 _09519_/X sky130_fd_sc_hd__or2_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _11658_/A _10791_/B vssd1 vssd1 vccd1 vccd1 _10791_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12530_ hold4107/X _12529_/X _12986_/S vssd1 vssd1 vccd1 vccd1 _12530_/X sky130_fd_sc_hd__mux2_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_61_wb_clk_i clkbuf_6_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18014_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12461_ hold679/X _12509_/A2 _12501_/A3 _12460_/X _12410_/A vssd1 vssd1 vccd1 vccd1
+ hold193/A sky130_fd_sc_hd__o311a_1
XFILLER_0_227_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14200_ _15545_/A _14202_/B vssd1 vssd1 vccd1 vccd1 _14200_/Y sky130_fd_sc_hd__nand2_1
X_11412_ _11697_/A _11412_/B vssd1 vssd1 vccd1 vccd1 _11412_/X sky130_fd_sc_hd__or2_1
X_15180_ hold1475/X _15167_/B _15179_/X _15404_/A vssd1 vssd1 vccd1 vccd1 _15180_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12392_ _15374_/A hold395/X vssd1 vssd1 vccd1 vccd1 _17289_/D sky130_fd_sc_hd__and2_1
XFILLER_0_163_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14131_ hold2029/X _14142_/B _14130_/X _14131_/C1 vssd1 vssd1 vccd1 vccd1 _14131_/X
+ sky130_fd_sc_hd__o211a_1
X_11343_ _11631_/A _11343_/B vssd1 vssd1 vccd1 vccd1 _11343_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14062_ _14850_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14062_/X sky130_fd_sc_hd__or2_1
XFILLER_0_240_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11274_ _11658_/A _11274_/B vssd1 vssd1 vccd1 vccd1 _11274_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13013_ hold945/X _13017_/B vssd1 vssd1 vccd1 vccd1 hold946/A sky130_fd_sc_hd__or2_1
Xhold5180 _11962_/X vssd1 vssd1 vccd1 vccd1 _17144_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10225_ hold3997/X _10649_/B _10224_/X _14691_/C1 vssd1 vssd1 vccd1 vccd1 _10225_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5191 _16971_/Q vssd1 vssd1 vccd1 vccd1 hold5191/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4490 _13885_/Y vssd1 vssd1 vccd1 vccd1 _17748_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17821_ _17853_/CLK _17821_/D vssd1 vssd1 vccd1 vccd1 _17821_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10156_ hold4537/X _10628_/B _10155_/X _14697_/C1 vssd1 vssd1 vccd1 vccd1 _10156_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__buf_4
XTAP_5962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17752_ _18462_/CLK _17752_/D vssd1 vssd1 vccd1 vccd1 _17752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10087_ hold3706/X _10568_/B _10086_/X _14769_/C1 vssd1 vssd1 vccd1 vccd1 _10087_/X
+ sky130_fd_sc_hd__o211a_1
X_14964_ _15233_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14964_/X sky130_fd_sc_hd__or2_1
XTAP_5984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16703_ _18229_/CLK _16703_/D vssd1 vssd1 vccd1 vccd1 _16703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13915_ _13935_/A _13915_/B vssd1 vssd1 vccd1 vccd1 _17765_/D sky130_fd_sc_hd__and2_1
XFILLER_0_233_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17683_ _17747_/CLK _17683_/D vssd1 vssd1 vccd1 vccd1 _17683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14895_ hold1283/X hold332/X _14894_/X _14895_/C1 vssd1 vssd1 vccd1 vccd1 _14895_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16634_ _18224_/CLK _16634_/D vssd1 vssd1 vccd1 vccd1 _16634_/Q sky130_fd_sc_hd__dfxtp_1
X_13846_ _13888_/A _13846_/B vssd1 vssd1 vccd1 vccd1 _13846_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16565_ _18181_/CLK _16565_/D vssd1 vssd1 vccd1 vccd1 _16565_/Q sky130_fd_sc_hd__dfxtp_1
X_13777_ hold5193/X _13856_/B _13776_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _13777_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10989_ _11091_/A _10989_/B vssd1 vssd1 vccd1 vccd1 _10989_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18304_ _18421_/CLK _18304_/D vssd1 vssd1 vccd1 vccd1 _18304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15516_ hold2881/X _15560_/A2 _15515_/X _12864_/A vssd1 vssd1 vccd1 vccd1 _15516_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12728_ hold4058/X _12727_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12729_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16496_ _18377_/CLK _16496_/D vssd1 vssd1 vccd1 vccd1 _16496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18235_ _18235_/CLK _18235_/D vssd1 vssd1 vccd1 vccd1 _18235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15447_ _16097_/Q _15487_/B1 _15488_/A2 _16049_/Q vssd1 vssd1 vccd1 vccd1 _15447_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12659_ hold3158/X _12658_/X _12851_/S vssd1 vssd1 vccd1 vccd1 _12660_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_155_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18166_ _18166_/CLK _18166_/D vssd1 vssd1 vccd1 vccd1 _18166_/Q sky130_fd_sc_hd__dfxtp_1
X_15378_ hold668/X _15484_/A2 _15441_/A2 hold781/X vssd1 vssd1 vccd1 vccd1 _15378_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17117_ _17277_/CLK _17117_/D vssd1 vssd1 vccd1 vccd1 _17117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14329_ hold1662/X _14326_/B _14328_/X _14462_/C1 vssd1 vssd1 vccd1 vccd1 _14329_/X
+ sky130_fd_sc_hd__o211a_1
Xhold405 hold405/A vssd1 vssd1 vccd1 vccd1 hold405/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18097_ _18115_/CLK _18097_/D vssd1 vssd1 vccd1 vccd1 _18097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold416 hold420/X vssd1 vssd1 vccd1 vccd1 hold421/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold427 hold427/A vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold438 hold41/X vssd1 vssd1 vccd1 vccd1 hold438/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold449 hold449/A vssd1 vssd1 vccd1 vccd1 hold449/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_6_38_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_38_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_17048_ _17936_/CLK _17048_/D vssd1 vssd1 vccd1 vccd1 _17048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09870_ _09954_/A _09870_/B vssd1 vssd1 vccd1 vccd1 _09870_/X sky130_fd_sc_hd__or2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout907 hold289/X vssd1 vssd1 vccd1 vccd1 _15557_/A sky130_fd_sc_hd__buf_12
XFILLER_0_81_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout918 hold991/X vssd1 vssd1 vccd1 vccd1 _14330_/A sky130_fd_sc_hd__buf_12
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout929 hold1253/X vssd1 vssd1 vccd1 vccd1 _15213_/A sky130_fd_sc_hd__buf_4
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _15254_/A _08821_/B vssd1 vssd1 vccd1 vccd1 _16029_/D sky130_fd_sc_hd__and2_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1105 hold1151/X vssd1 vssd1 vccd1 vccd1 hold1152/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 _08245_/X vssd1 vssd1 vccd1 vccd1 _15757_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08752_ _15344_/A _08752_/B vssd1 vssd1 vccd1 vccd1 _15996_/D sky130_fd_sc_hd__and2_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1127 _18068_/Q vssd1 vssd1 vccd1 vccd1 hold1127/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1138 hold1138/A vssd1 vssd1 vccd1 vccd1 _15173_/A sky130_fd_sc_hd__buf_12
XFILLER_0_174_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1149 _16261_/Q vssd1 vssd1 vccd1 vccd1 hold1149/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08683_ hold673/X hold856/X _08721_/S vssd1 vssd1 vccd1 vccd1 hold857/A sky130_fd_sc_hd__mux2_1
XFILLER_0_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09304_ hold3055/X _09323_/B _09303_/X _12906_/A vssd1 vssd1 vccd1 vccd1 _09304_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09235_ _14166_/A hold1269/X hold271/X vssd1 vssd1 vccd1 vccd1 _09235_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09166_ _15549_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09166_/X sky130_fd_sc_hd__or2_1
XFILLER_0_17_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08117_ _13933_/A _08117_/B vssd1 vssd1 vccd1 vccd1 _15697_/D sky130_fd_sc_hd__and2_1
X_09097_ hold1702/X _09102_/B _09096_/X _12978_/A vssd1 vssd1 vccd1 vccd1 _09097_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08048_ hold355/X _14627_/A vssd1 vssd1 vccd1 vccd1 _08048_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_222_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold950 hold967/X vssd1 vssd1 vccd1 vccd1 hold950/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold961 hold961/A vssd1 vssd1 vccd1 vccd1 hold961/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 hold972/A vssd1 vssd1 vccd1 vccd1 hold972/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 hold983/A vssd1 vssd1 vccd1 vccd1 hold983/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold994 hold994/A vssd1 vssd1 vccd1 vccd1 hold994/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3030 _09320_/X vssd1 vssd1 vccd1 vccd1 _16270_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10010_ _16494_/Q _10022_/B _10022_/C vssd1 vssd1 vccd1 vccd1 _10010_/X sky130_fd_sc_hd__and3_1
Xhold3041 _15615_/Q vssd1 vssd1 vccd1 vccd1 hold3041/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3052 _15015_/X vssd1 vssd1 vccd1 vccd1 _18293_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3063 _17783_/Q vssd1 vssd1 vccd1 vccd1 hold3063/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09999_ _13110_/A _11067_/A _09998_/X vssd1 vssd1 vccd1 vccd1 _09999_/Y sky130_fd_sc_hd__a21oi_1
Xhold3074 _15595_/Q vssd1 vssd1 vccd1 vccd1 hold3074/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2340 _15806_/Q vssd1 vssd1 vccd1 vccd1 hold2340/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3085 _13047_/X vssd1 vssd1 vccd1 vccd1 _13048_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2351 _18126_/Q vssd1 vssd1 vccd1 vccd1 hold2351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3096 _07957_/X vssd1 vssd1 vccd1 vccd1 _15621_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2362 _09296_/X vssd1 vssd1 vccd1 vccd1 _16258_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2373 _15649_/Q vssd1 vssd1 vccd1 vccd1 hold2373/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2384 _17863_/Q vssd1 vssd1 vccd1 vccd1 hold2384/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1650 _15627_/Q vssd1 vssd1 vccd1 vccd1 hold1650/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2395 _08489_/X vssd1 vssd1 vccd1 vccd1 _15873_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_230_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ _13749_/A _11961_/B vssd1 vssd1 vccd1 vccd1 _11961_/X sky130_fd_sc_hd__or2_1
XFILLER_0_58_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1661 _14045_/X vssd1 vssd1 vccd1 vccd1 _17828_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1672 _15748_/Q vssd1 vssd1 vccd1 vccd1 hold1672/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1683 _14293_/X vssd1 vssd1 vccd1 vccd1 _17946_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1694 _15750_/Q vssd1 vssd1 vccd1 vccd1 hold1694/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10912_ hold5618/X _11213_/B _10911_/X _14342_/A vssd1 vssd1 vccd1 vccd1 _10912_/X
+ sky130_fd_sc_hd__o211a_1
X_13700_ hold2406/X hold4943/X _13817_/C vssd1 vssd1 vccd1 vccd1 _13701_/B sky130_fd_sc_hd__mux2_1
X_14680_ _14681_/A _14843_/B vssd1 vssd1 vccd1 vccd1 _14680_/Y sky130_fd_sc_hd__nor2_2
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11892_ _12273_/A _11892_/B vssd1 vssd1 vccd1 vccd1 _11892_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13631_ hold1332/X hold4683/X _13862_/C vssd1 vssd1 vccd1 vccd1 _13632_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_184_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10843_ hold3824/X _11222_/B _10842_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _10843_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16350_ _18393_/CLK _16350_/D vssd1 vssd1 vccd1 vccd1 _16350_/Q sky130_fd_sc_hd__dfxtp_1
X_13562_ hold1084/X hold5533/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13563_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10774_ hold3324/X _10013_/B _10773_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _10774_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15301_ _16294_/Q _15477_/A2 _15487_/B1 hold567/X _15300_/X vssd1 vssd1 vccd1 vccd1
+ _15302_/D sky130_fd_sc_hd__a221o_1
X_12513_ _13048_/A hold2264/X _07809_/X _07789_/A vssd1 vssd1 vccd1 vccd1 _12513_/X
+ sky130_fd_sc_hd__a211o_1
X_16281_ _17750_/CLK _16281_/D vssd1 vssd1 vccd1 vccd1 _16281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13493_ hold1669/X hold4123/X _13877_/C vssd1 vssd1 vccd1 vccd1 _13494_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18020_ _18020_/CLK _18020_/D vssd1 vssd1 vccd1 vccd1 _18020_/Q sky130_fd_sc_hd__dfxtp_1
X_12444_ _15374_/A hold279/X vssd1 vssd1 vccd1 vccd1 _17315_/D sky130_fd_sc_hd__and2_1
X_15232_ hold1722/X _15219_/B _15231_/X _08954_/A vssd1 vssd1 vccd1 vccd1 _15232_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_267_wb_clk_i clkbuf_6_56_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18170_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15163_ _15163_/A _15167_/B vssd1 vssd1 vccd1 vccd1 _15163_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12375_ hold4387/X _13749_/A _12374_/X vssd1 vssd1 vccd1 vccd1 _12375_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14114_ hold911/X _14160_/B vssd1 vssd1 vccd1 vccd1 _14114_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11326_ hold5635/X _12305_/B _11325_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11326_/X
+ sky130_fd_sc_hd__o211a_1
X_15094_ hold3008/X hold340/X _15093_/X _15160_/C1 vssd1 vssd1 vccd1 vccd1 _15094_/X
+ sky130_fd_sc_hd__o211a_1
X_14045_ hold1660/X _14040_/B _14044_/X _14462_/C1 vssd1 vssd1 vccd1 vccd1 _14045_/X
+ sky130_fd_sc_hd__o211a_1
X_11257_ hold5639/X _11744_/B _11256_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _11257_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10208_ hold1455/X hold3684/X _10634_/C vssd1 vssd1 vccd1 vccd1 _10209_/B sky130_fd_sc_hd__mux2_1
XTAP_6460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11188_ _11206_/A _11188_/B vssd1 vssd1 vccd1 vccd1 _16886_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_235_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_234_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17804_ _17838_/CLK _17804_/D vssd1 vssd1 vccd1 vccd1 _17804_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10139_ hold1976/X hold3200/X _10595_/C vssd1 vssd1 vccd1 vccd1 _10140_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_175_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15996_ _18406_/CLK _15996_/D vssd1 vssd1 vccd1 vccd1 hold325/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17735_ _17735_/CLK _17735_/D vssd1 vssd1 vccd1 vccd1 _17735_/Q sky130_fd_sc_hd__dfxtp_1
X_14947_ hold2875/X _14946_/B _14946_/Y _15228_/C1 vssd1 vssd1 vccd1 vccd1 _14947_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17666_ _17730_/CLK _17666_/D vssd1 vssd1 vccd1 vccd1 _17666_/Q sky130_fd_sc_hd__dfxtp_1
X_14878_ _15217_/A hold332/X vssd1 vssd1 vccd1 vccd1 _14878_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_159_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_216_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16617_ _18205_/CLK _16617_/D vssd1 vssd1 vccd1 vccd1 _16617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13829_ _17730_/Q _13829_/B _13829_/C vssd1 vssd1 vccd1 vccd1 _13829_/X sky130_fd_sc_hd__and3_1
XFILLER_0_147_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17597_ _17626_/CLK _17597_/D vssd1 vssd1 vccd1 vccd1 _17597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16548_ _18106_/CLK _16548_/D vssd1 vssd1 vccd1 vccd1 _16548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16479_ _18296_/CLK _16479_/D vssd1 vssd1 vccd1 vccd1 _16479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09020_ hold23/X hold326/X _09060_/S vssd1 vssd1 vccd1 vccd1 _09021_/B sky130_fd_sc_hd__mux2_1
X_18218_ _18218_/CLK _18218_/D vssd1 vssd1 vccd1 vccd1 _18218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5905 hold6034/X vssd1 vssd1 vccd1 vccd1 _13081_/A sky130_fd_sc_hd__buf_1
XFILLER_0_170_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18149_ _18149_/CLK _18149_/D vssd1 vssd1 vccd1 vccd1 _18149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold202 hold449/X vssd1 vssd1 vccd1 vccd1 hold450/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5916 hold5916/A vssd1 vssd1 vccd1 vccd1 hold5916/X sky130_fd_sc_hd__buf_2
XFILLER_0_124_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5927 hold5927/A vssd1 vssd1 vccd1 vccd1 hold5927/X sky130_fd_sc_hd__buf_2
Xhold213 hold31/X vssd1 vssd1 vccd1 vccd1 input15/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5938 hold6103/X vssd1 vssd1 vccd1 vccd1 hold5938/X sky130_fd_sc_hd__clkbuf_4
Xhold224 hold25/X vssd1 vssd1 vccd1 vccd1 input5/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5949 _16285_/Q vssd1 vssd1 vccd1 vccd1 hold5949/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 hold97/X vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__clkbuf_8
Xhold246 hold246/A vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold257 hold257/A vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 hold268/A vssd1 vssd1 vccd1 vccd1 hold268/X sky130_fd_sc_hd__buf_1
XFILLER_0_106_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold279 hold279/A vssd1 vssd1 vccd1 vccd1 hold279/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09922_ hold5817/X _10022_/B _09921_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _09922_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout704 _09047_/A vssd1 vssd1 vccd1 vccd1 _15414_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout715 _14368_/A vssd1 vssd1 vccd1 vccd1 _14354_/A sky130_fd_sc_hd__buf_4
XFILLER_0_141_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout726 _12418_/A vssd1 vssd1 vccd1 vccd1 _12410_/A sky130_fd_sc_hd__buf_4
Xfanout737 _09907_/C1 vssd1 vssd1 vccd1 vccd1 _15473_/A sky130_fd_sc_hd__buf_4
X_09853_ hold4638/X _10031_/B _09852_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09853_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 _13777_/C1 vssd1 vssd1 vccd1 vccd1 _08387_/A sky130_fd_sc_hd__buf_4
XFILLER_0_237_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout759 _14131_/C1 vssd1 vssd1 vccd1 vccd1 _13931_/A sky130_fd_sc_hd__buf_4
XFILLER_0_225_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ hold226/X hold310/X _08860_/S vssd1 vssd1 vccd1 vccd1 hold311/A sky130_fd_sc_hd__mux2_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ hold5014/X _11204_/B _09783_/X _15160_/C1 vssd1 vssd1 vccd1 vccd1 _09784_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ hold131/X _15988_/Q _08735_/S vssd1 vssd1 vccd1 vccd1 hold132/A sky130_fd_sc_hd__mux2_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 _11203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_119 hold915/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _12416_/A hold744/X vssd1 vssd1 vccd1 vccd1 _15954_/D sky130_fd_sc_hd__and2_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08597_ _17519_/Q hold948/A vssd1 vssd1 vccd1 vccd1 _08597_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_221_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09218_ _15547_/A _09218_/B vssd1 vssd1 vccd1 vccd1 _09218_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10490_ hold2025/X _16654_/Q _10640_/C vssd1 vssd1 vccd1 vccd1 _10491_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_106_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_360_wb_clk_i clkbuf_6_35_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17270_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_162_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09149_ hold1909/X _09164_/B _09148_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _09149_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12160_ hold4739/X _12350_/B _12159_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _12160_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11111_ hold3017/X _16861_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _11112_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_31_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12091_ hold5156/X _13886_/B _12090_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _17187_/D
+ sky130_fd_sc_hd__o211a_1
Xhold780 hold780/A vssd1 vssd1 vccd1 vccd1 hold780/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 hold791/A vssd1 vssd1 vccd1 vccd1 hold791/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ hold2573/X hold5241/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11043_/B sky130_fd_sc_hd__mux2_1
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15850_ _17678_/CLK _15850_/D vssd1 vssd1 vccd1 vccd1 _15850_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2170 _14845_/X vssd1 vssd1 vccd1 vccd1 _18211_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ hold2664/X _14828_/B _14800_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14801_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2181 _16191_/Q vssd1 vssd1 vccd1 vccd1 hold2181/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2192 _15098_/X vssd1 vssd1 vccd1 vccd1 _18333_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _17648_/CLK _15781_/D vssd1 vssd1 vccd1 vccd1 _15781_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _15244_/A _12993_/B vssd1 vssd1 vccd1 vccd1 _17507_/D sky130_fd_sc_hd__and2_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17520_ _17520_/CLK _17520_/D vssd1 vssd1 vccd1 vccd1 _17520_/Q sky130_fd_sc_hd__dfxtp_2
Xhold1480 _15132_/X vssd1 vssd1 vccd1 vccd1 _18349_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1491 _18372_/Q vssd1 vssd1 vccd1 vccd1 hold1491/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ _14732_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14732_/X sky130_fd_sc_hd__or2_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ hold5731/X _12362_/B _11943_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _11944_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _17452_/CLK _17451_/D vssd1 vssd1 vccd1 vccd1 _17451_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14663_ hold2295/X _14666_/B _14662_/Y _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14663_/X
+ sky130_fd_sc_hd__o211a_1
X_11875_ hold4976/X _12356_/B _11874_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _11875_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_197_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _18315_/CLK _16402_/D vssd1 vssd1 vccd1 vccd1 _16402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10826_ hold1159/X hold4070/X _11210_/C vssd1 vssd1 vccd1 vccd1 _10827_/B sky130_fd_sc_hd__mux2_1
X_13614_ _13719_/A _13614_/B vssd1 vssd1 vccd1 vccd1 _13614_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17382_ _18437_/CLK _17382_/D vssd1 vssd1 vccd1 vccd1 _17382_/Q sky130_fd_sc_hd__dfxtp_1
X_14594_ _14988_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14594_/X sky130_fd_sc_hd__or2_1
XFILLER_0_172_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_448_wb_clk_i clkbuf_6_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17724_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16333_ _18382_/CLK _16333_/D vssd1 vssd1 vccd1 vccd1 _16333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10757_ hold1682/X _16743_/Q _11144_/C vssd1 vssd1 vccd1 vccd1 _10758_/B sky130_fd_sc_hd__mux2_1
X_13545_ _13737_/A _13545_/B vssd1 vssd1 vccd1 vccd1 _13545_/X sky130_fd_sc_hd__or2_1
XFILLER_0_165_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16264_ _17514_/CLK _16264_/D vssd1 vssd1 vccd1 vccd1 _16264_/Q sky130_fd_sc_hd__dfxtp_1
X_13476_ _13752_/A _13476_/B vssd1 vssd1 vccd1 vccd1 _13476_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10688_ hold651/X hold3523/X _11738_/C vssd1 vssd1 vccd1 vccd1 _10689_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18003_ _18066_/CLK hold995/X vssd1 vssd1 vccd1 vccd1 hold994/A sky130_fd_sc_hd__dfxtp_1
X_15215_ _15215_/A _15219_/B vssd1 vssd1 vccd1 vccd1 _15215_/Y sky130_fd_sc_hd__nand2_1
X_12427_ hold92/X hold126/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold127/A sky130_fd_sc_hd__mux2_1
XFILLER_0_2_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16195_ _17476_/CLK _16195_/D vssd1 vssd1 vccd1 vccd1 _16195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15146_ hold2259/X _15167_/B _15145_/X _15146_/C1 vssd1 vssd1 vccd1 vccd1 _15146_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12358_ _13819_/A _12358_/B vssd1 vssd1 vccd1 vccd1 _12358_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_168_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11309_ hold1097/X hold4390/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11310_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15077_ _15185_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15077_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12289_ hold4923/X _12353_/B _12288_/X _12289_/C1 vssd1 vssd1 vccd1 vccd1 _12289_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14028_ _15535_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14028_/X sky130_fd_sc_hd__or2_1
XFILLER_0_177_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15979_ _16098_/CLK _15979_/D vssd1 vssd1 vccd1 vccd1 hold812/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08520_ _18460_/Q _13057_/B vssd1 vssd1 vccd1 vccd1 _08868_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_222_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17718_ _17718_/CLK _17718_/D vssd1 vssd1 vccd1 vccd1 _17718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08451_ hold1647/X _08488_/B _08450_/X _13795_/C1 vssd1 vssd1 vccd1 vccd1 _15854_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17649_ _17745_/CLK _17649_/D vssd1 vssd1 vccd1 vccd1 _17649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08382_ _14330_/A hold1226/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08383_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_189_wb_clk_i clkbuf_6_52_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18387_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_118_wb_clk_i clkbuf_6_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17339_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_143_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09003_ _09003_/A hold619/X vssd1 vssd1 vccd1 vccd1 _16118_/D sky130_fd_sc_hd__and2_1
XFILLER_0_14_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5702 _11677_/X vssd1 vssd1 vccd1 vccd1 _17049_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5713 _12340_/Y vssd1 vssd1 vccd1 vccd1 _17270_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5724 _13809_/Y vssd1 vssd1 vccd1 vccd1 _13810_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5735 _17149_/Q vssd1 vssd1 vccd1 vccd1 hold5735/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5746 _12061_/X vssd1 vssd1 vccd1 vccd1 _17177_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5757 _17140_/Q vssd1 vssd1 vccd1 vccd1 hold5757/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5768 _13528_/X vssd1 vssd1 vccd1 vccd1 _17629_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5779 _17723_/Q vssd1 vssd1 vccd1 vccd1 hold5779/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout501 _10538_/S vssd1 vssd1 vccd1 vccd1 _10040_/C sky130_fd_sc_hd__clkbuf_8
X_09905_ hold1491/X _16459_/Q _10025_/C vssd1 vssd1 vccd1 vccd1 _09906_/B sky130_fd_sc_hd__mux2_1
Xfanout512 _09499_/Y vssd1 vssd1 vccd1 vccd1 _10475_/S sky130_fd_sc_hd__clkbuf_8
Xfanout523 _09340_/X vssd1 vssd1 vccd1 vccd1 _15481_/B1 sky130_fd_sc_hd__buf_4
XFILLER_0_10_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout534 _09124_/Y vssd1 vssd1 vccd1 vccd1 _09164_/B sky130_fd_sc_hd__buf_4
Xfanout545 _08445_/B vssd1 vssd1 vccd1 vccd1 _08439_/B sky130_fd_sc_hd__clkbuf_8
Xfanout556 _08215_/B vssd1 vssd1 vccd1 vccd1 _08225_/B sky130_fd_sc_hd__buf_8
XFILLER_0_77_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09836_ hold1479/X _16436_/Q _10028_/C vssd1 vssd1 vccd1 vccd1 _09837_/B sky130_fd_sc_hd__mux2_1
Xfanout567 _07990_/B vssd1 vssd1 vccd1 vccd1 _07986_/B sky130_fd_sc_hd__buf_6
XFILLER_0_226_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout578 _14572_/X vssd1 vssd1 vccd1 vccd1 _14610_/B sky130_fd_sc_hd__buf_6
Xfanout589 _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13199_/C1 sky130_fd_sc_hd__buf_8
XFILLER_0_226_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_214_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09767_ hold2345/X _16413_/Q _10049_/C vssd1 vssd1 vccd1 vccd1 _09768_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_241_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _12412_/A _08718_/B vssd1 vssd1 vccd1 vccd1 _15980_/D sky130_fd_sc_hd__and2_1
XFILLER_0_154_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _18303_/Q _16390_/Q _09992_/C vssd1 vssd1 vccd1 vccd1 _09699_/B sky130_fd_sc_hd__mux2_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ hold438/X hold528/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08650_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_166_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11660_ hold1321/X hold5321/X _11660_/S vssd1 vssd1 vccd1 vccd1 _11661_/B sky130_fd_sc_hd__mux2_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ hold4238/X _10515_/A _10610_/X vssd1 vssd1 vccd1 vccd1 _10612_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_166_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11591_ hold2029/X hold5655/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11592_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_135_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13330_ hold5801/X _13808_/B _13329_/X _12738_/A vssd1 vssd1 vccd1 vccd1 _13330_/X
+ sky130_fd_sc_hd__o211a_1
X_10542_ _10542_/A _10542_/B vssd1 vssd1 vccd1 vccd1 _10542_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13261_ _13260_/X hold3463/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13261_/X sky130_fd_sc_hd__mux2_1
X_10473_ _10476_/A _10473_/B vssd1 vssd1 vccd1 vccd1 _10473_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15000_ _15161_/A _15004_/B vssd1 vssd1 vccd1 vccd1 _15000_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12212_ hold1459/X hold3870/X _13796_/S vssd1 vssd1 vccd1 vccd1 _12213_/B sky130_fd_sc_hd__mux2_1
X_13192_ _13185_/X _13191_/X _13296_/B1 vssd1 vssd1 vccd1 vccd1 _17542_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_103_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12143_ hold2203/X _17205_/Q _12335_/C vssd1 vssd1 vccd1 vccd1 _12144_/B sky130_fd_sc_hd__mux2_1
X_12074_ hold1091/X hold5785/X _12362_/C vssd1 vssd1 vccd1 vccd1 _12075_/B sky130_fd_sc_hd__mux2_1
X_16951_ _17799_/CLK _16951_/D vssd1 vssd1 vccd1 vccd1 _16951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15902_ _17320_/CLK _15902_/D vssd1 vssd1 vccd1 vccd1 hold587/A sky130_fd_sc_hd__dfxtp_1
X_11025_ _11121_/A _11025_/B vssd1 vssd1 vccd1 vccd1 _11025_/X sky130_fd_sc_hd__or2_1
XFILLER_0_194_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16882_ _18020_/CLK _16882_/D vssd1 vssd1 vccd1 vccd1 _16882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15833_ _17628_/CLK _15833_/D vssd1 vssd1 vccd1 vccd1 _15833_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _17747_/CLK _15764_/D vssd1 vssd1 vccd1 vccd1 _15764_/Q sky130_fd_sc_hd__dfxtp_1
X_12976_ hold2611/X hold3624/X _12985_/S vssd1 vssd1 vccd1 vccd1 _12976_/X sky130_fd_sc_hd__mux2_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17503_ _17512_/CLK _17503_/D vssd1 vssd1 vccd1 vccd1 _17503_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ hold1871/X _14718_/B _14714_/Y _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14715_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11927_ hold2832/X _17133_/Q _12227_/S vssd1 vssd1 vccd1 vccd1 _11928_/B sky130_fd_sc_hd__mux2_1
X_15695_ _17868_/CLK _15695_/D vssd1 vssd1 vccd1 vccd1 _15695_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ _17434_/CLK _17434_/D vssd1 vssd1 vccd1 vccd1 _17434_/Q sky130_fd_sc_hd__dfxtp_1
X_14646_ _15201_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14646_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ _15702_/Q hold5711/X _13463_/S vssd1 vssd1 vccd1 vccd1 _11859_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_282_wb_clk_i clkbuf_6_50_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18063_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_117_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10809_ _11103_/A _10809_/B vssd1 vssd1 vccd1 vccd1 _10809_/X sky130_fd_sc_hd__or2_1
XANTENNA_19 _13164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17365_ _17516_/CLK _17365_/D vssd1 vssd1 vccd1 vccd1 _17365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14577_ hold1730/X _14612_/B _14576_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _14577_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11789_ _17087_/Q _11789_/B _11789_/C vssd1 vssd1 vccd1 vccd1 _11789_/X sky130_fd_sc_hd__and3_1
XFILLER_0_166_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_211_wb_clk_i clkbuf_6_54_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18235_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16316_ _16319_/CLK _16316_/D vssd1 vssd1 vccd1 vccd1 _16316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13528_ hold5767/X _13808_/B _13527_/X _12738_/A vssd1 vssd1 vccd1 vccd1 _13528_/X
+ sky130_fd_sc_hd__o211a_1
X_17296_ _18425_/CLK _17296_/D vssd1 vssd1 vccd1 vccd1 hold701/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16247_ _17425_/CLK hold273/X vssd1 vssd1 vccd1 vccd1 _16247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13459_ hold5597/X _13847_/B _13458_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13459_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5009 _09892_/X vssd1 vssd1 vccd1 vccd1 _16454_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput104 _10651_/A vssd1 vssd1 vccd1 vccd1 io_oeb sky130_fd_sc_hd__buf_12
XFILLER_0_140_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput115 hold5967/X vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_12
Xhold4308 _12343_/Y vssd1 vssd1 vccd1 vccd1 _17271_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16178_ _17462_/CLK _16178_/D vssd1 vssd1 vccd1 vccd1 _16178_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4319 _11187_/Y vssd1 vssd1 vccd1 vccd1 _11188_/B sky130_fd_sc_hd__dlygate4sd3_1
Xoutput126 hold5941/X vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_12
Xoutput137 hold5918/X vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_12
X_15129_ _15183_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15129_/X sky130_fd_sc_hd__or2_1
Xhold3607 _09580_/X vssd1 vssd1 vccd1 vccd1 _16350_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3618 _09673_/X vssd1 vssd1 vccd1 vccd1 _16381_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3629 _09871_/X vssd1 vssd1 vccd1 vccd1 _16447_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07951_ hold1091/X _07991_/A2 _07950_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _07951_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2906 _18181_/Q vssd1 vssd1 vccd1 vccd1 hold2906/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2917 _09075_/X vssd1 vssd1 vccd1 vccd1 _16152_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2928 _18194_/Q vssd1 vssd1 vccd1 vccd1 hold2928/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2939 _08055_/X vssd1 vssd1 vccd1 vccd1 _15667_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07882_ hold1429/X _07865_/B _07881_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _15586_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09621_ _09933_/A _09621_/B vssd1 vssd1 vccd1 vccd1 _09621_/X sky130_fd_sc_hd__or2_1
XFILLER_0_177_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09552_ _09954_/A _09552_/B vssd1 vssd1 vccd1 vccd1 _09552_/X sky130_fd_sc_hd__or2_1
XFILLER_0_214_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08503_ _08504_/A _14897_/A vssd1 vssd1 vccd1 vccd1 _08503_/Y sky130_fd_sc_hd__nor2_2
X_09483_ _09483_/A _09483_/B _09483_/C vssd1 vssd1 vccd1 vccd1 _09483_/X sky130_fd_sc_hd__and3_1
XFILLER_0_194_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08434_ hold2451/X _08433_/B _08433_/Y _13684_/C1 vssd1 vssd1 vccd1 vccd1 _08434_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08365_ _12738_/A _08365_/B vssd1 vssd1 vccd1 vccd1 _15814_/D sky130_fd_sc_hd__and2_1
XFILLER_0_129_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ hold1049/X _08336_/A2 _08295_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _08296_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_229_1383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5510 _11845_/X vssd1 vssd1 vccd1 vccd1 _17105_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5521 _17676_/Q vssd1 vssd1 vccd1 vccd1 hold5521/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5532 _11374_/X vssd1 vssd1 vccd1 vccd1 _16948_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5543 _17195_/Q vssd1 vssd1 vccd1 vccd1 hold5543/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5554 _13747_/X vssd1 vssd1 vccd1 vccd1 _17702_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4820 _10822_/X vssd1 vssd1 vccd1 vccd1 _16764_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5565 _16975_/Q vssd1 vssd1 vccd1 vccd1 hold5565/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4831 _17625_/Q vssd1 vssd1 vccd1 vccd1 hold4831/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5576 _11953_/X vssd1 vssd1 vccd1 vccd1 _17141_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5587 _17652_/Q vssd1 vssd1 vccd1 vccd1 hold5587/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4842 _13717_/X vssd1 vssd1 vccd1 vccd1 _17692_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_86_wb_clk_i clkbuf_6_17_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18400_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4853 _16755_/Q vssd1 vssd1 vccd1 vccd1 hold4853/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5598 _13459_/X vssd1 vssd1 vccd1 vccd1 _17606_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4864 _11956_/X vssd1 vssd1 vccd1 vccd1 _17142_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4875 _17016_/Q vssd1 vssd1 vccd1 vccd1 hold4875/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout320 _10413_/A vssd1 vssd1 vccd1 vccd1 _10515_/A sky130_fd_sc_hd__buf_4
Xhold4886 _12163_/X vssd1 vssd1 vccd1 vccd1 _17211_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4897 _16886_/Q vssd1 vssd1 vccd1 vccd1 hold4897/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_15_wb_clk_i clkbuf_6_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18452_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout331 _10470_/A vssd1 vssd1 vccd1 vccd1 _10554_/A sky130_fd_sc_hd__buf_4
XFILLER_0_121_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout342 _09369_/X vssd1 vssd1 vccd1 vccd1 _15483_/B sky130_fd_sc_hd__clkbuf_8
Xfanout353 _08735_/S vssd1 vssd1 vccd1 vccd1 _08779_/S sky130_fd_sc_hd__buf_8
XFILLER_0_121_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout364 _15181_/Y vssd1 vssd1 vccd1 vccd1 _15221_/B sky130_fd_sc_hd__buf_6
XFILLER_0_195_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout375 hold446/X vssd1 vssd1 vccd1 vccd1 hold447/A sky130_fd_sc_hd__clkbuf_2
Xfanout386 _14780_/B vssd1 vssd1 vccd1 vccd1 _14786_/B sky130_fd_sc_hd__buf_6
XFILLER_0_22_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09819_ _09981_/A _09819_/B vssd1 vssd1 vccd1 vccd1 _09819_/X sky130_fd_sc_hd__or2_1
Xfanout397 _14501_/Y vssd1 vssd1 vccd1 vccd1 _14541_/B sky130_fd_sc_hd__buf_6
XFILLER_0_199_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12830_ hold3390/X _12829_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12830_/X sky130_fd_sc_hd__mux2_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12761_ hold3767/X _12760_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12761_/X sky130_fd_sc_hd__mux2_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14500_ hold636/X _14487_/B _14499_/X _14552_/C1 vssd1 vssd1 vccd1 vccd1 hold637/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _12093_/A _11712_/B vssd1 vssd1 vccd1 vccd1 _11712_/X sky130_fd_sc_hd__or2_1
X_15480_ _15480_/A _15480_/B _15480_/C _15480_/D vssd1 vssd1 vccd1 vccd1 _15480_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_167_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ hold3383/X _12691_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12692_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14431_ _15165_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _14431_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11643_ _11649_/A _11643_/B vssd1 vssd1 vccd1 vccd1 _11643_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17150_ _17278_/CLK _17150_/D vssd1 vssd1 vccd1 vccd1 _17150_/Q sky130_fd_sc_hd__dfxtp_1
X_14362_ _14362_/A _14362_/B vssd1 vssd1 vccd1 vccd1 _17980_/D sky130_fd_sc_hd__and2_1
XFILLER_0_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11574_ _11670_/A _11574_/B vssd1 vssd1 vccd1 vccd1 _11574_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput17 input17/A vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_2
Xinput28 input28/A vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_6
X_16101_ _16125_/CLK _16101_/D vssd1 vssd1 vccd1 vccd1 hold737/A sky130_fd_sc_hd__dfxtp_1
X_10525_ hold3261/X _10619_/B _10524_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10525_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput39 input39/A vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_1
X_13313_ hold2041/X hold4676/X _13409_/S vssd1 vssd1 vccd1 vccd1 _13314_/B sky130_fd_sc_hd__mux2_1
X_14293_ hold1682/X _14333_/A2 _14292_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _14293_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17081_ _17865_/CLK _17081_/D vssd1 vssd1 vccd1 vccd1 _17081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16032_ _17284_/CLK _16032_/D vssd1 vssd1 vccd1 vccd1 hold461/A sky130_fd_sc_hd__dfxtp_1
X_13244_ hold3450/X _13243_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13244_/X sky130_fd_sc_hd__mux2_4
X_10456_ hold4602/X _10646_/B _10455_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _10456_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ _13199_/A1 _13173_/X _13174_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13175_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10387_ hold3282/X _10601_/B _10386_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10387_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12126_ _12285_/A _12126_/B vssd1 vssd1 vccd1 vccd1 _12126_/X sky130_fd_sc_hd__or2_1
XFILLER_0_241_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17983_ _17983_/CLK _17983_/D vssd1 vssd1 vccd1 vccd1 _17983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_236_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12057_ _13749_/A _12057_/B vssd1 vssd1 vccd1 vccd1 _12057_/X sky130_fd_sc_hd__or2_1
X_16934_ _17877_/CLK _16934_/D vssd1 vssd1 vccd1 vccd1 _16934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11008_ hold4991/X _11213_/B _11007_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _11008_/X
+ sky130_fd_sc_hd__o211a_1
X_16865_ _18070_/CLK _16865_/D vssd1 vssd1 vccd1 vccd1 _16865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15816_ _17729_/CLK _15816_/D vssd1 vssd1 vccd1 vccd1 _15816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16796_ _18031_/CLK _16796_/D vssd1 vssd1 vccd1 vccd1 _16796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_463_wb_clk_i clkbuf_6_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17435_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15747_ _17718_/CLK _15747_/D vssd1 vssd1 vccd1 vccd1 _15747_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ hold3239/X _12958_/X _12971_/S vssd1 vssd1 vccd1 vccd1 _12960_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15678_ _17209_/CLK _15678_/D vssd1 vssd1 vccd1 vccd1 _15678_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17417_ _17429_/CLK _17417_/D vssd1 vssd1 vccd1 vccd1 _17417_/Q sky130_fd_sc_hd__dfxtp_1
X_14629_ hold1905/X _14664_/B _14628_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _14629_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18397_ _18399_/CLK _18397_/D vssd1 vssd1 vccd1 vccd1 _18397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08150_ _14960_/A hold1079/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08150_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17348_ _18400_/CLK _17348_/D vssd1 vssd1 vccd1 vccd1 _17348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08081_ hold1544/X _08097_/A2 _08080_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _08081_/X
+ sky130_fd_sc_hd__o211a_1
X_17279_ _17279_/CLK _17279_/D vssd1 vssd1 vccd1 vccd1 _17279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4105 _16935_/Q vssd1 vssd1 vccd1 vccd1 hold4105/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4116 _11515_/X vssd1 vssd1 vccd1 vccd1 _16995_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4127 _16778_/Q vssd1 vssd1 vccd1 vccd1 hold4127/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4138 _16784_/Q vssd1 vssd1 vccd1 vccd1 hold4138/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3404 _16354_/Q vssd1 vssd1 vccd1 vccd1 _13302_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold4149 _17017_/Q vssd1 vssd1 vccd1 vccd1 hold4149/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3415 _10008_/Y vssd1 vssd1 vccd1 vccd1 _10009_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3426 _10026_/Y vssd1 vssd1 vccd1 vccd1 _10027_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3437 _10582_/Y vssd1 vssd1 vccd1 vccd1 _16684_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08983_ hold143/X hold145/X _08991_/S vssd1 vssd1 vccd1 vccd1 _08984_/B sky130_fd_sc_hd__mux2_1
Xhold3448 _09990_/Y vssd1 vssd1 vccd1 vccd1 _09991_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2703 _15599_/Q vssd1 vssd1 vccd1 vccd1 hold2703/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2714 _15583_/Q vssd1 vssd1 vccd1 vccd1 hold2714/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3459 _16544_/Q vssd1 vssd1 vccd1 vccd1 hold3459/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2725 _17842_/Q vssd1 vssd1 vccd1 vccd1 hold2725/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2736 _14863_/X vssd1 vssd1 vccd1 vccd1 _18220_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07934_ _15557_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07934_/X sky130_fd_sc_hd__or2_1
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2747 _16212_/Q vssd1 vssd1 vccd1 vccd1 hold2747/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2758 _15733_/Q vssd1 vssd1 vccd1 vccd1 hold2758/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2769 _16159_/Q vssd1 vssd1 vccd1 vccd1 hold2769/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07865_ _15163_/A _07865_/B vssd1 vssd1 vccd1 vccd1 _07865_/Y sky130_fd_sc_hd__nand2_1
X_09604_ hold4833/X _09992_/B _09603_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _09604_/X
+ sky130_fd_sc_hd__o211a_1
X_07796_ _11158_/A _07796_/B vssd1 vssd1 vccd1 vccd1 _18462_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09535_ hold3218/X _10004_/B _09534_/X _15048_/A vssd1 vssd1 vccd1 vccd1 _09535_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_133_wb_clk_i clkbuf_6_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17325_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09466_ _09472_/C _09472_/D _09478_/B vssd1 vssd1 vccd1 vccd1 _09466_/Y sky130_fd_sc_hd__o21ai_1
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08417_ _15531_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08417_/X sky130_fd_sc_hd__or2_1
X_09397_ hold5950/A _09342_/B _09342_/Y _09396_/X _12412_/A vssd1 vssd1 vccd1 vccd1
+ _09397_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_171_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08348_ _14457_/A hold2340/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08349_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_62_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08279_ hold1267/X _08268_/B _08278_/X _12753_/A vssd1 vssd1 vccd1 vccd1 _08279_/X
+ sky130_fd_sc_hd__o211a_1
Xhold6030 _17556_/Q vssd1 vssd1 vccd1 vccd1 hold6030/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6041 data_in[13] vssd1 vssd1 vccd1 vccd1 hold166/A sky130_fd_sc_hd__dlygate4sd3_1
X_10310_ hold1058/X hold3670/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10311_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_105_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6052 _18369_/Q vssd1 vssd1 vccd1 vccd1 hold6052/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11290_ hold5213/X _11789_/B _11289_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _11290_/X
+ sky130_fd_sc_hd__o211a_1
Xhold6063 _18394_/Q vssd1 vssd1 vccd1 vccd1 hold6063/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6074 _18073_/Q vssd1 vssd1 vccd1 vccd1 hold6074/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6085 _18459_/Q vssd1 vssd1 vccd1 vccd1 hold6085/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5340 _11020_/X vssd1 vssd1 vccd1 vccd1 _16830_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold6096 data_in[4] vssd1 vssd1 vccd1 vccd1 hold257/A sky130_fd_sc_hd__dlygate4sd3_1
X_10241_ hold2637/X hold3700/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10242_/B sky130_fd_sc_hd__mux2_1
Xhold5351 _17647_/Q vssd1 vssd1 vccd1 vccd1 hold5351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5362 _17012_/Q vssd1 vssd1 vccd1 vccd1 hold5362/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5373 _10735_/X vssd1 vssd1 vccd1 vccd1 _16735_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5384 _17269_/Q vssd1 vssd1 vccd1 vccd1 hold5384/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4650 _16458_/Q vssd1 vssd1 vccd1 vccd1 hold4650/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5395 _13492_/X vssd1 vssd1 vccd1 vccd1 _17617_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10172_ hold959/X hold3595/X _10634_/C vssd1 vssd1 vccd1 vccd1 _10173_/B sky130_fd_sc_hd__mux2_1
Xhold4661 _13618_/X vssd1 vssd1 vccd1 vccd1 _17659_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4672 _17601_/Q vssd1 vssd1 vccd1 vccd1 hold4672/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4683 _17664_/Q vssd1 vssd1 vccd1 vccd1 hold4683/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4694 _09712_/X vssd1 vssd1 vccd1 vccd1 _16394_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3960 _16759_/Q vssd1 vssd1 vccd1 vccd1 hold3960/X sky130_fd_sc_hd__dlygate4sd3_1
X_14980_ _14980_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14980_/X sky130_fd_sc_hd__or2_1
Xhold3971 _10393_/X vssd1 vssd1 vccd1 vccd1 _16621_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3982 _16418_/Q vssd1 vssd1 vccd1 vccd1 hold3982/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout150 _12626_/S vssd1 vssd1 vccd1 vccd1 _12749_/S sky130_fd_sc_hd__buf_4
Xhold3993 _16443_/Q vssd1 vssd1 vccd1 vccd1 hold3993/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_156_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout161 _13817_/B vssd1 vssd1 vccd1 vccd1 _13814_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_233_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout172 _11717_/B vssd1 vssd1 vccd1 vccd1 _12299_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_199_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout183 fanout210/X vssd1 vssd1 vccd1 vccd1 _11071_/A2 sky130_fd_sc_hd__clkbuf_4
X_13931_ _13931_/A hold309/X vssd1 vssd1 vccd1 vccd1 _17773_/D sky130_fd_sc_hd__and2_1
Xfanout194 fanout210/X vssd1 vssd1 vccd1 vccd1 _13877_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_233_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16650_ _18063_/CLK _16650_/D vssd1 vssd1 vccd1 vccd1 _16650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13862_ _13862_/A _13862_/B _13862_/C vssd1 vssd1 vccd1 vccd1 _13862_/X sky130_fd_sc_hd__and3_1
XFILLER_0_57_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15601_ _17279_/CLK _15601_/D vssd1 vssd1 vccd1 vccd1 _15601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12813_ _12837_/A _12813_/B vssd1 vssd1 vccd1 vccd1 _17447_/D sky130_fd_sc_hd__and2_1
XFILLER_0_241_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_232_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16581_ _18177_/CLK _16581_/D vssd1 vssd1 vccd1 vccd1 _16581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13793_ hold1291/X hold4658/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13794_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_69_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18320_ _18352_/CLK hold291/X vssd1 vssd1 vccd1 vccd1 _18320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15532_ hold1453/X _15547_/B _15531_/X _12822_/A vssd1 vssd1 vccd1 vccd1 _15532_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_1302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _12750_/A _12744_/B vssd1 vssd1 vccd1 vccd1 _17424_/D sky130_fd_sc_hd__and2_1
XFILLER_0_201_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18251_ _18383_/CLK _18251_/D vssd1 vssd1 vccd1 vccd1 _18251_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15463_ _15481_/A1 _15455_/X _15462_/X _15490_/B1 hold5957/A vssd1 vssd1 vccd1 vccd1
+ _15463_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_166_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _12873_/A _12675_/B vssd1 vssd1 vccd1 vccd1 _17401_/D sky130_fd_sc_hd__and2_1
XFILLER_0_182_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17202_ _17202_/CLK _17202_/D vssd1 vssd1 vccd1 vccd1 _17202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14414_ hold2973/X _14446_/A2 _14413_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _14414_/X
+ sky130_fd_sc_hd__o211a_1
X_18182_ _18214_/CLK _18182_/D vssd1 vssd1 vccd1 vccd1 _18182_/Q sky130_fd_sc_hd__dfxtp_1
X_11626_ hold5651/X _12299_/B _11625_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _11626_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_182_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15394_ _15394_/A _15394_/B vssd1 vssd1 vccd1 vccd1 _18415_/D sky130_fd_sc_hd__and2_1
XFILLER_0_65_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17133_ _17261_/CLK _17133_/D vssd1 vssd1 vccd1 vccd1 _17133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14345_ hold911/X _17972_/Q _14391_/S vssd1 vssd1 vccd1 vccd1 _14345_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11557_ hold5253/X _11165_/B _11556_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _11557_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold609 hold609/A vssd1 vssd1 vccd1 vccd1 hold609/X sky130_fd_sc_hd__dlygate4sd3_1
X_10508_ hold1089/X hold3642/X _10646_/C vssd1 vssd1 vccd1 vccd1 _10509_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17064_ _18448_/CLK _17064_/D vssd1 vssd1 vccd1 vccd1 _17064_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_28_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_28_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_150_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14276_ _14330_/A _14282_/B vssd1 vssd1 vccd1 vccd1 _14276_/X sky130_fd_sc_hd__or2_1
X_11488_ hold5271/X _11786_/B _11487_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _11488_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_204_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16015_ _18424_/CLK _16015_/D vssd1 vssd1 vccd1 vccd1 hold565/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10439_ hold2888/X _16637_/Q _10637_/C vssd1 vssd1 vccd1 vccd1 _10440_/B sky130_fd_sc_hd__mux2_1
X_13227_ _13226_/X hold4717/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13227_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_141_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13158_ _13158_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13158_/X sky130_fd_sc_hd__or2_1
XFILLER_0_236_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ hold5681/X _12299_/B _12108_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _12109_/X
+ sky130_fd_sc_hd__o211a_1
X_13089_ _13089_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13089_/X sky130_fd_sc_hd__and2_1
XFILLER_0_178_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17966_ _18345_/CLK _17966_/D vssd1 vssd1 vccd1 vccd1 _17966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1309 _16278_/Q vssd1 vssd1 vccd1 vccd1 hold1309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_236_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16917_ _17831_/CLK _16917_/D vssd1 vssd1 vccd1 vccd1 _16917_/Q sky130_fd_sc_hd__dfxtp_1
X_17897_ _17897_/CLK _17897_/D vssd1 vssd1 vccd1 vccd1 _17897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_1371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16848_ _18051_/CLK _16848_/D vssd1 vssd1 vccd1 vccd1 _16848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_233_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16779_ _18047_/CLK _16779_/D vssd1 vssd1 vccd1 vccd1 _16779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09320_ hold3029/X _09323_/B _09319_/Y _12894_/A vssd1 vssd1 vccd1 vccd1 _09320_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09251_ hold951/X _16237_/Q _09283_/S vssd1 vssd1 vccd1 vccd1 hold952/A sky130_fd_sc_hd__mux2_1
XFILLER_0_8_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18449_ _18451_/CLK _18449_/D vssd1 vssd1 vccd1 vccd1 _18449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08202_ hold2017/X _08213_/B _08201_/X _13765_/C1 vssd1 vssd1 vccd1 vccd1 _08202_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09182_ _15511_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09182_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08133_ _08133_/A _08133_/B vssd1 vssd1 vccd1 vccd1 _15705_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08064_ hold933/X _08094_/B vssd1 vssd1 vccd1 vccd1 _08064_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3201 _10620_/Y vssd1 vssd1 vccd1 vccd1 _10621_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3212 _17498_/Q vssd1 vssd1 vccd1 vccd1 hold3212/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3223 _12971_/X vssd1 vssd1 vccd1 vccd1 _12972_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3234 _09925_/X vssd1 vssd1 vccd1 vccd1 _16465_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3245 _16377_/Q vssd1 vssd1 vccd1 vccd1 hold3245/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2500 _08330_/X vssd1 vssd1 vccd1 vccd1 _15798_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3256 _10540_/X vssd1 vssd1 vccd1 vccd1 _16670_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2511 _17992_/Q vssd1 vssd1 vccd1 vccd1 hold2511/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2522 _18189_/Q vssd1 vssd1 vccd1 vccd1 hold2522/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3267 _09877_/X vssd1 vssd1 vccd1 vccd1 _16449_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08966_ _15482_/A hold348/X vssd1 vssd1 vccd1 vccd1 _16100_/D sky130_fd_sc_hd__and2_1
Xhold2533 _13969_/X vssd1 vssd1 vccd1 vccd1 _17791_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3278 _16513_/Q vssd1 vssd1 vccd1 vccd1 _10067_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2544 _18177_/Q vssd1 vssd1 vccd1 vccd1 hold2544/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3289 _12866_/X vssd1 vssd1 vccd1 vccd1 _12867_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_385_wb_clk_i clkbuf_6_35_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17209_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1810 _13991_/X vssd1 vssd1 vccd1 vccd1 _17802_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2555 _17852_/Q vssd1 vssd1 vccd1 vccd1 hold2555/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1821 _18385_/Q vssd1 vssd1 vccd1 vccd1 hold1821/X sky130_fd_sc_hd__dlygate4sd3_1
X_07917_ hold1678/X _07918_/B _07916_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _07917_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2566 _15544_/X vssd1 vssd1 vccd1 vccd1 _18450_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1832 _07935_/X vssd1 vssd1 vccd1 vccd1 _15611_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2577 _17837_/Q vssd1 vssd1 vccd1 vccd1 hold2577/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2588 _14719_/X vssd1 vssd1 vccd1 vccd1 _18151_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08897_ _12416_/A hold562/X vssd1 vssd1 vccd1 vccd1 _16066_/D sky130_fd_sc_hd__and2_1
Xhold1843 _18010_/Q vssd1 vssd1 vccd1 vccd1 hold1843/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1854 _14919_/X vssd1 vssd1 vccd1 vccd1 _18246_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2599 _15604_/Q vssd1 vssd1 vccd1 vccd1 hold2599/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_314_wb_clk_i clkbuf_6_47_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18069_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1865 _15576_/Q vssd1 vssd1 vccd1 vccd1 hold1865/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1876 _14317_/X vssd1 vssd1 vccd1 vccd1 _17958_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07848_ hold3116/X _07869_/B _07847_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _07848_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1887 _15561_/Q vssd1 vssd1 vccd1 vccd1 hold1887/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1898 _14418_/X vssd1 vssd1 vccd1 vccd1 _18007_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09518_ hold2497/X _13110_/A _09992_/C vssd1 vssd1 vccd1 vccd1 _09519_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10790_ hold1501/X hold4016/X _11210_/C vssd1 vssd1 vccd1 vccd1 _10791_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_211_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09456_/D _09449_/B vssd1 vssd1 vccd1 vccd1 _16309_/D sky130_fd_sc_hd__nor2_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12460_ _17323_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12460_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ hold2205/X _16961_/Q _11774_/C vssd1 vssd1 vccd1 vccd1 _11412_/B sky130_fd_sc_hd__mux2_1
X_12391_ hold147/X _17289_/Q _12443_/S vssd1 vssd1 vccd1 vccd1 hold395/A sky130_fd_sc_hd__mux2_1
XFILLER_0_191_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14130_ _15203_/A _14140_/B vssd1 vssd1 vccd1 vccd1 _14130_/X sky130_fd_sc_hd__or2_1
X_11342_ hold1656/X hold5434/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11343_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_201_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_wb_clk_i clkbuf_6_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18013_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14061_ hold2989/X _14094_/B _14060_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _14061_/X
+ sky130_fd_sc_hd__o211a_1
X_11273_ hold2256/X hold4751/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11274_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5170 _13702_/X vssd1 vssd1 vccd1 vccd1 _17687_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10224_ _10536_/A _10224_/B vssd1 vssd1 vccd1 vccd1 _10224_/X sky130_fd_sc_hd__or2_1
Xhold5181 _16757_/Q vssd1 vssd1 vccd1 vccd1 hold5181/X sky130_fd_sc_hd__dlygate4sd3_1
X_13012_ hold2404/X _13003_/Y _13011_/X _14358_/A vssd1 vssd1 vccd1 vccd1 _13012_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5192 _11347_/X vssd1 vssd1 vccd1 vccd1 _16939_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4480 _17213_/Q vssd1 vssd1 vccd1 vccd1 hold4480/X sky130_fd_sc_hd__dlygate4sd3_1
X_17820_ _17820_/CLK _17820_/D vssd1 vssd1 vccd1 vccd1 _17820_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10155_ _10515_/A _10155_/B vssd1 vssd1 vccd1 vccd1 _10155_/X sky130_fd_sc_hd__or2_1
Xhold4491 _17138_/Q vssd1 vssd1 vccd1 vccd1 hold4491/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17751_ _18460_/CLK _17751_/D vssd1 vssd1 vccd1 vccd1 _17751_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3790 _11785_/Y vssd1 vssd1 vccd1 vccd1 _17085_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14963_ hold6066/X _14946_/B hold408/X _15228_/C1 vssd1 vssd1 vccd1 vccd1 hold409/A
+ sky130_fd_sc_hd__o211a_1
X_10086_ _10476_/A _10086_/B vssd1 vssd1 vccd1 vccd1 _10086_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16702_ _18164_/CLK _16702_/D vssd1 vssd1 vccd1 vccd1 _16702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13914_ _15203_/A _17765_/Q hold297/X vssd1 vssd1 vccd1 vccd1 _13914_/X sky130_fd_sc_hd__mux2_1
X_17682_ _17705_/CLK _17682_/D vssd1 vssd1 vccd1 vccd1 _17682_/Q sky130_fd_sc_hd__dfxtp_1
X_14894_ _15233_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14894_/X sky130_fd_sc_hd__or2_1
X_16633_ _18191_/CLK _16633_/D vssd1 vssd1 vccd1 vccd1 _16633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13845_ hold4303/X _13407_/A _13844_/X vssd1 vssd1 vccd1 vccd1 _13845_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_202_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16564_ _18154_/CLK _16564_/D vssd1 vssd1 vccd1 vccd1 _16564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13776_ _13776_/A _13776_/B vssd1 vssd1 vccd1 vccd1 _13776_/X sky130_fd_sc_hd__or2_1
X_10988_ hold2066/X _16820_/Q _11186_/C vssd1 vssd1 vccd1 vccd1 _10989_/B sky130_fd_sc_hd__mux2_1
X_18303_ _18411_/CLK hold369/X vssd1 vssd1 vccd1 vccd1 _18303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15515_ _15515_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15515_/X sky130_fd_sc_hd__or2_1
X_12727_ hold2459/X hold3165/X _12766_/S vssd1 vssd1 vccd1 vccd1 _12727_/X sky130_fd_sc_hd__mux2_1
X_16495_ _18250_/CLK _16495_/D vssd1 vssd1 vccd1 vccd1 _16495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18234_ _18234_/CLK _18234_/D vssd1 vssd1 vccd1 vccd1 _18234_/Q sky130_fd_sc_hd__dfxtp_1
X_15446_ _17320_/Q _15487_/A2 _15446_/B1 hold399/X vssd1 vssd1 vccd1 vccd1 _15446_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_182_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12658_ hold2201/X hold3133/X _12850_/S vssd1 vssd1 vccd1 vccd1 _12658_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18165_ _18215_/CLK _18165_/D vssd1 vssd1 vccd1 vccd1 _18165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11609_ hold3039/X _17027_/Q _11774_/C vssd1 vssd1 vccd1 vccd1 _11610_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15377_ hold545/X _09357_/A _09386_/D hold659/X _15376_/X vssd1 vssd1 vccd1 vccd1
+ _15382_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12589_ hold2495/X hold3118/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12589_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_142_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17116_ _17614_/CLK _17116_/D vssd1 vssd1 vccd1 vccd1 _17116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14328_ _14543_/A _14334_/B vssd1 vssd1 vccd1 vccd1 _14328_/X sky130_fd_sc_hd__or2_1
X_18096_ _18180_/CLK _18096_/D vssd1 vssd1 vccd1 vccd1 _18096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold406 hold406/A vssd1 vssd1 vccd1 vccd1 hold406/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold417 hold422/X vssd1 vssd1 vccd1 vccd1 hold423/A sky130_fd_sc_hd__buf_6
Xhold428 hold52/X vssd1 vssd1 vccd1 vccd1 input19/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold439 hold439/A vssd1 vssd1 vccd1 vccd1 hold439/X sky130_fd_sc_hd__dlygate4sd3_1
X_17047_ _17895_/CLK _17047_/D vssd1 vssd1 vccd1 vccd1 _17047_/Q sky130_fd_sc_hd__dfxtp_1
X_14259_ hold2623/X _14268_/B _14258_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14259_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout908 hold289/X vssd1 vssd1 vccd1 vccd1 _14443_/A sky130_fd_sc_hd__buf_6
Xfanout919 hold991/X vssd1 vssd1 vccd1 vccd1 _15225_/A sky130_fd_sc_hd__buf_6
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ hold452/X hold844/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08821_/B sky130_fd_sc_hd__mux2_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 hold1153/X vssd1 vssd1 vccd1 vccd1 hold1106/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 _17915_/Q vssd1 vssd1 vccd1 vccd1 hold1117/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ hold23/X hold325/X _08779_/S vssd1 vssd1 vccd1 vccd1 _08752_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_174_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1128 _14544_/X vssd1 vssd1 vccd1 vccd1 _18068_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17949_ _17949_/CLK hold538/X vssd1 vssd1 vccd1 vccd1 hold537/A sky130_fd_sc_hd__dfxtp_1
Xhold1139 _15173_/X vssd1 vssd1 vccd1 vccd1 hold1139/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08682_ _15491_/A _08682_/B vssd1 vssd1 vccd1 vccd1 _15962_/D sky130_fd_sc_hd__and2_1
XFILLER_0_174_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09303_ _15199_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09303_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09234_ _12843_/A _09234_/B vssd1 vssd1 vccd1 vccd1 _16228_/D sky130_fd_sc_hd__and2_1
XFILLER_0_145_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_228_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09165_ hold2464/X _09164_/B _09164_/Y _12906_/A vssd1 vssd1 vccd1 vccd1 _09165_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08116_ _14461_/A hold2787/X hold108/X vssd1 vssd1 vccd1 vccd1 _08117_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_185_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09096_ _15103_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _09096_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08047_ hold444/X hold405/X hold337/X hold509/X vssd1 vssd1 vccd1 vccd1 _14627_/A
+ sky130_fd_sc_hd__or4bb_4
Xhold940 hold940/A vssd1 vssd1 vccd1 vccd1 hold940/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold951 hold951/A vssd1 vssd1 vccd1 vccd1 hold951/X sky130_fd_sc_hd__buf_12
Xhold962 hold962/A vssd1 vssd1 vccd1 vccd1 hold962/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 hold973/A vssd1 vssd1 vccd1 vccd1 hold973/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold984 hold984/A vssd1 vssd1 vccd1 vccd1 hold984/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3020 _14516_/X vssd1 vssd1 vccd1 vccd1 _18054_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 hold995/A vssd1 vssd1 vccd1 vccd1 hold995/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3031 _18012_/Q vssd1 vssd1 vccd1 vccd1 hold3031/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3042 _07945_/X vssd1 vssd1 vccd1 vccd1 _15615_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3053 _15629_/Q vssd1 vssd1 vccd1 vccd1 hold3053/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09998_ _16490_/Q _11162_/B _11162_/C vssd1 vssd1 vccd1 vccd1 _09998_/X sky130_fd_sc_hd__and3_1
Xhold3064 _13953_/X vssd1 vssd1 vccd1 vccd1 _17783_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2330 _16250_/Q vssd1 vssd1 vccd1 vccd1 hold2330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3075 _07903_/X vssd1 vssd1 vccd1 vccd1 _15595_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3086 _13048_/X vssd1 vssd1 vccd1 vccd1 _17525_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2341 _15780_/Q vssd1 vssd1 vccd1 vccd1 hold2341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3097 _18115_/Q vssd1 vssd1 vccd1 vccd1 hold3097/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2352 _14667_/X vssd1 vssd1 vccd1 vccd1 _18126_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08949_ hold679/X hold882/X _08991_/S vssd1 vssd1 vccd1 vccd1 hold883/A sky130_fd_sc_hd__mux2_1
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2363 _17800_/Q vssd1 vssd1 vccd1 vccd1 hold2363/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2374 _08016_/X vssd1 vssd1 vccd1 vccd1 _15649_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1640 _09119_/X vssd1 vssd1 vccd1 vccd1 _16174_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2385 _14119_/X vssd1 vssd1 vccd1 vccd1 _17863_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1651 _07969_/X vssd1 vssd1 vccd1 vccd1 _15627_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2396 _15651_/Q vssd1 vssd1 vccd1 vccd1 hold2396/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1662 _17964_/Q vssd1 vssd1 vccd1 vccd1 hold1662/X sky130_fd_sc_hd__dlygate4sd3_1
X_11960_ hold2359/X hold3976/X _13748_/S vssd1 vssd1 vccd1 vccd1 _11961_/B sky130_fd_sc_hd__mux2_1
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1673 _08224_/X vssd1 vssd1 vccd1 vccd1 _15748_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_230_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1684 _18061_/Q vssd1 vssd1 vccd1 vccd1 hold1684/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_233_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911_ _11103_/A _10911_/B vssd1 vssd1 vccd1 vccd1 _10911_/X sky130_fd_sc_hd__or2_1
Xhold1695 _08231_/X vssd1 vssd1 vccd1 vccd1 _15750_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ hold2654/X hold3505/X _12371_/C vssd1 vssd1 vccd1 vccd1 _11892_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_211_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13630_ hold4589/X _13829_/B _13629_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13630_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_212_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10842_ _11124_/A _10842_/B vssd1 vssd1 vccd1 vccd1 _10842_/X sky130_fd_sc_hd__or2_1
XFILLER_0_184_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13561_ hold5355/X _13868_/B _13560_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _13561_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10773_ _11061_/A _10773_/B vssd1 vssd1 vccd1 vccd1 _10773_/X sky130_fd_sc_hd__or2_1
X_15300_ hold470/X _15448_/A2 _15446_/B1 hold285/X vssd1 vssd1 vccd1 vccd1 _15300_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12512_ _09342_/A hold2264/X _07802_/Y _12511_/X vssd1 vssd1 vccd1 vccd1 _12512_/X
+ sky130_fd_sc_hd__o211a_1
X_16280_ _17750_/CLK _16280_/D vssd1 vssd1 vccd1 vccd1 _16280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13492_ hold5394/X _13883_/B _13491_/X _13684_/C1 vssd1 vssd1 vccd1 vccd1 _13492_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15231_ _15231_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15231_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12443_ hold278/X _17315_/Q _12443_/S vssd1 vssd1 vccd1 vccd1 hold279/A sky130_fd_sc_hd__mux2_1
XFILLER_0_191_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15162_ hold1503/X _15165_/B _15161_/Y _15212_/C1 vssd1 vssd1 vccd1 vccd1 _15162_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12374_ _17282_/Q _12374_/B _13748_/S vssd1 vssd1 vccd1 vccd1 _12374_/X sky130_fd_sc_hd__and3_1
XFILLER_0_205_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14113_ hold2117/X _14142_/B _14112_/X _14462_/C1 vssd1 vssd1 vccd1 vccd1 _14113_/X
+ sky130_fd_sc_hd__o211a_1
X_11325_ _12093_/A _11325_/B vssd1 vssd1 vccd1 vccd1 _11325_/X sky130_fd_sc_hd__or2_1
X_15093_ _15201_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15093_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14044_ _14330_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14044_/X sky130_fd_sc_hd__or2_1
X_11256_ _11649_/A _11256_/B vssd1 vssd1 vccd1 vccd1 _11256_/X sky130_fd_sc_hd__or2_1
XFILLER_0_205_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_236_wb_clk_i clkbuf_6_62_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18212_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ hold3320/X _10589_/B _10206_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10207_/X
+ sky130_fd_sc_hd__o211a_1
X_11187_ hold4318/X _11091_/A _11186_/X vssd1 vssd1 vccd1 vccd1 _11187_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10138_ hold5142/X _11225_/B _10137_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _10138_/X
+ sky130_fd_sc_hd__o211a_1
X_17803_ _17887_/CLK _17803_/D vssd1 vssd1 vccd1 vccd1 _17803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15995_ _18409_/CLK _15995_/D vssd1 vssd1 vccd1 vccd1 hold779/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17734_ _17734_/CLK _17734_/D vssd1 vssd1 vccd1 vccd1 _17734_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14946_ _15215_/A _14946_/B vssd1 vssd1 vccd1 vccd1 _14946_/Y sky130_fd_sc_hd__nand2_1
X_10069_ _10603_/A _10069_/B vssd1 vssd1 vccd1 vccd1 _16513_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17665_ _17697_/CLK _17665_/D vssd1 vssd1 vccd1 vccd1 _17665_/Q sky130_fd_sc_hd__dfxtp_1
X_14877_ hold1863/X _14880_/B _14876_/Y _14877_/C1 vssd1 vssd1 vccd1 vccd1 _14877_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_230_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16616_ _18206_/CLK _16616_/D vssd1 vssd1 vccd1 vccd1 _16616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13828_ _13864_/A _13828_/B vssd1 vssd1 vccd1 vccd1 _13828_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_106_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_230_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17596_ _17628_/CLK _17596_/D vssd1 vssd1 vccd1 vccd1 _17596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16547_ _18181_/CLK _16547_/D vssd1 vssd1 vccd1 vccd1 _16547_/Q sky130_fd_sc_hd__dfxtp_1
X_13759_ hold5414/X _13883_/B _13758_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13759_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16478_ _18391_/CLK _16478_/D vssd1 vssd1 vccd1 vccd1 _16478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18217_ _18217_/CLK _18217_/D vssd1 vssd1 vccd1 vccd1 _18217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15429_ hold189/X _09386_/A _15427_/X vssd1 vssd1 vccd1 vccd1 _15432_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_170_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18148_ _18154_/CLK _18148_/D vssd1 vssd1 vccd1 vccd1 _18148_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5906 output97/X vssd1 vssd1 vccd1 vccd1 data_out[3] sky130_fd_sc_hd__buf_12
XFILLER_0_14_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5917 _18408_/Q vssd1 vssd1 vccd1 vccd1 hold5917/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 hold451/X vssd1 vssd1 vccd1 vccd1 hold452/A sky130_fd_sc_hd__buf_1
XFILLER_0_223_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5928 _18410_/Q vssd1 vssd1 vccd1 vccd1 hold5928/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 input15/X vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__buf_1
XFILLER_0_198_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5939 hold5939/A vssd1 vssd1 vccd1 vccd1 load_status[5] sky130_fd_sc_hd__buf_12
XFILLER_0_124_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold225 input5/X vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__dlygate4sd3_1
X_18079_ _18265_/CLK _18079_/D vssd1 vssd1 vccd1 vccd1 _18079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold236 hold236/A vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 hold247/A vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold258 hold70/X vssd1 vssd1 vccd1 vccd1 input31/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09921_ _09981_/A _09921_/B vssd1 vssd1 vccd1 vccd1 _09921_/X sky130_fd_sc_hd__or2_1
XFILLER_0_141_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold269 hold362/X vssd1 vssd1 vccd1 vccd1 hold363/A sky130_fd_sc_hd__buf_6
Xfanout705 _09047_/A vssd1 vssd1 vccd1 vccd1 _12438_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout716 _14368_/A vssd1 vssd1 vccd1 vccd1 _14552_/C1 sky130_fd_sc_hd__buf_4
X_09852_ _09912_/A _09852_/B vssd1 vssd1 vccd1 vccd1 _09852_/X sky130_fd_sc_hd__or2_1
Xfanout727 _12418_/A vssd1 vssd1 vccd1 vccd1 _12426_/A sky130_fd_sc_hd__buf_4
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout738 fanout739/X vssd1 vssd1 vccd1 vccd1 _09907_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_226_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout749 fanout843/X vssd1 vssd1 vccd1 vccd1 _13777_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08803_ _08868_/B _12380_/B _13046_/D vssd1 vssd1 vccd1 vccd1 _08858_/S sky130_fd_sc_hd__or3_4
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09783_ _11109_/A _09783_/B vssd1 vssd1 vccd1 vccd1 _09783_/X sky130_fd_sc_hd__or2_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08734_ _12426_/A hold855/X vssd1 vssd1 vccd1 vccd1 _15987_/D sky130_fd_sc_hd__and2_1
XFILLER_0_206_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 _15219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ hold226/X hold743/X _08721_/S vssd1 vssd1 vccd1 vccd1 hold744/A sky130_fd_sc_hd__mux2_1
XFILLER_0_230_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _17519_/Q hold937/X vssd1 vssd1 vccd1 vccd1 _13034_/D sky130_fd_sc_hd__and2_1
XFILLER_0_193_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09217_ hold2571/X _09218_/B _09216_/Y _12837_/A vssd1 vssd1 vccd1 vccd1 _09217_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09148_ _14596_/A _09156_/B vssd1 vssd1 vccd1 vccd1 _09148_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09079_ hold1163/X _09106_/B _09078_/X _12987_/A vssd1 vssd1 vccd1 vccd1 _09079_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11110_ hold5040/X _11204_/B _11109_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _11110_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12090_ _13407_/A _12090_/B vssd1 vssd1 vccd1 vccd1 _12090_/X sky130_fd_sc_hd__or2_1
XFILLER_0_202_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold770 hold770/A vssd1 vssd1 vccd1 vccd1 hold770/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 hold781/A vssd1 vssd1 vccd1 vccd1 hold781/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 hold792/A vssd1 vssd1 vccd1 vccd1 hold792/X sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ hold4861/X _11153_/B _11040_/X _14552_/C1 vssd1 vssd1 vccd1 vccd1 _11041_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2160 _09318_/X vssd1 vssd1 vccd1 vccd1 _16269_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2171 _18022_/Q vssd1 vssd1 vccd1 vccd1 hold2171/X sky130_fd_sc_hd__dlygate4sd3_1
X_14800_ _15193_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14800_/X sky130_fd_sc_hd__or2_1
XFILLER_0_216_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2182 _09157_/X vssd1 vssd1 vccd1 vccd1 _16191_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_232_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _17672_/CLK _15780_/D vssd1 vssd1 vccd1 vccd1 _15780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12992_ hold4770/X _12991_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12993_/B sky130_fd_sc_hd__mux2_1
Xhold2193 _16189_/Q vssd1 vssd1 vccd1 vccd1 hold2193/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1470 _18317_/Q vssd1 vssd1 vccd1 vccd1 hold1470/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14731_ hold1712/X _14718_/B _14730_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14731_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1481 _17814_/Q vssd1 vssd1 vccd1 vccd1 hold1481/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1492 _15178_/X vssd1 vssd1 vccd1 vccd1 _18372_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ _12267_/A _11943_/B vssd1 vssd1 vccd1 vccd1 _11943_/X sky130_fd_sc_hd__or2_1
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _17450_/CLK _17450_/D vssd1 vssd1 vccd1 vccd1 _17450_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _15163_/A _14666_/B vssd1 vssd1 vccd1 vccd1 _14662_/Y sky130_fd_sc_hd__nand2_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11874_ _13482_/A _11874_/B vssd1 vssd1 vccd1 vccd1 _11874_/X sky130_fd_sc_hd__or2_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16401_ _18323_/CLK _16401_/D vssd1 vssd1 vccd1 vccd1 _16401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13613_ hold2011/X hold3967/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13614_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_211_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17381_ _17484_/CLK _17381_/D vssd1 vssd1 vccd1 vccd1 _17381_/Q sky130_fd_sc_hd__dfxtp_1
X_10825_ hold5279/X _11195_/B _10824_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _10825_/X
+ sky130_fd_sc_hd__o211a_1
X_14593_ hold2737/X _14612_/B _14592_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _14593_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16332_ _18349_/CLK _16332_/D vssd1 vssd1 vccd1 vccd1 _16332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13544_ _15820_/Q _17635_/Q _13862_/C vssd1 vssd1 vccd1 vccd1 _13545_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_223_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10756_ hold4068/X _11732_/B _10755_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _10756_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16263_ _18013_/CLK _16263_/D vssd1 vssd1 vccd1 vccd1 _16263_/Q sky130_fd_sc_hd__dfxtp_1
X_13475_ hold1436/X hold5470/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13476_/B sky130_fd_sc_hd__mux2_1
X_10687_ hold5631/X _11165_/B _10686_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _10687_/X
+ sky130_fd_sc_hd__o211a_1
X_18002_ _18194_/CLK _18002_/D vssd1 vssd1 vccd1 vccd1 _18002_/Q sky130_fd_sc_hd__dfxtp_1
X_15214_ hold1949/X _15221_/B _15213_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _15214_/X
+ sky130_fd_sc_hd__o211a_1
X_12426_ _12426_/A _12426_/B vssd1 vssd1 vccd1 vccd1 _17306_/D sky130_fd_sc_hd__and2_1
X_16194_ _17477_/CLK _16194_/D vssd1 vssd1 vccd1 vccd1 _16194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_417_wb_clk_i clkbuf_6_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17259_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_106_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15145_ _15145_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15145_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12357_ hold4370/X _13482_/A _12356_/X vssd1 vssd1 vccd1 vccd1 _12357_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ hold4131/X _12329_/B _11307_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11308_/X
+ sky130_fd_sc_hd__o211a_1
X_15076_ hold1941/X hold341/X _15075_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _15076_/X
+ sky130_fd_sc_hd__o211a_1
X_12288_ _13314_/A _12288_/B vssd1 vssd1 vccd1 vccd1 _12288_/X sky130_fd_sc_hd__or2_1
XFILLER_0_205_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14027_ hold2960/X _14038_/B _14026_/X _13895_/A vssd1 vssd1 vccd1 vccd1 _14027_/X
+ sky130_fd_sc_hd__o211a_1
X_11239_ hold4105/X _11717_/B _11238_/X _12588_/A vssd1 vssd1 vccd1 vccd1 _11239_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_219_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15978_ _17297_/CLK _15978_/D vssd1 vssd1 vccd1 vccd1 hold174/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14929_ hold1960/X _14952_/B _14928_/X _15202_/C1 vssd1 vssd1 vccd1 vccd1 _14929_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17717_ _17746_/CLK _17717_/D vssd1 vssd1 vccd1 vccd1 _17717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08450_ _15509_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08450_/X sky130_fd_sc_hd__or2_1
X_17648_ _17648_/CLK _17648_/D vssd1 vssd1 vccd1 vccd1 _17648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_212_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08381_ _08381_/A _08381_/B vssd1 vssd1 vccd1 vccd1 _15822_/D sky130_fd_sc_hd__and2_1
X_17579_ _17606_/CLK _17579_/D vssd1 vssd1 vccd1 vccd1 _17579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09002_ hold618/X _16118_/Q _09056_/S vssd1 vssd1 vccd1 vccd1 hold619/A sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5703 _17031_/Q vssd1 vssd1 vccd1 vccd1 hold5703/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5714 _17114_/Q vssd1 vssd1 vccd1 vccd1 hold5714/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_158_wb_clk_i clkbuf_6_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16139_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5725 _13810_/Y vssd1 vssd1 vccd1 vccd1 _17723_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5736 _11881_/X vssd1 vssd1 vccd1 vccd1 _17117_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5747 _16334_/Q vssd1 vssd1 vccd1 vccd1 _13142_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5758 _11854_/X vssd1 vssd1 vccd1 vccd1 _17108_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5769 _17142_/Q vssd1 vssd1 vccd1 vccd1 hold5769/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout502 _10538_/S vssd1 vssd1 vccd1 vccd1 _10634_/C sky130_fd_sc_hd__clkbuf_8
X_09904_ hold4652/X _11201_/B _09903_/X _14372_/A vssd1 vssd1 vccd1 vccd1 _09904_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout513 _10385_/S vssd1 vssd1 vccd1 vccd1 _10049_/C sky130_fd_sc_hd__buf_6
XFILLER_0_217_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout524 _09315_/B vssd1 vssd1 vccd1 vccd1 _09337_/B sky130_fd_sc_hd__buf_4
Xfanout535 _09098_/B vssd1 vssd1 vccd1 vccd1 _09118_/B sky130_fd_sc_hd__buf_4
Xfanout546 _08393_/Y vssd1 vssd1 vccd1 vccd1 _08442_/A2 sky130_fd_sc_hd__buf_6
X_09835_ hold4606/X _10031_/B _09834_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09835_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout557 _08213_/B vssd1 vssd1 vccd1 vccd1 _08209_/B sky130_fd_sc_hd__buf_6
Xfanout568 _07991_/A2 vssd1 vssd1 vccd1 vccd1 _07978_/B sky130_fd_sc_hd__buf_6
Xfanout579 _14843_/B vssd1 vssd1 vccd1 vccd1 _15182_/B sky130_fd_sc_hd__buf_6
XFILLER_0_214_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_225_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09766_ hold4152/X _10052_/B _09765_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09766_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08717_ hold315/X hold869/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08718_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09697_ hold3601/X _10025_/B _09696_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _16389_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08648_ _15254_/A _08648_/B vssd1 vssd1 vccd1 vccd1 _15946_/D sky130_fd_sc_hd__and2_1
XFILLER_0_16_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08579_ _12390_/A hold621/X vssd1 vssd1 vccd1 vccd1 _15913_/D sky130_fd_sc_hd__and2_1
XFILLER_0_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _10610_/A _10628_/B _10628_/C vssd1 vssd1 vccd1 vccd1 _10610_/X sky130_fd_sc_hd__and3_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11590_ hold5661/X _12323_/B _11589_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _11590_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10541_ hold2620/X hold3890/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10542_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_187_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13260_ hold4399/X _13259_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13260_/X sky130_fd_sc_hd__mux2_2
X_10472_ hold2096/X _16648_/Q _10571_/C vssd1 vssd1 vccd1 vccd1 _10473_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12211_ hold5442/X _12299_/B _12210_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _12211_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13191_ _13199_/A1 _13189_/X _13190_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13191_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_1340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12142_ hold4563/X _12350_/B _12141_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _12142_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12073_ hold4480/X _12362_/B _12072_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _12073_/X
+ sky130_fd_sc_hd__o211a_1
X_16950_ _17936_/CLK _16950_/D vssd1 vssd1 vccd1 vccd1 _16950_/Q sky130_fd_sc_hd__dfxtp_1
X_15901_ _17322_/CLK _15901_/D vssd1 vssd1 vccd1 vccd1 hold281/A sky130_fd_sc_hd__dfxtp_1
X_11024_ hold1901/X hold5064/X _11216_/C vssd1 vssd1 vccd1 vccd1 _11025_/B sky130_fd_sc_hd__mux2_1
X_16881_ _18052_/CLK _16881_/D vssd1 vssd1 vccd1 vccd1 _16881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15832_ _17721_/CLK _15832_/D vssd1 vssd1 vccd1 vccd1 _15832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_218_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _17705_/CLK _15763_/D vssd1 vssd1 vccd1 vccd1 _15763_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _12978_/A _12975_/B vssd1 vssd1 vccd1 vccd1 _17501_/D sky130_fd_sc_hd__and2_1
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_234_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14714_ _15161_/A _14718_/B vssd1 vssd1 vccd1 vccd1 _14714_/Y sky130_fd_sc_hd__nand2_1
X_17502_ _17513_/CLK _17502_/D vssd1 vssd1 vccd1 vccd1 _17502_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ hold3935/X _13817_/B _11925_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _11926_/X
+ sky130_fd_sc_hd__o211a_1
X_15694_ _17262_/CLK _15694_/D vssd1 vssd1 vccd1 vccd1 _15694_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17433_ _17440_/CLK _17433_/D vssd1 vssd1 vccd1 vccd1 _17433_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14645_ hold3097/X _14664_/B _14644_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _14645_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11857_ hold5462/X _12335_/B _11856_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _11857_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_213_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10808_ hold2507/X _16760_/Q _11213_/C vssd1 vssd1 vccd1 vccd1 _10809_/B sky130_fd_sc_hd__mux2_1
X_17364_ _18013_/CLK _17364_/D vssd1 vssd1 vccd1 vccd1 _17364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14576_ hold915/X _14624_/B vssd1 vssd1 vccd1 vccd1 _14576_/X sky130_fd_sc_hd__or2_1
X_11788_ _12331_/A _11788_/B vssd1 vssd1 vccd1 vccd1 _11788_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_126_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16315_ _16315_/CLK _16315_/D vssd1 vssd1 vccd1 vccd1 _16315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13527_ _13719_/A _13527_/B vssd1 vssd1 vccd1 vccd1 _13527_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17295_ _17295_/CLK _17295_/D vssd1 vssd1 vccd1 vccd1 hold749/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10739_ hold2729/X hold3476/X _11219_/C vssd1 vssd1 vccd1 vccd1 _10740_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16246_ _17425_/CLK _16246_/D vssd1 vssd1 vccd1 vccd1 _16246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13458_ _13752_/A _13458_/B vssd1 vssd1 vccd1 vccd1 _13458_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_251_wb_clk_i clkbuf_6_59_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18218_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12409_ hold172/X hold781/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12410_/B sky130_fd_sc_hd__mux2_1
X_16177_ _17462_/CLK _16177_/D vssd1 vssd1 vccd1 vccd1 _16177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13389_ _13581_/A _13389_/B vssd1 vssd1 vccd1 vccd1 _13389_/X sky130_fd_sc_hd__or2_1
XFILLER_0_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput105 _17524_/Q vssd1 vssd1 vccd1 vccd1 io_out sky130_fd_sc_hd__buf_12
XFILLER_0_140_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput116 hold5952/X vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_12
Xhold4309 _16719_/Q vssd1 vssd1 vccd1 vccd1 hold4309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput127 hold5937/X vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_12
X_15128_ _15128_/A _15182_/B vssd1 vssd1 vccd1 vccd1 _15157_/B sky130_fd_sc_hd__or2_4
Xoutput138 hold5946/X vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_12
Xhold3608 _16617_/Q vssd1 vssd1 vccd1 vccd1 hold3608/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3619 _17438_/Q vssd1 vssd1 vccd1 vccd1 hold3619/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15059_ hold235/X _18315_/Q _15071_/S vssd1 vssd1 vccd1 vccd1 hold236/A sky130_fd_sc_hd__mux2_1
X_07950_ _15085_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07950_/X sky130_fd_sc_hd__or2_1
Xhold2907 _14781_/X vssd1 vssd1 vccd1 vccd1 _18181_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2918 _18119_/Q vssd1 vssd1 vccd1 vccd1 hold2918/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2929 _14809_/X vssd1 vssd1 vccd1 vccd1 _18194_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07881_ _15559_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07881_/X sky130_fd_sc_hd__or2_1
XFILLER_0_235_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_235_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09620_ hold1072/X _16364_/Q _10028_/C vssd1 vssd1 vccd1 vccd1 _09621_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_37_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09551_ hold1576/X _16341_/Q _10049_/C vssd1 vssd1 vccd1 vccd1 _09552_/B sky130_fd_sc_hd__mux2_1
X_08502_ hold444/X hold509/A hold337/X hold405/X vssd1 vssd1 vccd1 vccd1 _14897_/A
+ sky130_fd_sc_hd__or4bb_4
XFILLER_0_222_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09482_ _09483_/A _09482_/B vssd1 vssd1 vccd1 vccd1 _09484_/C sky130_fd_sc_hd__or2_1
XFILLER_0_176_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08433_ _15221_/A _08433_/B vssd1 vssd1 vccd1 vccd1 _08433_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_187_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08364_ _15533_/A hold2478/X hold115/X vssd1 vssd1 vccd1 vccd1 _08365_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_339_wb_clk_i clkbuf_6_43_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17280_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08295_ _15085_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08295_/X sky130_fd_sc_hd__or2_1
XFILLER_0_144_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5500 _16963_/Q vssd1 vssd1 vccd1 vccd1 hold5500/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5511 _16668_/Q vssd1 vssd1 vccd1 vccd1 hold5511/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5522 _13573_/X vssd1 vssd1 vccd1 vccd1 _17644_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5533 _17641_/Q vssd1 vssd1 vccd1 vccd1 hold5533/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5544 _12019_/X vssd1 vssd1 vccd1 vccd1 _17163_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5555 _17714_/Q vssd1 vssd1 vccd1 vccd1 hold5555/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4810 _12175_/X vssd1 vssd1 vccd1 vccd1 _17215_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4821 _16845_/Q vssd1 vssd1 vccd1 vccd1 hold4821/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5566 _11359_/X vssd1 vssd1 vccd1 vccd1 _16943_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4832 _13420_/X vssd1 vssd1 vccd1 vccd1 _17593_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5577 _17037_/Q vssd1 vssd1 vccd1 vccd1 hold5577/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5588 _13501_/X vssd1 vssd1 vccd1 vccd1 _17620_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4843 _17275_/Q vssd1 vssd1 vccd1 vccd1 hold4843/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4854 _10699_/X vssd1 vssd1 vccd1 vccd1 _16723_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5599 _16973_/Q vssd1 vssd1 vccd1 vccd1 hold5599/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4865 _17215_/Q vssd1 vssd1 vccd1 vccd1 hold4865/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4876 _11482_/X vssd1 vssd1 vccd1 vccd1 _16984_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout310 _11061_/A vssd1 vssd1 vccd1 vccd1 _09912_/A sky130_fd_sc_hd__buf_4
XFILLER_0_79_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout321 _10413_/A vssd1 vssd1 vccd1 vccd1 _10551_/A sky130_fd_sc_hd__buf_4
XFILLER_0_61_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4887 _16951_/Q vssd1 vssd1 vccd1 vccd1 hold4887/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout332 fanout335/A vssd1 vssd1 vccd1 vccd1 _10470_/A sky130_fd_sc_hd__buf_4
Xhold4898 _11092_/X vssd1 vssd1 vccd1 vccd1 _16854_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout343 _09369_/X vssd1 vssd1 vccd1 vccd1 _15474_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_233_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout354 _08721_/S vssd1 vssd1 vccd1 vccd1 _08727_/S sky130_fd_sc_hd__buf_8
Xfanout365 _15181_/Y vssd1 vssd1 vccd1 vccd1 _15219_/B sky130_fd_sc_hd__buf_6
XFILLER_0_226_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout376 hold446/X vssd1 vssd1 vccd1 vccd1 _15004_/B sky130_fd_sc_hd__buf_6
XFILLER_0_195_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout387 _14774_/B vssd1 vssd1 vccd1 vccd1 _14772_/B sky130_fd_sc_hd__buf_6
X_09818_ hold2220/X hold5821/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09819_/B sky130_fd_sc_hd__mux2_1
Xfanout398 _14479_/B vssd1 vssd1 vccd1 vccd1 _14499_/B sky130_fd_sc_hd__buf_8
XFILLER_0_94_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_55_wb_clk_i clkbuf_6_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18016_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_213_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09749_ _18320_/Q _16407_/Q _10385_/S vssd1 vssd1 vccd1 vccd1 _09750_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12760_ hold980/X _17431_/Q _12766_/S vssd1 vssd1 vccd1 vccd1 _12760_/X sky130_fd_sc_hd__mux2_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ hold1736/X hold5630/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11712_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_166_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12691_ hold1654/X _17408_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12691_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ hold2975/X _14433_/B _14429_/Y _14364_/A vssd1 vssd1 vccd1 vccd1 _14430_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11642_ hold1698/X hold5315/X _11738_/C vssd1 vssd1 vccd1 vccd1 _11643_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_181_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14361_ _14988_/A hold2593/X _14381_/S vssd1 vssd1 vccd1 vccd1 _14362_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11573_ hold2384/X hold5004/X _11765_/C vssd1 vssd1 vccd1 vccd1 _11574_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_181_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput18 input18/A vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_2
X_16100_ _18424_/CLK _16100_/D vssd1 vssd1 vccd1 vccd1 hold347/A sky130_fd_sc_hd__dfxtp_1
X_13312_ _13305_/X _13311_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17557_/D sky130_fd_sc_hd__o21a_1
Xinput29 input29/A vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_6
X_10524_ _10524_/A _10524_/B vssd1 vssd1 vccd1 vccd1 _10524_/X sky130_fd_sc_hd__or2_1
X_17080_ _17936_/CLK _17080_/D vssd1 vssd1 vccd1 vccd1 _17080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14292_ _14972_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14292_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_18_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_18_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_16031_ _18410_/CLK _16031_/D vssd1 vssd1 vccd1 vccd1 hold527/A sky130_fd_sc_hd__dfxtp_1
X_13243_ _13242_/X _16923_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13243_/X sky130_fd_sc_hd__mux2_2
X_10455_ _10551_/A _10455_/B vssd1 vssd1 vccd1 vccd1 _10455_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13174_ _13174_/A _13294_/B vssd1 vssd1 vccd1 vccd1 _13174_/X sky130_fd_sc_hd__or2_1
X_10386_ _10386_/A _10386_/B vssd1 vssd1 vccd1 vccd1 _10386_/X sky130_fd_sc_hd__or2_1
XFILLER_0_241_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12125_ hold2453/X _17199_/Q _12317_/C vssd1 vssd1 vccd1 vccd1 _12126_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17982_ _18047_/CLK _17982_/D vssd1 vssd1 vccd1 vccd1 _17982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12056_ hold969/X _17176_/Q _13748_/S vssd1 vssd1 vccd1 vccd1 _12057_/B sky130_fd_sc_hd__mux2_1
X_16933_ _18427_/CLK _16933_/D vssd1 vssd1 vccd1 vccd1 _16933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_237_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11007_ _11103_/A _11007_/B vssd1 vssd1 vccd1 vccd1 _11007_/X sky130_fd_sc_hd__or2_1
X_16864_ _18067_/CLK _16864_/D vssd1 vssd1 vccd1 vccd1 _16864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15815_ _17630_/CLK _15815_/D vssd1 vssd1 vccd1 vccd1 _15815_/Q sky130_fd_sc_hd__dfxtp_1
X_16795_ _18030_/CLK _16795_/D vssd1 vssd1 vccd1 vccd1 _16795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15746_ _17746_/CLK _15746_/D vssd1 vssd1 vccd1 vccd1 _15746_/Q sky130_fd_sc_hd__dfxtp_1
X_12958_ hold1446/X hold3232/X _12970_/S vssd1 vssd1 vccd1 vccd1 _12958_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11909_ hold2938/X _17127_/Q _12293_/C vssd1 vssd1 vccd1 vccd1 _11910_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15677_ _17902_/CLK _15677_/D vssd1 vssd1 vccd1 vccd1 _15677_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ hold2092/X _17474_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12889_/X sky130_fd_sc_hd__mux2_1
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_57_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_57_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_14628_ hold927/X _14678_/B vssd1 vssd1 vccd1 vccd1 _14628_/X sky130_fd_sc_hd__or2_1
XFILLER_0_135_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17416_ _17430_/CLK _17416_/D vssd1 vssd1 vccd1 vccd1 _17416_/Q sky130_fd_sc_hd__dfxtp_1
X_18396_ _18396_/CLK _18396_/D vssd1 vssd1 vccd1 vccd1 _18396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17347_ _17347_/CLK hold69/X vssd1 vssd1 vccd1 vccd1 _17347_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_432_wb_clk_i clkbuf_6_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17730_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14559_ hold927/X _14557_/Y _14558_/X _15218_/C1 vssd1 vssd1 vccd1 vccd1 hold928/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08080_ _14604_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08080_/X sky130_fd_sc_hd__or2_1
X_17278_ _17278_/CLK _17278_/D vssd1 vssd1 vccd1 vccd1 _17278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16229_ _17437_/CLK _16229_/D vssd1 vssd1 vccd1 vccd1 _16229_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4106 _11239_/X vssd1 vssd1 vccd1 vccd1 _16903_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4117 _16770_/Q vssd1 vssd1 vccd1 vccd1 hold4117/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4128 _10768_/X vssd1 vssd1 vccd1 vccd1 _16746_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4139 _10786_/X vssd1 vssd1 vccd1 vccd1 _16752_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3405 _10071_/Y vssd1 vssd1 vccd1 vccd1 _10072_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3416 _10009_/Y vssd1 vssd1 vccd1 vccd1 _16493_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3427 _10027_/Y vssd1 vssd1 vccd1 vccd1 _16499_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08982_ _12438_/A hold93/X vssd1 vssd1 vccd1 vccd1 _16108_/D sky130_fd_sc_hd__and2_1
Xhold3438 _16353_/Q vssd1 vssd1 vccd1 vccd1 _13294_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3449 _09991_/Y vssd1 vssd1 vccd1 vccd1 _16487_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2704 _07911_/X vssd1 vssd1 vccd1 vccd1 _15599_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2715 _07876_/X vssd1 vssd1 vccd1 vccd1 _15583_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07933_ hold1664/X _07924_/B _07932_/X _12199_/C1 vssd1 vssd1 vccd1 vccd1 _07933_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2726 _14075_/X vssd1 vssd1 vccd1 vccd1 _17842_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2737 _18090_/Q vssd1 vssd1 vccd1 vccd1 hold2737/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2748 _09201_/X vssd1 vssd1 vccd1 vccd1 _16212_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2759 _08194_/X vssd1 vssd1 vccd1 vccd1 _15733_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07864_ hold3043/X _07865_/B _07863_/Y _12265_/C1 vssd1 vssd1 vccd1 vccd1 _07864_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09603_ _09987_/A _09603_/B vssd1 vssd1 vccd1 vccd1 _09603_/X sky130_fd_sc_hd__or2_1
X_07795_ _18461_/Q hold1119/X _09342_/A _09438_/B vssd1 vssd1 vccd1 vccd1 _07795_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_09534_ _11061_/A _09534_/B vssd1 vssd1 vccd1 vccd1 _09534_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09465_ _09465_/A _09465_/B vssd1 vssd1 vccd1 vccd1 _16315_/D sky130_fd_sc_hd__nor2_1
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08416_ hold2591/X _08442_/A2 _08415_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08416_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09396_ _09386_/B _09369_/B _07809_/B vssd1 vssd1 vccd1 vccd1 _09396_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_173_wb_clk_i clkbuf_6_48_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18315_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08347_ _08347_/A _08347_/B vssd1 vssd1 vccd1 vccd1 _15805_/D sky130_fd_sc_hd__and2_1
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_102_wb_clk_i clkbuf_6_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18417_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08278_ _15557_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08278_/X sky130_fd_sc_hd__or2_1
Xhold6020 _17547_/Q vssd1 vssd1 vccd1 vccd1 hold6020/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6031 _17530_/Q vssd1 vssd1 vccd1 vccd1 hold6031/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6042 data_in[24] vssd1 vssd1 vccd1 vccd1 hold140/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6053 _18193_/Q vssd1 vssd1 vccd1 vccd1 hold6053/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6064 _18362_/Q vssd1 vssd1 vccd1 vccd1 hold6064/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5330 _11638_/X vssd1 vssd1 vccd1 vccd1 _17036_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6075 _18273_/Q vssd1 vssd1 vccd1 vccd1 hold6075/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6086 data_in[22] vssd1 vssd1 vccd1 vccd1 hold427/A sky130_fd_sc_hd__dlygate4sd3_1
X_10240_ hold3954/X _10649_/B _10239_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10240_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5341 _17610_/Q vssd1 vssd1 vccd1 vccd1 hold5341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6097 data_in[5] vssd1 vssd1 vccd1 vccd1 hold392/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5352 _13486_/X vssd1 vssd1 vccd1 vccd1 _17615_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5363 _11470_/X vssd1 vssd1 vccd1 vccd1 _16980_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5374 _17033_/Q vssd1 vssd1 vccd1 vccd1 hold5374/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4640 _16453_/Q vssd1 vssd1 vccd1 vccd1 hold4640/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5385 _12241_/X vssd1 vssd1 vccd1 vccd1 _17237_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10171_ hold3972/X _10649_/B _10170_/X _14691_/C1 vssd1 vssd1 vccd1 vccd1 _10171_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4651 _09808_/X vssd1 vssd1 vccd1 vccd1 _16426_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5396 _17711_/Q vssd1 vssd1 vccd1 vccd1 hold5396/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4662 _16482_/Q vssd1 vssd1 vccd1 vccd1 hold4662/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4673 _13348_/X vssd1 vssd1 vccd1 vccd1 _17569_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4684 _13537_/X vssd1 vssd1 vccd1 vccd1 _17632_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3950 _16480_/Q vssd1 vssd1 vccd1 vccd1 hold3950/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4695 _17180_/Q vssd1 vssd1 vccd1 vccd1 hold4695/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3961 _10711_/X vssd1 vssd1 vccd1 vccd1 _16727_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3972 _16579_/Q vssd1 vssd1 vccd1 vccd1 hold3972/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout151 _12851_/S vssd1 vssd1 vccd1 vccd1 _12848_/S sky130_fd_sc_hd__buf_6
Xhold3983 _09688_/X vssd1 vssd1 vccd1 vccd1 _16386_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout162 _13817_/B vssd1 vssd1 vccd1 vccd1 _13811_/B sky130_fd_sc_hd__buf_4
Xhold3994 _09763_/X vssd1 vssd1 vccd1 vccd1 _16411_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13930_ hold220/X _17773_/Q _13942_/S vssd1 vssd1 vccd1 vccd1 hold309/A sky130_fd_sc_hd__mux2_1
Xfanout173 _11717_/B vssd1 vssd1 vccd1 vccd1 _12305_/B sky130_fd_sc_hd__buf_4
XFILLER_0_96_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout184 _13868_/B vssd1 vssd1 vccd1 vccd1 _13856_/B sky130_fd_sc_hd__buf_4
Xfanout195 _12365_/B vssd1 vssd1 vccd1 vccd1 _12374_/B sky130_fd_sc_hd__buf_4
XFILLER_0_198_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13861_ _13888_/A _13861_/B vssd1 vssd1 vccd1 vccd1 _13861_/Y sky130_fd_sc_hd__nor2_1
X_15600_ _17280_/CLK _15600_/D vssd1 vssd1 vccd1 vccd1 _15600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12812_ hold3373/X _12811_/X _12812_/S vssd1 vssd1 vccd1 vccd1 _12812_/X sky130_fd_sc_hd__mux2_1
X_16580_ _18170_/CLK _16580_/D vssd1 vssd1 vccd1 vccd1 _16580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13792_ hold5603/X _13877_/B _13791_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13792_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_232_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15531_ _15531_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15531_/X sky130_fd_sc_hd__or2_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ hold3173/X _12742_/X _12749_/S vssd1 vssd1 vccd1 vccd1 _12743_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18250_ _18250_/CLK _18250_/D vssd1 vssd1 vccd1 vccd1 _18250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15462_ _15480_/A _15462_/B _15462_/C _15462_/D vssd1 vssd1 vccd1 vccd1 _15462_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12674_ hold3125/X _12673_/X _12851_/S vssd1 vssd1 vccd1 vccd1 _12674_/X sky130_fd_sc_hd__mux2_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _17266_/CLK _17201_/D vssd1 vssd1 vccd1 vccd1 _17201_/Q sky130_fd_sc_hd__dfxtp_1
X_14413_ _14413_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14413_/X sky130_fd_sc_hd__or2_1
XFILLER_0_38_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18181_ _18181_/CLK _18181_/D vssd1 vssd1 vccd1 vccd1 _18181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11625_ _12210_/A _11625_/B vssd1 vssd1 vccd1 vccd1 _11625_/X sky130_fd_sc_hd__or2_1
X_15393_ _15490_/A1 _15385_/X _15392_/X _15481_/B1 hold5914/A vssd1 vssd1 vccd1 vccd1
+ _15393_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_5_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17132_ _17260_/CLK _17132_/D vssd1 vssd1 vccd1 vccd1 _17132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14344_ _14344_/A _14344_/B vssd1 vssd1 vccd1 vccd1 _17971_/D sky130_fd_sc_hd__and2_1
XFILLER_0_163_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11556_ _11556_/A _11556_/B vssd1 vssd1 vccd1 vccd1 _11556_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10507_ _10601_/A _10601_/B _10506_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _16659_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17063_ _18448_/CLK _17063_/D vssd1 vssd1 vccd1 vccd1 _17063_/Q sky130_fd_sc_hd__dfxtp_1
X_14275_ hold1915/X _14272_/B _14274_/X _14342_/A vssd1 vssd1 vccd1 vccd1 _14275_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11487_ _11667_/A _11487_/B vssd1 vssd1 vccd1 vccd1 _11487_/X sky130_fd_sc_hd__or2_1
X_16014_ _18421_/CLK _16014_/D vssd1 vssd1 vccd1 vccd1 hold463/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13226_ _17579_/Q _17113_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13226_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10438_ hold5511/X _11213_/B _10437_/X _14342_/A vssd1 vssd1 vccd1 vccd1 _10438_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13157_ _13156_/X hold3468/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13157_/X sky130_fd_sc_hd__mux2_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10369_ hold3690/X _10601_/B _10368_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10369_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12108_ _12210_/A _12108_/B vssd1 vssd1 vccd1 vccd1 _12108_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _13081_/X _13087_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17529_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_209_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17965_ _17973_/CLK _17965_/D vssd1 vssd1 vccd1 vccd1 _17965_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12039_ _12267_/A _12039_/B vssd1 vssd1 vccd1 vccd1 _12039_/X sky130_fd_sc_hd__or2_1
X_16916_ _17894_/CLK _16916_/D vssd1 vssd1 vccd1 vccd1 _16916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17896_ _17936_/CLK _17896_/D vssd1 vssd1 vccd1 vccd1 _17896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16847_ _18050_/CLK _16847_/D vssd1 vssd1 vccd1 vccd1 _16847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16778_ _17981_/CLK _16778_/D vssd1 vssd1 vccd1 vccd1 _16778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15729_ _17732_/CLK _15729_/D vssd1 vssd1 vccd1 vccd1 _15729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_wb_clk_i clkbuf_6_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17456_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09250_ _12810_/A _09250_/B vssd1 vssd1 vccd1 vccd1 _16236_/D sky130_fd_sc_hd__and2_1
XFILLER_0_186_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18448_ _18448_/CLK _18448_/D vssd1 vssd1 vccd1 vccd1 _18448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08201_ _14529_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08201_/X sky130_fd_sc_hd__or2_1
XFILLER_0_111_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09181_ hold6050/X _09218_/B _09180_/X _12777_/A vssd1 vssd1 vccd1 vccd1 _09181_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18379_ _18379_/CLK _18379_/D vssd1 vssd1 vccd1 vccd1 _18379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08132_ _15537_/A hold1129/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08133_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08063_ hold2811/X _08097_/A2 _08062_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _08063_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3202 _16355_/Q vssd1 vssd1 vccd1 vccd1 _13310_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3213 _12965_/X vssd1 vssd1 vccd1 vccd1 _12966_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3224 _16375_/Q vssd1 vssd1 vccd1 vccd1 hold3224/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3235 _17368_/Q vssd1 vssd1 vccd1 vccd1 hold3235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3246 _09565_/X vssd1 vssd1 vccd1 vccd1 _16345_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2501 _18040_/Q vssd1 vssd1 vccd1 vccd1 hold2501/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08965_ hold180/X hold347/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold348/A sky130_fd_sc_hd__mux2_1
Xhold3257 _16656_/Q vssd1 vssd1 vccd1 vccd1 hold3257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2512 _15606_/Q vssd1 vssd1 vccd1 vccd1 hold2512/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2523 _14799_/X vssd1 vssd1 vccd1 vccd1 _18189_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3268 _17380_/Q vssd1 vssd1 vccd1 vccd1 hold3268/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2534 _18340_/Q vssd1 vssd1 vccd1 vccd1 hold2534/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3279 _09973_/X vssd1 vssd1 vccd1 vccd1 _16481_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2545 _14773_/X vssd1 vssd1 vccd1 vccd1 _18177_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1800 _14480_/X vssd1 vssd1 vccd1 vccd1 _18037_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1811 _17512_/Q vssd1 vssd1 vccd1 vccd1 hold1811/X sky130_fd_sc_hd__dlygate4sd3_1
X_07916_ _14604_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07916_/X sky130_fd_sc_hd__or2_1
Xhold2556 _14095_/X vssd1 vssd1 vccd1 vccd1 _17852_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1822 _15206_/X vssd1 vssd1 vccd1 vccd1 _18385_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08896_ hold169/X hold561/X _08930_/S vssd1 vssd1 vccd1 vccd1 hold562/A sky130_fd_sc_hd__mux2_1
Xhold2567 _15597_/Q vssd1 vssd1 vccd1 vccd1 hold2567/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1833 _18348_/Q vssd1 vssd1 vccd1 vccd1 hold1833/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2578 _14065_/X vssd1 vssd1 vccd1 vccd1 _17837_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1844 _14424_/X vssd1 vssd1 vccd1 vccd1 _18010_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2589 _15772_/Q vssd1 vssd1 vccd1 vccd1 hold2589/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1855 _18050_/Q vssd1 vssd1 vccd1 vccd1 hold1855/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1866 _07862_/X vssd1 vssd1 vccd1 vccd1 _15576_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07847_ _15525_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07847_/X sky130_fd_sc_hd__or2_1
XFILLER_0_230_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1877 _15725_/Q vssd1 vssd1 vccd1 vccd1 hold1877/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1888 _07832_/X vssd1 vssd1 vccd1 vccd1 _15561_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1899 _18186_/Q vssd1 vssd1 vccd1 vccd1 hold1899/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09517_ hold3750/X _10004_/B _09516_/X _15042_/A vssd1 vssd1 vccd1 vccd1 _09517_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_354_wb_clk_i clkbuf_6_40_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17740_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _09447_/A _09444_/X _09478_/B vssd1 vssd1 vccd1 vccd1 _09449_/B sky130_fd_sc_hd__o21ai_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09379_ _17326_/Q _15487_/A2 _09392_/C hold431/X _09378_/X vssd1 vssd1 vccd1 vccd1
+ _09383_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_192_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11410_ hold5426/X _11792_/B _11409_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _11410_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12390_ _12390_/A _12390_/B vssd1 vssd1 vccd1 vccd1 _17288_/D sky130_fd_sc_hd__and2_1
XFILLER_0_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11341_ hold5359/X _11726_/B _11340_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _11341_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14060_ _15513_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14060_/X sky130_fd_sc_hd__or2_1
X_11272_ hold5103/X _11753_/B _11271_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _11272_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5160 _10789_/X vssd1 vssd1 vccd1 vccd1 _16753_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13011_ _15515_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13011_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10223_ hold2991/X hold3811/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10224_/B sky130_fd_sc_hd__mux2_1
Xhold5171 _17281_/Q vssd1 vssd1 vccd1 vccd1 hold5171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5182 _10705_/X vssd1 vssd1 vccd1 vccd1 _16725_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5193 _17744_/Q vssd1 vssd1 vccd1 vccd1 hold5193/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_70_wb_clk_i clkbuf_6_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17500_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4470 _11151_/Y vssd1 vssd1 vccd1 vccd1 _11152_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10154_ hold2380/X hold3441/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10155_/B sky130_fd_sc_hd__mux2_1
Xhold4481 _12073_/X vssd1 vssd1 vccd1 vccd1 _17181_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4492 _11848_/X vssd1 vssd1 vccd1 vccd1 _17106_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3780 _10141_/X vssd1 vssd1 vccd1 vccd1 _16537_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14962_ hold289/X hold407/X vssd1 vssd1 vccd1 vccd1 hold408/A sky130_fd_sc_hd__or2_1
X_17750_ _17750_/CLK _17750_/D vssd1 vssd1 vccd1 vccd1 _17750_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3791 _16872_/Q vssd1 vssd1 vccd1 vccd1 hold3791/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ hold2279/X hold3417/X _10571_/C vssd1 vssd1 vccd1 vccd1 _10086_/B sky130_fd_sc_hd__mux2_1
XTAP_5964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16701_ _18227_/CLK _16701_/D vssd1 vssd1 vccd1 vccd1 _16701_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13913_ _13923_/A _13913_/B vssd1 vssd1 vccd1 vccd1 _17764_/D sky130_fd_sc_hd__and2_1
X_14893_ hold1829/X _14880_/B _14892_/X _14893_/C1 vssd1 vssd1 vccd1 vccd1 _14893_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17681_ _17745_/CLK _17681_/D vssd1 vssd1 vccd1 vccd1 _17681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16632_ _18194_/CLK _16632_/D vssd1 vssd1 vccd1 vccd1 _16632_/Q sky130_fd_sc_hd__dfxtp_1
X_13844_ _17735_/Q _13886_/B _13886_/C vssd1 vssd1 vccd1 vccd1 _13844_/X sky130_fd_sc_hd__and3_1
XFILLER_0_226_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16563_ _18177_/CLK _16563_/D vssd1 vssd1 vccd1 vccd1 _16563_/Q sky130_fd_sc_hd__dfxtp_1
X_13775_ hold2304/X _17712_/Q _13871_/C vssd1 vssd1 vccd1 vccd1 _13776_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10987_ hold3808/X _11204_/B _10986_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _10987_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18302_ _18423_/CLK _18302_/D vssd1 vssd1 vccd1 vccd1 _18302_/Q sky130_fd_sc_hd__dfxtp_1
X_12726_ _12753_/A _12726_/B vssd1 vssd1 vccd1 vccd1 _17418_/D sky130_fd_sc_hd__and2_1
X_15514_ hold2863/X _15560_/A2 _15513_/X _12864_/A vssd1 vssd1 vccd1 vccd1 _15514_/X
+ sky130_fd_sc_hd__o211a_1
X_16494_ _18375_/CLK _16494_/D vssd1 vssd1 vccd1 vccd1 _16494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15445_ hold463/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15445_/X sky130_fd_sc_hd__or2_1
X_18233_ _18233_/CLK _18233_/D vssd1 vssd1 vccd1 vccd1 _18233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12657_ _12873_/A _12657_/B vssd1 vssd1 vccd1 vccd1 _17395_/D sky130_fd_sc_hd__and2_1
XFILLER_0_210_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11608_ hold3866/X _11798_/B _11607_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _11608_/X
+ sky130_fd_sc_hd__o211a_1
X_15376_ _17341_/Q _15486_/B1 _09362_/D _16118_/Q vssd1 vssd1 vccd1 vccd1 _15376_/X
+ sky130_fd_sc_hd__a22o_1
X_18164_ _18164_/CLK _18164_/D vssd1 vssd1 vccd1 vccd1 _18164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12588_ _12588_/A _12588_/B vssd1 vssd1 vccd1 vccd1 _17372_/D sky130_fd_sc_hd__and2_1
XFILLER_0_111_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14327_ hold2507/X _14326_/B _14326_/Y _14342_/A vssd1 vssd1 vccd1 vccd1 _14327_/X
+ sky130_fd_sc_hd__o211a_1
X_17115_ _17741_/CLK _17115_/D vssd1 vssd1 vccd1 vccd1 _17115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18095_ _18223_/CLK _18095_/D vssd1 vssd1 vccd1 vccd1 _18095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11539_ hold5002/X _11726_/B _11538_/X _13895_/A vssd1 vssd1 vccd1 vccd1 _11539_/X
+ sky130_fd_sc_hd__o211a_1
Xhold407 hold407/A vssd1 vssd1 vccd1 vccd1 hold407/X sky130_fd_sc_hd__buf_4
Xhold418 hold418/A vssd1 vssd1 vccd1 vccd1 hold418/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17046_ _17894_/CLK _17046_/D vssd1 vssd1 vccd1 vccd1 _17046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold429 input19/X vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__buf_1
X_14258_ _15099_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14258_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13209_ _13209_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13209_/X sky130_fd_sc_hd__and2_1
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ hold2053/X _14202_/B _14188_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _14189_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout909 hold289/X vssd1 vssd1 vccd1 vccd1 _15231_/A sky130_fd_sc_hd__buf_12
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08750_ _15414_/A hold780/X vssd1 vssd1 vccd1 vccd1 _15995_/D sky130_fd_sc_hd__and2_1
Xhold1107 hold1107/A vssd1 vssd1 vccd1 vccd1 _15203_/A sky130_fd_sc_hd__buf_12
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _18014_/CLK _17948_/D vssd1 vssd1 vccd1 vccd1 _17948_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1118 _14227_/X vssd1 vssd1 vccd1 vccd1 _17915_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1129 _15705_/Q vssd1 vssd1 vccd1 vccd1 hold1129/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_240_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08681_ hold452/X hold865/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08682_/B sky130_fd_sc_hd__mux2_1
X_17879_ _18448_/CLK _17879_/D vssd1 vssd1 vccd1 vccd1 _17879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_232_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_215_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09302_ hold1149/X _09325_/B _09301_/X _12906_/A vssd1 vssd1 vccd1 vccd1 _09302_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09233_ _14164_/A hold1654/X hold271/X vssd1 vssd1 vccd1 vccd1 _09233_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09164_ _15547_/A _09164_/B vssd1 vssd1 vccd1 vccd1 _09164_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_161_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08115_ _08115_/A _08115_/B vssd1 vssd1 vccd1 vccd1 _15696_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09095_ hold2002/X _09102_/B _09094_/X _12978_/A vssd1 vssd1 vccd1 vccd1 _09095_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08046_ hold969/X _08033_/B _08045_/X _08151_/A vssd1 vssd1 vccd1 vccd1 hold970/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold930 hold930/A vssd1 vssd1 vccd1 vccd1 input66/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_222_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold941 hold941/A vssd1 vssd1 vccd1 vccd1 hold941/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold952 hold952/A vssd1 vssd1 vccd1 vccd1 hold952/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 hold963/A vssd1 vssd1 vccd1 vccd1 hold963/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold974 la_data_in[4] vssd1 vssd1 vccd1 vccd1 hold974/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3010 _16186_/Q vssd1 vssd1 vccd1 vccd1 hold3010/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold985 hold985/A vssd1 vssd1 vccd1 vccd1 hold985/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 hold996/A vssd1 vssd1 vccd1 vccd1 hold996/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3021 _16192_/Q vssd1 vssd1 vccd1 vccd1 hold3021/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3032 _14428_/X vssd1 vssd1 vccd1 vccd1 _18012_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3043 _15577_/Q vssd1 vssd1 vccd1 vccd1 hold3043/X sky130_fd_sc_hd__dlygate4sd3_1
X_09997_ _11203_/A _09997_/B vssd1 vssd1 vccd1 vccd1 _09997_/Y sky130_fd_sc_hd__nor2_1
XTAP_5216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3054 _07973_/X vssd1 vssd1 vccd1 vccd1 _15629_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3065 _18253_/Q vssd1 vssd1 vccd1 vccd1 hold3065/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2320 _15882_/Q vssd1 vssd1 vccd1 vccd1 hold2320/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2331 _18437_/Q vssd1 vssd1 vccd1 vccd1 hold2331/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3076 _15836_/Q vssd1 vssd1 vccd1 vccd1 hold3076/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08948_ _15274_/A _08948_/B vssd1 vssd1 vccd1 vccd1 _16091_/D sky130_fd_sc_hd__and2_1
Xhold3087 _18383_/Q vssd1 vssd1 vccd1 vccd1 hold3087/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2342 _08294_/X vssd1 vssd1 vccd1 vccd1 _15780_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3098 _14645_/X vssd1 vssd1 vccd1 vccd1 _18115_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2353 _18067_/Q vssd1 vssd1 vccd1 vccd1 hold2353/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2364 _13987_/X vssd1 vssd1 vccd1 vccd1 _17800_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2375 _15721_/Q vssd1 vssd1 vccd1 vccd1 hold2375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1630 _15585_/Q vssd1 vssd1 vccd1 vccd1 hold1630/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1641 _16196_/Q vssd1 vssd1 vccd1 vccd1 hold1641/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2386 _15872_/Q vssd1 vssd1 vccd1 vccd1 hold2386/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1652 _18108_/Q vssd1 vssd1 vccd1 vccd1 hold1652/X sky130_fd_sc_hd__dlygate4sd3_1
X_08879_ _12390_/A _08879_/B vssd1 vssd1 vccd1 vccd1 _16057_/D sky130_fd_sc_hd__and2_1
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2397 _08020_/X vssd1 vssd1 vccd1 vccd1 _15651_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1663 _14329_/X vssd1 vssd1 vccd1 vccd1 _17964_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1674 _17953_/Q vssd1 vssd1 vccd1 vccd1 hold1674/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10910_ hold2083/X hold5549/X _11213_/C vssd1 vssd1 vccd1 vccd1 _10911_/B sky130_fd_sc_hd__mux2_1
Xhold1685 _14530_/X vssd1 vssd1 vccd1 vccd1 _18061_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_230_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1696 _16275_/Q vssd1 vssd1 vccd1 vccd1 hold1696/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ hold5251/X _13886_/B _11889_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _11890_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10841_ hold2292/X _16771_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _10842_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13560_ _13752_/A _13560_/B vssd1 vssd1 vccd1 vccd1 _13560_/X sky130_fd_sc_hd__or2_1
X_10772_ hold1588/X _16748_/Q _10964_/S vssd1 vssd1 vccd1 vccd1 _10773_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_136_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12511_ _07809_/X _12510_/Y _13048_/A hold2264/X vssd1 vssd1 vccd1 vccd1 _12511_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_176_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13491_ _13788_/A _13491_/B vssd1 vssd1 vccd1 vccd1 _13491_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15230_ hold2933/X _15221_/B _15229_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _15230_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12442_ _15314_/A _12442_/B vssd1 vssd1 vccd1 vccd1 _17314_/D sky130_fd_sc_hd__and2_1
XFILLER_0_136_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15161_ _15161_/A _15165_/B vssd1 vssd1 vccd1 vccd1 _15161_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_140_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12373_ _13888_/A _12373_/B vssd1 vssd1 vccd1 vccd1 _12373_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_105_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14112_ hold915/X _14160_/B vssd1 vssd1 vccd1 vccd1 _14112_/X sky130_fd_sc_hd__or2_1
XFILLER_0_205_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11324_ hold1238/X hold4111/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11325_/B sky130_fd_sc_hd__mux2_1
X_15092_ hold2257/X hold341/X _15091_/X _15228_/C1 vssd1 vssd1 vccd1 vccd1 _15092_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14043_ hold1409/X _14040_/B _14042_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _14043_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11255_ hold2903/X hold4636/X _11738_/C vssd1 vssd1 vccd1 vccd1 _11256_/B sky130_fd_sc_hd__mux2_1
X_10206_ _10470_/A _10206_/B vssd1 vssd1 vccd1 vccd1 _10206_/X sky130_fd_sc_hd__or2_1
XTAP_6440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11186_ _16886_/Q _11186_/B _11186_/C vssd1 vssd1 vccd1 vccd1 _11186_/X sky130_fd_sc_hd__and3_1
XTAP_6451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17802_ _17894_/CLK _17802_/D vssd1 vssd1 vccd1 vccd1 _17802_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10137_ _11121_/A _10137_/B vssd1 vssd1 vccd1 vccd1 _10137_/X sky130_fd_sc_hd__or2_1
XTAP_6484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15994_ _16058_/CLK _15994_/D vssd1 vssd1 vccd1 vccd1 hold873/A sky130_fd_sc_hd__dfxtp_1
XTAP_5761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_276_wb_clk_i clkbuf_6_51_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18391_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17733_ _17733_/CLK _17733_/D vssd1 vssd1 vccd1 vccd1 _17733_/Q sky130_fd_sc_hd__dfxtp_1
X_10068_ _13294_/A _09978_/A _10067_/X vssd1 vssd1 vccd1 vccd1 _10069_/B sky130_fd_sc_hd__a21oi_1
X_14945_ hold2143/X _14952_/B _14944_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _14945_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_238_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_205_wb_clk_i clkbuf_6_55_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18296_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17664_ _17728_/CLK _17664_/D vssd1 vssd1 vccd1 vccd1 _17664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14876_ _15161_/A _14880_/B vssd1 vssd1 vccd1 vccd1 _14876_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16615_ _18203_/CLK _16615_/D vssd1 vssd1 vccd1 vccd1 _16615_/Q sky130_fd_sc_hd__dfxtp_1
X_13827_ hold4230/X _13737_/A _13826_/X vssd1 vssd1 vccd1 vccd1 _13827_/Y sky130_fd_sc_hd__a21oi_1
X_17595_ _17689_/CLK _17595_/D vssd1 vssd1 vccd1 vccd1 _17595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16546_ _18168_/CLK _16546_/D vssd1 vssd1 vccd1 vccd1 _16546_/Q sky130_fd_sc_hd__dfxtp_1
X_13758_ _13758_/A _13758_/B vssd1 vssd1 vccd1 vccd1 _13758_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12709_ hold2337/X hold3826/X _12766_/S vssd1 vssd1 vccd1 vccd1 _12709_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16477_ _18390_/CLK _16477_/D vssd1 vssd1 vccd1 vccd1 _16477_/Q sky130_fd_sc_hd__dfxtp_1
X_13689_ _13788_/A _13689_/B vssd1 vssd1 vccd1 vccd1 _13689_/X sky130_fd_sc_hd__or2_1
XFILLER_0_72_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18216_ _18222_/CLK _18216_/D vssd1 vssd1 vccd1 vccd1 _18216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15428_ hold207/X _09367_/A _09362_/C _17346_/Q vssd1 vssd1 vccd1 vccd1 _15428_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18147_ _18215_/CLK _18147_/D vssd1 vssd1 vccd1 vccd1 _18147_/Q sky130_fd_sc_hd__dfxtp_1
X_15359_ hold533/X _15485_/A2 _09392_/C hold601/X _15358_/X vssd1 vssd1 vccd1 vccd1
+ _15362_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5907 _18400_/Q vssd1 vssd1 vccd1 vccd1 hold5907/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5918 hold5918/A vssd1 vssd1 vccd1 vccd1 hold5918/X sky130_fd_sc_hd__buf_2
XFILLER_0_223_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold204 hold204/A vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5929 hold5929/A vssd1 vssd1 vccd1 vccd1 hold5929/X sky130_fd_sc_hd__buf_2
XFILLER_0_111_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold215 hold32/X vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__buf_4
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold226 hold26/X vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__buf_4
X_18078_ _18393_/CLK _18078_/D vssd1 vssd1 vccd1 vccd1 _18078_/Q sky130_fd_sc_hd__dfxtp_1
Xhold237 hold237/A vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold248 hold76/X vssd1 vssd1 vccd1 vccd1 input8/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09920_ hold3186/X hold5080/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09921_/B sky130_fd_sc_hd__mux2_1
Xhold259 input31/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17029_ _17877_/CLK _17029_/D vssd1 vssd1 vccd1 vccd1 _17029_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout706 _09047_/A vssd1 vssd1 vccd1 vccd1 _09057_/A sky130_fd_sc_hd__buf_2
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09851_ hold1903/X _16441_/Q _10031_/C vssd1 vssd1 vccd1 vccd1 _09852_/B sky130_fd_sc_hd__mux2_1
Xfanout717 _09907_/C1 vssd1 vssd1 vccd1 vccd1 _14368_/A sky130_fd_sc_hd__clkbuf_4
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout728 _09907_/C1 vssd1 vssd1 vccd1 vccd1 _12418_/A sky130_fd_sc_hd__clkbuf_4
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 _07787_/Y vssd1 vssd1 vccd1 vccd1 fanout739/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_237_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _12440_/A hold432/X vssd1 vssd1 vccd1 vccd1 _16020_/D sky130_fd_sc_hd__and2_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ hold3008/X hold3982/X _11204_/C vssd1 vssd1 vccd1 vccd1 _09783_/B sky130_fd_sc_hd__mux2_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ hold618/X hold854/X _08779_/S vssd1 vssd1 vccd1 vccd1 hold855/A sky130_fd_sc_hd__mux2_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08664_ _08730_/A _12380_/B vssd1 vssd1 vccd1 vccd1 _08723_/S sky130_fd_sc_hd__or2_2
XFILLER_0_212_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08595_ _15324_/A hold491/X vssd1 vssd1 vccd1 vccd1 _15921_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09216_ _15545_/A _09218_/B vssd1 vssd1 vccd1 vccd1 _09216_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09147_ hold3010/X _09164_/B _09146_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _09147_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09078_ _15519_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09078_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08029_ _15543_/A _08029_/B vssd1 vssd1 vccd1 vccd1 _08029_/Y sky130_fd_sc_hd__nand2_1
Xhold760 hold760/A vssd1 vssd1 vccd1 vccd1 hold760/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold771 hold771/A vssd1 vssd1 vccd1 vccd1 hold771/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold782 hold782/A vssd1 vssd1 vccd1 vccd1 hold782/X sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ _11136_/A _11040_/B vssd1 vssd1 vccd1 vccd1 _11040_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold793 hold793/A vssd1 vssd1 vccd1 vccd1 hold793/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2150 _14223_/X vssd1 vssd1 vccd1 vccd1 _17913_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2161 _18180_/Q vssd1 vssd1 vccd1 vccd1 hold2161/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2172 _14450_/X vssd1 vssd1 vccd1 vccd1 _18022_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12991_ hold2580/X hold4747/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12991_/X sky130_fd_sc_hd__mux2_1
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2183 _17945_/Q vssd1 vssd1 vccd1 vccd1 hold2183/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2194 _09153_/X vssd1 vssd1 vccd1 vccd1 _16189_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_232_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1460 _07937_/X vssd1 vssd1 vccd1 vccd1 _15612_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14730_ _15231_/A _14730_/B vssd1 vssd1 vccd1 vccd1 _14730_/X sky130_fd_sc_hd__or2_1
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1471 _15775_/Q vssd1 vssd1 vccd1 vccd1 hold1471/X sky130_fd_sc_hd__dlygate4sd3_1
X_11942_ hold1275/X hold4491/X _12362_/C vssd1 vssd1 vccd1 vccd1 _11943_/B sky130_fd_sc_hd__mux2_1
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1482 _14017_/X vssd1 vssd1 vccd1 vccd1 _17814_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1493 hold6131/X vssd1 vssd1 vccd1 vccd1 _09463_/B sky130_fd_sc_hd__buf_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ hold2991/X _14664_/B _14660_/Y _14877_/C1 vssd1 vssd1 vccd1 vccd1 _14661_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11873_ hold535/X hold4273/X _13481_/S vssd1 vssd1 vccd1 vccd1 _11874_/B sky130_fd_sc_hd__mux2_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16400_ _18345_/CLK _16400_/D vssd1 vssd1 vccd1 vccd1 _16400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13612_ hold5797/X _13808_/B _13611_/X _12738_/A vssd1 vssd1 vccd1 vccd1 _13612_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ _11661_/A _10824_/B vssd1 vssd1 vccd1 vccd1 _10824_/X sky130_fd_sc_hd__or2_1
XFILLER_0_200_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14592_ _15201_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14592_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17380_ _17380_/CLK _17380_/D vssd1 vssd1 vccd1 vccd1 _17380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16331_ _17535_/CLK _16331_/D vssd1 vssd1 vccd1 vccd1 _16331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13543_ hold4541/X _13829_/B _13542_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13543_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10755_ _11637_/A _10755_/B vssd1 vssd1 vccd1 vccd1 _10755_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16262_ _17374_/CLK _16262_/D vssd1 vssd1 vccd1 vccd1 _16262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13474_ hold5513/X _13847_/B _13473_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13474_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10686_ _11655_/A _10686_/B vssd1 vssd1 vccd1 vccd1 _10686_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15213_ _15213_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15213_/X sky130_fd_sc_hd__or2_1
X_18001_ _18053_/CLK _18001_/D vssd1 vssd1 vccd1 vccd1 _18001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12425_ hold53/X hold457/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12426_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16193_ _17476_/CLK _16193_/D vssd1 vssd1 vccd1 vccd1 _16193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15144_ hold984/X _15167_/B _15143_/X _15064_/A vssd1 vssd1 vccd1 vccd1 hold985/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12356_ _17276_/Q _12356_/B _13481_/S vssd1 vssd1 vccd1 vccd1 _12356_/X sky130_fd_sc_hd__and3_1
XFILLER_0_65_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11307_ _11667_/A _11307_/B vssd1 vssd1 vccd1 vccd1 _11307_/X sky130_fd_sc_hd__or2_1
X_15075_ _15183_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15075_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12287_ hold1630/X _17253_/Q _13409_/S vssd1 vssd1 vccd1 vccd1 _12288_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14026_ _15533_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14026_/X sky130_fd_sc_hd__or2_1
XFILLER_0_205_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_457_wb_clk_i clkbuf_6_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17445_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11238_ _11622_/A _11238_/B vssd1 vssd1 vccd1 vccd1 _11238_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11169_ hold3523/X _11649_/A _11168_/X vssd1 vssd1 vccd1 vccd1 _11169_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15977_ _18425_/CLK _15977_/D vssd1 vssd1 vccd1 vccd1 hold533/A sky130_fd_sc_hd__dfxtp_1
XTAP_5580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17716_ _17716_/CLK _17716_/D vssd1 vssd1 vccd1 vccd1 _17716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14928_ _15197_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14928_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17647_ _17672_/CLK _17647_/D vssd1 vssd1 vccd1 vccd1 _17647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14859_ hold1089/X hold332/X _14858_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14859_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_230_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08380_ _14543_/A hold1066/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08381_/B sky130_fd_sc_hd__mux2_1
X_17578_ _17738_/CLK _17578_/D vssd1 vssd1 vccd1 vccd1 _17578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16529_ _18149_/CLK _16529_/D vssd1 vssd1 vccd1 vccd1 _16529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09001_ _09057_/A hold265/X vssd1 vssd1 vccd1 vccd1 _16117_/D sky130_fd_sc_hd__and2_1
XFILLER_0_147_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_1293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5704 _11527_/X vssd1 vssd1 vccd1 vccd1 _16999_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5715 _12351_/Y vssd1 vssd1 vccd1 vccd1 _12352_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5726 _17565_/Q vssd1 vssd1 vccd1 vccd1 hold5726/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5737 _17277_/Q vssd1 vssd1 vccd1 vccd1 hold5737/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5748 _10011_/Y vssd1 vssd1 vccd1 vccd1 _10012_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5759 _17273_/Q vssd1 vssd1 vccd1 vccd1 hold5759/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_198_wb_clk_i clkbuf_6_53_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18380_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09903_ _11067_/A _09903_/B vssd1 vssd1 vccd1 vccd1 _09903_/X sky130_fd_sc_hd__or2_1
Xfanout503 _11183_/C vssd1 vssd1 vccd1 vccd1 _11213_/C sky130_fd_sc_hd__buf_6
Xfanout514 _10385_/S vssd1 vssd1 vccd1 vccd1 _10601_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_201_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout525 _09285_/Y vssd1 vssd1 vccd1 vccd1 _09325_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout536 _09102_/B vssd1 vssd1 vccd1 vccd1 _09106_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09834_ _09948_/A _09834_/B vssd1 vssd1 vccd1 vccd1 _09834_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_127_wb_clk_i clkbuf_6_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18410_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout547 _08393_/Y vssd1 vssd1 vccd1 vccd1 _08433_/B sky130_fd_sc_hd__clkbuf_8
Xfanout558 _08173_/Y vssd1 vssd1 vccd1 vccd1 _08213_/B sky130_fd_sc_hd__buf_8
Xfanout569 _07938_/Y vssd1 vssd1 vccd1 vccd1 _07991_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_77_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09765_ _09957_/A _09765_/B vssd1 vssd1 vccd1 vccd1 _09765_/X sky130_fd_sc_hd__or2_1
XFILLER_0_225_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_214_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08716_ _12418_/A _08716_/B vssd1 vssd1 vccd1 vccd1 _15979_/D sky130_fd_sc_hd__and2_1
XFILLER_0_55_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09696_ _09912_/A _09696_/B vssd1 vssd1 vccd1 vccd1 _09696_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08647_ hold143/X hold592/X _08657_/S vssd1 vssd1 vccd1 vccd1 _08648_/B sky130_fd_sc_hd__mux2_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08578_ hold92/X hold620/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold621/A sky130_fd_sc_hd__mux2_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10540_ _10634_/A _10598_/B _10539_/X _10564_/C1 vssd1 vssd1 vccd1 vccd1 _10540_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10471_ _10565_/A _10568_/B _10470_/X _14893_/C1 vssd1 vssd1 vccd1 vccd1 _10471_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12210_ _12210_/A _12210_/B vssd1 vssd1 vccd1 vccd1 _12210_/X sky130_fd_sc_hd__or2_1
XFILLER_0_228_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13190_ _13190_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13190_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12141_ _12255_/A _12141_/B vssd1 vssd1 vccd1 vccd1 _12141_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12072_ _12267_/A _12072_/B vssd1 vssd1 vccd1 vccd1 _12072_/X sky130_fd_sc_hd__or2_1
Xhold590 hold590/A vssd1 vssd1 vccd1 vccd1 hold590/X sky130_fd_sc_hd__dlygate4sd3_1
X_15900_ _17303_/CLK _15900_/D vssd1 vssd1 vccd1 vccd1 hold411/A sky130_fd_sc_hd__dfxtp_1
X_11023_ hold3956/X _10616_/B _11022_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _11023_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16880_ _18039_/CLK _16880_/D vssd1 vssd1 vccd1 vccd1 _16880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15831_ _17626_/CLK _15831_/D vssd1 vssd1 vccd1 vccd1 _15831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ hold4137/X _12973_/X _12986_/S vssd1 vssd1 vccd1 vccd1 _12975_/B sky130_fd_sc_hd__mux2_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15762_ _17620_/CLK _15762_/D vssd1 vssd1 vccd1 vccd1 _15762_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ _17513_/CLK _17501_/D vssd1 vssd1 vccd1 vccd1 _17501_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1290 _13973_/X vssd1 vssd1 vccd1 vccd1 _17793_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14713_ hold2021/X _14720_/B _14712_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _14713_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_213_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11925_ _13800_/A _11925_/B vssd1 vssd1 vccd1 vccd1 _11925_/X sky130_fd_sc_hd__or2_1
XFILLER_0_234_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _17229_/CLK _15693_/D vssd1 vssd1 vccd1 vccd1 _15693_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17432_ _17440_/CLK _17432_/D vssd1 vssd1 vccd1 vccd1 _17432_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_47_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_47_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_14644_ _15199_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14644_/X sky130_fd_sc_hd__or2_1
X_11856_ _12240_/A _11856_/B vssd1 vssd1 vccd1 vccd1 _11856_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10807_ hold5303/X _11225_/B _10806_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10807_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14575_ hold1947/X _14610_/B _14574_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _14575_/X
+ sky130_fd_sc_hd__o211a_1
X_17363_ _17374_/CLK _17363_/D vssd1 vssd1 vccd1 vccd1 _17363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11787_ hold4449/X _11667_/A _11786_/X vssd1 vssd1 vccd1 vccd1 _11787_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16314_ _16315_/CLK _16314_/D vssd1 vssd1 vccd1 vccd1 _16314_/Q sky130_fd_sc_hd__dfxtp_1
X_10738_ hold5227/X _11225_/B _10737_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _10738_/X
+ sky130_fd_sc_hd__o211a_1
X_13526_ hold2478/X _17629_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13527_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_83_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17294_ _17337_/CLK _17294_/D vssd1 vssd1 vccd1 vccd1 hold357/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13457_ hold1791/X hold5502/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13458_/B sky130_fd_sc_hd__mux2_1
X_16245_ _17425_/CLK _16245_/D vssd1 vssd1 vccd1 vccd1 _16245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10669_ hold4899/X _11144_/B _10668_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _10669_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_1406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12408_ _12438_/A hold170/X vssd1 vssd1 vccd1 vccd1 _17297_/D sky130_fd_sc_hd__and2_1
XFILLER_0_24_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13388_ hold2386/X hold3493/X _13463_/S vssd1 vssd1 vccd1 vccd1 _13389_/B sky130_fd_sc_hd__mux2_1
X_16176_ _17468_/CLK _16176_/D vssd1 vssd1 vccd1 vccd1 _16176_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput106 hold5971/X vssd1 vssd1 vccd1 vccd1 ki sky130_fd_sc_hd__buf_12
XFILLER_0_112_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput117 hold5960/X vssd1 vssd1 vccd1 vccd1 hold5961/A sky130_fd_sc_hd__buf_6
X_15127_ _15128_/A _15182_/B vssd1 vssd1 vccd1 vccd1 _15127_/Y sky130_fd_sc_hd__nor2_2
Xoutput128 hold5947/X vssd1 vssd1 vccd1 vccd1 hold5948/A sky130_fd_sc_hd__buf_6
X_12339_ hold5711/X _12255_/A _12338_/X vssd1 vssd1 vccd1 vccd1 _12339_/Y sky130_fd_sc_hd__a21oi_1
Xoutput139 _09339_/A vssd1 vssd1 vccd1 vccd1 load_data sky130_fd_sc_hd__buf_12
XFILLER_0_107_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3609 _10285_/X vssd1 vssd1 vccd1 vccd1 _16585_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15058_ _15068_/A hold789/X vssd1 vssd1 vccd1 vccd1 _18314_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_291_wb_clk_i clkbuf_6_37_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17859_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2908 _17950_/Q vssd1 vssd1 vccd1 vccd1 hold2908/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2919 _14653_/X vssd1 vssd1 vccd1 vccd1 _18119_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14009_ hold2711/X _14040_/B _14008_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _14009_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_220_wb_clk_i clkbuf_6_61_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18217_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07880_ hold1630/X _07865_/B _07879_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _07880_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09550_ hold4512/X _10028_/B _09549_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09550_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08501_ hold1161/X _08488_/B _08500_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _08501_/X
+ sky130_fd_sc_hd__o211a_1
X_09481_ _09482_/B _09484_/B _09481_/C vssd1 vssd1 vccd1 vccd1 _16321_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_76_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08432_ hold1330/X _08433_/B _08431_/Y _08389_/A vssd1 vssd1 vccd1 vccd1 _08432_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_1333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08363_ _08363_/A _08363_/B vssd1 vssd1 vccd1 vccd1 _15813_/D sky130_fd_sc_hd__and2_1
XFILLER_0_191_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08294_ hold2341/X _08336_/A2 _08293_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _08294_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_379_wb_clk_i clkbuf_6_33_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17614_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5501 _11323_/X vssd1 vssd1 vccd1 vccd1 _16931_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5512 _10438_/X vssd1 vssd1 vccd1 vccd1 _16636_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5523 _16848_/Q vssd1 vssd1 vccd1 vccd1 hold5523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5534 _13468_/X vssd1 vssd1 vccd1 vccd1 _17609_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4800 _10657_/X vssd1 vssd1 vccd1 vccd1 _16709_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5545 _17748_/Q vssd1 vssd1 vccd1 vccd1 hold5545/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_308_wb_clk_i clkbuf_6_45_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17968_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_160_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5556 _13687_/X vssd1 vssd1 vccd1 vccd1 _17682_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4811 _17226_/Q vssd1 vssd1 vccd1 vccd1 hold4811/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4822 _10969_/X vssd1 vssd1 vccd1 vccd1 _16813_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5567 _17062_/Q vssd1 vssd1 vccd1 vccd1 hold5567/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4833 _16390_/Q vssd1 vssd1 vccd1 vccd1 hold4833/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5578 _11545_/X vssd1 vssd1 vccd1 vccd1 _17005_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4844 _12259_/X vssd1 vssd1 vccd1 vccd1 _17243_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5589 _17088_/Q vssd1 vssd1 vccd1 vccd1 hold5589/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4855 _17264_/Q vssd1 vssd1 vccd1 vccd1 hold4855/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout300 _11049_/A vssd1 vssd1 vccd1 vccd1 _11136_/A sky130_fd_sc_hd__buf_4
Xhold4866 _12079_/X vssd1 vssd1 vccd1 vccd1 _17183_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout311 wire337/X vssd1 vssd1 vccd1 vccd1 _11061_/A sky130_fd_sc_hd__clkbuf_8
Xhold4877 _16943_/Q vssd1 vssd1 vccd1 vccd1 hold4877/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4888 _11287_/X vssd1 vssd1 vccd1 vccd1 _16919_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout322 _10539_/A vssd1 vssd1 vccd1 vccd1 _10413_/A sky130_fd_sc_hd__buf_2
Xhold4899 _16745_/Q vssd1 vssd1 vccd1 vccd1 hold4899/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout333 _10542_/A vssd1 vssd1 vccd1 vccd1 _10524_/A sky130_fd_sc_hd__buf_4
XFILLER_0_61_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout344 _15489_/A vssd1 vssd1 vccd1 vccd1 _15480_/A sky130_fd_sc_hd__buf_4
Xfanout355 _08723_/S vssd1 vssd1 vccd1 vccd1 _08721_/S sky130_fd_sc_hd__buf_8
XFILLER_0_219_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout366 _15157_/B vssd1 vssd1 vccd1 vccd1 _15179_/B sky130_fd_sc_hd__buf_6
X_09817_ hold3574/X _10031_/B _09816_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09817_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout377 hold407/X vssd1 vssd1 vccd1 vccd1 _14964_/B sky130_fd_sc_hd__buf_6
XFILLER_0_226_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout388 _14734_/Y vssd1 vssd1 vccd1 vccd1 _14774_/B sky130_fd_sc_hd__buf_8
Xfanout399 _14447_/Y vssd1 vssd1 vccd1 vccd1 _14487_/B sky130_fd_sc_hd__buf_8
XFILLER_0_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09748_ hold4169/X _10052_/B _09747_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09748_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_213_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ hold3216/X _10601_/B _09678_/X _15204_/C1 vssd1 vssd1 vccd1 vccd1 _09679_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_95_wb_clk_i clkbuf_6_19_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17300_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_139_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ hold5225/X _12317_/B _11709_/X _14211_/C1 vssd1 vssd1 vccd1 vccd1 _11710_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12849_/A _12690_/B vssd1 vssd1 vccd1 vccd1 _17406_/D sky130_fd_sc_hd__and2_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_wb_clk_i clkbuf_6_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17380_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11641_ hold5583/X _11744_/B _11640_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _11641_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14360_ _14364_/A _14360_/B vssd1 vssd1 vccd1 vccd1 _17979_/D sky130_fd_sc_hd__and2_1
X_11572_ hold5428/X _11195_/B _11571_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _11572_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13311_ _13311_/A1 _13309_/X _13310_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13311_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput19 input19/A vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_2
X_10523_ hold2958/X _16665_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10524_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_181_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14291_ hold2183/X _14333_/A2 _14290_/X _13895_/A vssd1 vssd1 vccd1 vccd1 _14291_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16030_ _18409_/CLK _16030_/D vssd1 vssd1 vccd1 vccd1 hold830/A sky130_fd_sc_hd__dfxtp_1
X_13242_ _17581_/Q _17115_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13242_/X sky130_fd_sc_hd__mux2_1
X_10454_ hold2058/X hold4482/X _10646_/C vssd1 vssd1 vccd1 vccd1 _10455_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13173_ _13172_/X hold4340/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13173_/X sky130_fd_sc_hd__mux2_1
X_10385_ hold2544/X _16619_/Q _10385_/S vssd1 vssd1 vccd1 vccd1 _10386_/B sky130_fd_sc_hd__mux2_1
X_12124_ hold5456/X _12323_/B _12123_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _12124_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17981_ _17981_/CLK _17981_/D vssd1 vssd1 vccd1 vccd1 _17981_/Q sky130_fd_sc_hd__dfxtp_1
X_12055_ hold4030/X _12365_/B _12054_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _12055_/X
+ sky130_fd_sc_hd__o211a_1
X_16932_ _18428_/CLK _16932_/D vssd1 vssd1 vccd1 vccd1 _16932_/Q sky130_fd_sc_hd__dfxtp_1
X_11006_ hold1027/X _16826_/Q _11213_/C vssd1 vssd1 vccd1 vccd1 _11007_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_217_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16863_ _18066_/CLK _16863_/D vssd1 vssd1 vccd1 vccd1 _16863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15814_ _17690_/CLK _15814_/D vssd1 vssd1 vccd1 vccd1 _15814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16794_ _17997_/CLK _16794_/D vssd1 vssd1 vccd1 vccd1 _16794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_232_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15745_ _17716_/CLK _15745_/D vssd1 vssd1 vccd1 vccd1 _15745_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _14358_/A _12957_/B vssd1 vssd1 vccd1 vccd1 _17495_/D sky130_fd_sc_hd__and2_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11908_ hold4873/X _12308_/B _11907_/X _08167_/A vssd1 vssd1 vccd1 vccd1 _11908_/X
+ sky130_fd_sc_hd__o211a_1
X_15676_ _17229_/CLK _15676_/D vssd1 vssd1 vccd1 vccd1 _15676_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _12888_/A _12888_/B vssd1 vssd1 vccd1 vccd1 _17472_/D sky130_fd_sc_hd__and2_1
XFILLER_0_201_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17415_ _17430_/CLK _17415_/D vssd1 vssd1 vccd1 vccd1 _17415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14627_ _14627_/A _15182_/B vssd1 vssd1 vccd1 vccd1 _14672_/B sky130_fd_sc_hd__or2_4
X_18395_ _18395_/CLK _18395_/D vssd1 vssd1 vccd1 vccd1 _18395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11839_ hold5380/X _12323_/B _11838_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _11839_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17346_ _17347_/CLK hold45/X vssd1 vssd1 vccd1 vccd1 _17346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14558_ _15492_/A _14573_/B _18074_/Q vssd1 vssd1 vccd1 vccd1 _14558_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13509_ _13800_/A _13509_/B vssd1 vssd1 vccd1 vccd1 _13509_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17277_ _17277_/CLK _17277_/D vssd1 vssd1 vccd1 vccd1 _17277_/Q sky130_fd_sc_hd__dfxtp_1
X_14489_ _15169_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14489_/X sky130_fd_sc_hd__or2_1
XFILLER_0_141_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16228_ _18458_/CLK _16228_/D vssd1 vssd1 vccd1 vccd1 _16228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4107 _17353_/Q vssd1 vssd1 vccd1 vccd1 hold4107/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_401_wb_clk_i clkbuf_6_37_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17825_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16159_ _17500_/CLK _16159_/D vssd1 vssd1 vccd1 vccd1 _16159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4118 _10744_/X vssd1 vssd1 vccd1 vccd1 _16738_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4129 _17685_/Q vssd1 vssd1 vccd1 vccd1 hold4129/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3406 hold4527/X vssd1 vssd1 vccd1 vccd1 _10604_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08981_ hold92/X _16108_/Q _08991_/S vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__mux2_1
Xhold3417 hold6117/X vssd1 vssd1 vccd1 vccd1 hold3417/X sky130_fd_sc_hd__buf_2
Xhold3428 _16520_/Q vssd1 vssd1 vccd1 vccd1 hold3428/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_228_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3439 _16352_/Q vssd1 vssd1 vccd1 vccd1 _13286_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2705 _15669_/Q vssd1 vssd1 vccd1 vccd1 hold2705/X sky130_fd_sc_hd__dlygate4sd3_1
X_07932_ _15555_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07932_/X sky130_fd_sc_hd__or2_1
Xhold2716 _15863_/Q vssd1 vssd1 vccd1 vccd1 hold2716/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2727 _18214_/Q vssd1 vssd1 vccd1 vccd1 hold2727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2738 _14593_/X vssd1 vssd1 vccd1 vccd1 _18090_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2749 _15740_/Q vssd1 vssd1 vccd1 vccd1 hold2749/X sky130_fd_sc_hd__dlygate4sd3_1
X_07863_ _15215_/A _07865_/B vssd1 vssd1 vccd1 vccd1 _07863_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_78_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09602_ hold2185/X _16358_/Q _09992_/C vssd1 vssd1 vccd1 vccd1 _09603_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_3_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07794_ _11158_/A _07794_/B vssd1 vssd1 vccd1 vccd1 _18461_/D sky130_fd_sc_hd__nor2_1
X_09533_ hold2369/X _13150_/A _10964_/S vssd1 vssd1 vccd1 vccd1 _09534_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_78_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09464_ _09463_/A _09461_/X _09478_/B vssd1 vssd1 vccd1 vccd1 _09465_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08415_ _15529_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08415_/X sky130_fd_sc_hd__or2_1
XFILLER_0_148_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09395_ _12412_/A _09395_/B vssd1 vssd1 vccd1 vccd1 _16284_/D sky130_fd_sc_hd__and2_1
XFILLER_0_148_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08346_ _14850_/A hold2718/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08347_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_19_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08277_ hold1568/X _08268_/B _08276_/X _12753_/A vssd1 vssd1 vccd1 vccd1 _08277_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6010 _17553_/Q vssd1 vssd1 vccd1 vccd1 hold6010/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6021 _17532_/Q vssd1 vssd1 vccd1 vccd1 hold6021/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6032 _17531_/Q vssd1 vssd1 vccd1 vccd1 hold6032/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6043 data_in[25] vssd1 vssd1 vccd1 vccd1 hold435/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6054 _18250_/Q vssd1 vssd1 vccd1 vccd1 hold6054/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_225_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6065 _18370_/Q vssd1 vssd1 vccd1 vccd1 hold6065/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5320 _13549_/X vssd1 vssd1 vccd1 vccd1 _17636_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_142_wb_clk_i clkbuf_6_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17535_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold6076 _18275_/Q vssd1 vssd1 vccd1 vccd1 hold6076/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5331 _17154_/Q vssd1 vssd1 vccd1 vccd1 hold5331/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6087 data_in[12] vssd1 vssd1 vccd1 vccd1 hold247/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5342 _13375_/X vssd1 vssd1 vccd1 vccd1 _17578_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5353 _16800_/Q vssd1 vssd1 vccd1 vccd1 hold5353/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6098 la_data_in[29] vssd1 vssd1 vccd1 vccd1 hold506/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5364 _16804_/Q vssd1 vssd1 vccd1 vccd1 hold5364/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4630 _17600_/Q vssd1 vssd1 vccd1 vccd1 hold4630/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5375 _11533_/X vssd1 vssd1 vccd1 vccd1 _17001_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4641 _09793_/X vssd1 vssd1 vccd1 vccd1 _16421_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10170_ _10554_/A _10170_/B vssd1 vssd1 vccd1 vccd1 _10170_/X sky130_fd_sc_hd__or2_1
Xhold5386 _17707_/Q vssd1 vssd1 vccd1 vccd1 hold5386/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4652 _16490_/Q vssd1 vssd1 vccd1 vccd1 hold4652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5397 _13678_/X vssd1 vssd1 vccd1 vccd1 _17679_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4663 _09880_/X vssd1 vssd1 vccd1 vccd1 _16450_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4674 _16904_/Q vssd1 vssd1 vccd1 vccd1 hold4674/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3940 _16686_/Q vssd1 vssd1 vccd1 vccd1 hold3940/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4685 _17663_/Q vssd1 vssd1 vccd1 vccd1 hold4685/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3951 _09874_/X vssd1 vssd1 vccd1 vccd1 _16448_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4696 _11974_/X vssd1 vssd1 vccd1 vccd1 _17148_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3962 _17726_/Q vssd1 vssd1 vccd1 vccd1 _13817_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3973 _10171_/X vssd1 vssd1 vccd1 vccd1 _16547_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_238_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3984 _16687_/Q vssd1 vssd1 vccd1 vccd1 hold3984/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout152 hold2272/X vssd1 vssd1 vccd1 vccd1 _12851_/S sky130_fd_sc_hd__buf_6
Xfanout163 _13817_/B vssd1 vssd1 vccd1 vccd1 _12293_/B sky130_fd_sc_hd__buf_2
Xhold3995 _16589_/Q vssd1 vssd1 vccd1 vccd1 hold3995/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout174 fanout210/X vssd1 vssd1 vccd1 vccd1 _11717_/B sky130_fd_sc_hd__clkbuf_4
Xfanout185 _13868_/B vssd1 vssd1 vccd1 vccd1 _13871_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout196 _12365_/B vssd1 vssd1 vccd1 vccd1 _13886_/B sky130_fd_sc_hd__buf_4
X_13860_ hold4458/X _13788_/A _13859_/X vssd1 vssd1 vccd1 vccd1 _13860_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_198_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12811_ hold1666/X _17448_/Q _12811_/S vssd1 vssd1 vccd1 vccd1 _12811_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13791_ _13791_/A _13791_/B vssd1 vssd1 vccd1 vccd1 _13791_/X sky130_fd_sc_hd__or2_1
XFILLER_0_215_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ hold2904/X _15547_/B _15529_/X _12822_/A vssd1 vssd1 vccd1 vccd1 _15530_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _16245_/Q _17425_/Q _12811_/S vssd1 vssd1 vccd1 vccd1 _12742_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15461_ hold775/X _09362_/D _09392_/D hold457/X _15460_/X vssd1 vssd1 vccd1 vccd1
+ _15462_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_182_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ hold2000/X _17402_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _12673_/X sky130_fd_sc_hd__mux2_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17200_ _17229_/CLK _17200_/D vssd1 vssd1 vccd1 vccd1 _17200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ hold2123/X hold4179/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11625_/B sky130_fd_sc_hd__mux2_1
X_14412_ hold3091/X _14446_/A2 _14411_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _14412_/X
+ sky130_fd_sc_hd__o211a_1
X_18180_ _18180_/CLK _18180_/D vssd1 vssd1 vccd1 vccd1 _18180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15392_ _15480_/A _15392_/B _15392_/C _15392_/D vssd1 vssd1 vccd1 vccd1 _15392_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17131_ _17878_/CLK _17131_/D vssd1 vssd1 vccd1 vccd1 _17131_/Q sky130_fd_sc_hd__dfxtp_1
X_14343_ hold915/X hold1620/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14344_/B sky130_fd_sc_hd__mux2_1
X_11555_ hold1393/X hold5127/X _11654_/S vssd1 vssd1 vccd1 vccd1 _11556_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_208_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10506_ _10542_/A _10506_/B vssd1 vssd1 vccd1 vccd1 _10506_/X sky130_fd_sc_hd__or2_1
X_14274_ _15169_/A _14282_/B vssd1 vssd1 vccd1 vccd1 _14274_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17062_ _17910_/CLK _17062_/D vssd1 vssd1 vccd1 vccd1 _17062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11486_ hold1742/X hold4020/X _12242_/S vssd1 vssd1 vccd1 vccd1 _11487_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_122_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13225_ _13225_/A _13225_/B vssd1 vssd1 vccd1 vccd1 _13225_/X sky130_fd_sc_hd__and2_1
X_16013_ _18423_/CLK _16013_/D vssd1 vssd1 vccd1 vccd1 hold154/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10437_ _11103_/A _10437_/B vssd1 vssd1 vccd1 vccd1 _10437_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13156_ hold3523/X _13155_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13156_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10368_ _10482_/A _10368_/B vssd1 vssd1 vccd1 vccd1 _10368_/X sky130_fd_sc_hd__or2_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ hold3053/X _17193_/Q _12299_/C vssd1 vssd1 vccd1 vccd1 _12108_/B sky130_fd_sc_hd__mux2_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13087_ _13199_/A1 _13085_/X _13086_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13087_/X
+ sky130_fd_sc_hd__o211a_1
X_17964_ _17964_/CLK _17964_/D vssd1 vssd1 vccd1 vccd1 _17964_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ _10413_/A _10299_/B vssd1 vssd1 vccd1 vccd1 _10299_/X sky130_fd_sc_hd__or2_1
XFILLER_0_236_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12038_ hold2433/X hold5731/X _12362_/C vssd1 vssd1 vccd1 vccd1 _12039_/B sky130_fd_sc_hd__mux2_1
X_16915_ _17892_/CLK _16915_/D vssd1 vssd1 vccd1 vccd1 _16915_/Q sky130_fd_sc_hd__dfxtp_1
X_17895_ _17895_/CLK _17895_/D vssd1 vssd1 vccd1 vccd1 _17895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_233_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16846_ _18049_/CLK _16846_/D vssd1 vssd1 vccd1 vccd1 _16846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16777_ _18461_/CLK _16777_/D vssd1 vssd1 vccd1 vccd1 _16777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13989_ hold1676/X _13986_/B _13988_/X _14131_/C1 vssd1 vssd1 vccd1 vccd1 _13989_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15728_ _17697_/CLK _15728_/D vssd1 vssd1 vccd1 vccd1 _15728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18447_ _18447_/CLK _18447_/D vssd1 vssd1 vccd1 vccd1 _18447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15659_ _17897_/CLK _15659_/D vssd1 vssd1 vccd1 vccd1 _15659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08200_ hold2790/X _08213_/B _08199_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08200_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09180_ _15509_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09180_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18378_ _18378_/CLK _18378_/D vssd1 vssd1 vccd1 vccd1 _18378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08131_ _08131_/A _08131_/B vssd1 vssd1 vccd1 vccd1 _15704_/D sky130_fd_sc_hd__and2_1
XFILLER_0_83_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17329_ _18405_/CLK hold60/X vssd1 vssd1 vccd1 vccd1 _17329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08062_ _15521_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08062_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3203 _10074_/Y vssd1 vssd1 vccd1 vccd1 _10075_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3214 _16495_/Q vssd1 vssd1 vccd1 vccd1 hold3214/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3225 _09559_/X vssd1 vssd1 vccd1 vccd1 _16343_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3236 _12575_/X vssd1 vssd1 vccd1 vccd1 _12576_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_228_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3247 _16555_/Q vssd1 vssd1 vccd1 vccd1 hold3247/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2502 _14486_/X vssd1 vssd1 vccd1 vccd1 _18040_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08964_ _15434_/A _08964_/B vssd1 vssd1 vccd1 vccd1 _16099_/D sky130_fd_sc_hd__and2_1
Xhold3258 _10402_/X vssd1 vssd1 vccd1 vccd1 _16624_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2513 _07925_/X vssd1 vssd1 vccd1 vccd1 _15606_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2524 _16231_/Q vssd1 vssd1 vccd1 vccd1 hold2524/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3269 _12611_/X vssd1 vssd1 vccd1 vccd1 _12612_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2535 _15112_/X vssd1 vssd1 vccd1 vccd1 _18340_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1801 _18232_/Q vssd1 vssd1 vccd1 vccd1 hold1801/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2546 _18070_/Q vssd1 vssd1 vccd1 vccd1 hold2546/X sky130_fd_sc_hd__dlygate4sd3_1
X_07915_ hold1556/X _07918_/B _07914_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _07915_/X
+ sky130_fd_sc_hd__o211a_1
X_08895_ _15324_/A _08895_/B vssd1 vssd1 vccd1 vccd1 _16065_/D sky130_fd_sc_hd__and2_1
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1812 _13008_/X vssd1 vssd1 vccd1 vccd1 _17512_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2557 _16221_/Q vssd1 vssd1 vccd1 vccd1 hold2557/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1823 _16217_/Q vssd1 vssd1 vccd1 vccd1 hold1823/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2568 _07907_/X vssd1 vssd1 vccd1 vccd1 _15597_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1834 _15130_/X vssd1 vssd1 vccd1 vccd1 _18348_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2579 _18308_/Q vssd1 vssd1 vccd1 vccd1 hold2579/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1845 _18199_/Q vssd1 vssd1 vccd1 vccd1 hold1845/X sky130_fd_sc_hd__dlygate4sd3_1
X_07846_ hold1039/X _07869_/B _07845_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _07846_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1856 _14508_/X vssd1 vssd1 vccd1 vccd1 _18050_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1867 _18042_/Q vssd1 vssd1 vccd1 vccd1 hold1867/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1878 _08178_/X vssd1 vssd1 vccd1 vccd1 _15725_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1889 _18121_/Q vssd1 vssd1 vccd1 vccd1 hold1889/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09516_ _09984_/A _09516_/B vssd1 vssd1 vccd1 vccd1 _09516_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09447_ _09447_/A _09447_/B _09447_/C _09447_/D vssd1 vssd1 vccd1 vccd1 _09456_/D
+ sky130_fd_sc_hd__and4_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_394_wb_clk_i clkbuf_6_36_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17900_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09378_ _15936_/Q _15448_/A2 _09386_/D hold547/X vssd1 vssd1 vccd1 vccd1 _09378_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08329_ _15553_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08329_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_323_wb_clk_i clkbuf_6_46_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17907_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_151_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11340_ _11631_/A _11340_/B vssd1 vssd1 vccd1 vccd1 _11340_/X sky130_fd_sc_hd__or2_1
XFILLER_0_201_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11271_ _11658_/A _11271_/B vssd1 vssd1 vccd1 vccd1 _11271_/X sky130_fd_sc_hd__or2_1
X_13010_ hold1635/X _13003_/Y _13009_/X _14358_/A vssd1 vssd1 vccd1 vccd1 _13010_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5150 _17648_/Q vssd1 vssd1 vccd1 vccd1 hold5150/X sky130_fd_sc_hd__dlygate4sd3_1
X_10222_ hold4504/X _10604_/B _10221_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _10222_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5161 _17050_/Q vssd1 vssd1 vccd1 vccd1 hold5161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5172 _12277_/X vssd1 vssd1 vccd1 vccd1 _17249_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5183 _16983_/Q vssd1 vssd1 vccd1 vccd1 hold5183/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5194 _13777_/X vssd1 vssd1 vccd1 vccd1 _17712_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4460 _13861_/Y vssd1 vssd1 vccd1 vccd1 _17740_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10153_ hold3799/X _10631_/B _10152_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10153_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4471 _17099_/Q vssd1 vssd1 vccd1 vccd1 hold4471/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4482 _16642_/Q vssd1 vssd1 vccd1 vccd1 hold4482/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4493 _16606_/Q vssd1 vssd1 vccd1 vccd1 hold4493/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3770 _12764_/X vssd1 vssd1 vccd1 vccd1 _12765_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3781 _16627_/Q vssd1 vssd1 vccd1 vccd1 hold3781/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10084_ hold3740/X _10598_/B _10083_/X _15019_/C1 vssd1 vssd1 vccd1 vccd1 _10084_/X
+ sky130_fd_sc_hd__o211a_1
X_14961_ hold1299/X _14952_/B _14960_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _14961_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3792 _11050_/X vssd1 vssd1 vccd1 vccd1 _16840_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__buf_4
XTAP_5965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16700_ _18162_/CLK _16700_/D vssd1 vssd1 vccd1 vccd1 _16700_/Q sky130_fd_sc_hd__dfxtp_1
X_13912_ _14413_/A hold2930/X hold297/X vssd1 vssd1 vccd1 vccd1 _13913_/B sky130_fd_sc_hd__mux2_1
XTAP_5987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17680_ _17744_/CLK _17680_/D vssd1 vssd1 vccd1 vccd1 _17680_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14892_ _15231_/A _14892_/B vssd1 vssd1 vccd1 vccd1 _14892_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16631_ _18221_/CLK _16631_/D vssd1 vssd1 vccd1 vccd1 _16631_/Q sky130_fd_sc_hd__dfxtp_1
X_13843_ _13873_/A _13843_/B vssd1 vssd1 vccd1 vccd1 _13843_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_230_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16562_ _18124_/CLK _16562_/D vssd1 vssd1 vccd1 vccd1 _16562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10986_ _10986_/A _10986_/B vssd1 vssd1 vccd1 vccd1 _10986_/X sky130_fd_sc_hd__or2_1
X_13774_ hold5492/X _13871_/B _13773_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13774_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18301_ _18375_/CLK _18301_/D vssd1 vssd1 vccd1 vccd1 _18301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15513_ _15513_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15513_/X sky130_fd_sc_hd__or2_1
X_12725_ hold3400/X _12724_/X _12812_/S vssd1 vssd1 vccd1 vccd1 _12725_/X sky130_fd_sc_hd__mux2_1
X_16493_ _18334_/CLK _16493_/D vssd1 vssd1 vccd1 vccd1 _16493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18232_ _18232_/CLK _18232_/D vssd1 vssd1 vccd1 vccd1 _18232_/Q sky130_fd_sc_hd__dfxtp_1
X_15444_ _15473_/A _15444_/B vssd1 vssd1 vccd1 vccd1 _18420_/D sky130_fd_sc_hd__and2_1
XFILLER_0_183_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12656_ hold3143/X _12655_/X _12851_/S vssd1 vssd1 vccd1 vccd1 _12656_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_143_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18163_ _18227_/CLK _18163_/D vssd1 vssd1 vccd1 vccd1 _18163_/Q sky130_fd_sc_hd__dfxtp_1
X_11607_ _11697_/A _11607_/B vssd1 vssd1 vccd1 vccd1 _11607_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15375_ hold400/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15375_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12587_ hold3131/X _12586_/X _12923_/S vssd1 vssd1 vccd1 vccd1 _12587_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_142_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17114_ _17576_/CLK _17114_/D vssd1 vssd1 vccd1 vccd1 _17114_/Q sky130_fd_sc_hd__dfxtp_1
X_14326_ _15221_/A _14326_/B vssd1 vssd1 vccd1 vccd1 _14326_/Y sky130_fd_sc_hd__nand2_1
X_18094_ _18200_/CLK _18094_/D vssd1 vssd1 vccd1 vccd1 _18094_/Q sky130_fd_sc_hd__dfxtp_1
X_11538_ _11631_/A _11538_/B vssd1 vssd1 vccd1 vccd1 _11538_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold408 hold408/A vssd1 vssd1 vccd1 vccd1 hold408/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 hold419/A vssd1 vssd1 vccd1 vccd1 hold419/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17045_ _17861_/CLK _17045_/D vssd1 vssd1 vccd1 vccd1 _17045_/Q sky130_fd_sc_hd__dfxtp_1
X_14257_ hold1670/X _14272_/B _14256_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14257_/X
+ sky130_fd_sc_hd__o211a_1
X_11469_ _11661_/A _11469_/B vssd1 vssd1 vccd1 vccd1 _11469_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13208_ _13201_/X _13207_/X _13296_/B1 vssd1 vssd1 vccd1 vccd1 _17544_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_237_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14188_ _15207_/A _14204_/B vssd1 vssd1 vccd1 vccd1 _14188_/X sky130_fd_sc_hd__or2_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13139_ _13138_/X hold6002/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13139_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_238_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 _15149_/X vssd1 vssd1 vccd1 vccd1 hold1108/X sky130_fd_sc_hd__dlygate4sd3_1
X_17947_ _18045_/CLK _17947_/D vssd1 vssd1 vccd1 vccd1 _17947_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1119 _17750_/Q vssd1 vssd1 vccd1 vccd1 hold1119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08680_ _12426_/A hold852/X vssd1 vssd1 vccd1 vccd1 _15961_/D sky130_fd_sc_hd__and2_1
XFILLER_0_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17878_ _17878_/CLK _17878_/D vssd1 vssd1 vccd1 vccd1 _17878_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_6_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_215_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16829_ _17973_/CLK _16829_/D vssd1 vssd1 vccd1 vccd1 _16829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09301_ hold933/X _09337_/B vssd1 vssd1 vccd1 vccd1 _09301_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09232_ hold113/X hold363/A vssd1 vssd1 vccd1 vccd1 hold364/A sky130_fd_sc_hd__or2_1
XFILLER_0_75_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09163_ hold2479/X _09164_/B _09162_/Y _12906_/A vssd1 vssd1 vccd1 vccd1 _09163_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08114_ _15085_/A hold1015/X hold108/X vssd1 vssd1 vccd1 vccd1 _08114_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09094_ _15535_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09094_/X sky130_fd_sc_hd__or2_1
XFILLER_0_71_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08045_ _14732_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08045_/X sky130_fd_sc_hd__or2_1
Xhold920 hold920/A vssd1 vssd1 vccd1 vccd1 hold920/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold931 input66/X vssd1 vssd1 vccd1 vccd1 hold931/X sky130_fd_sc_hd__buf_1
XFILLER_0_222_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold942 hold942/A vssd1 vssd1 vccd1 vccd1 hold942/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold953 hold953/A vssd1 vssd1 vccd1 vccd1 hold953/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 hold964/A vssd1 vssd1 vccd1 vccd1 hold964/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 hold975/A vssd1 vssd1 vccd1 vccd1 input63/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3000 _16205_/Q vssd1 vssd1 vccd1 vccd1 hold3000/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold986 hold986/A vssd1 vssd1 vccd1 vccd1 hold986/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3011 _09147_/X vssd1 vssd1 vccd1 vccd1 _16186_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3022 _09159_/X vssd1 vssd1 vccd1 vccd1 _16192_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3033 _18087_/Q vssd1 vssd1 vccd1 vccd1 hold3033/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold997 hold997/A vssd1 vssd1 vccd1 vccd1 hold997/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09996_ _13102_/A _09984_/A _09995_/X vssd1 vssd1 vccd1 vccd1 _09997_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3044 _07864_/X vssd1 vssd1 vccd1 vccd1 _15577_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3055 _16262_/Q vssd1 vssd1 vccd1 vccd1 hold3055/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2310 _15617_/Q vssd1 vssd1 vccd1 vccd1 hold2310/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3066 _14933_/X vssd1 vssd1 vccd1 vccd1 _18253_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2321 _08510_/X vssd1 vssd1 vccd1 vccd1 _15882_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3077 _08412_/X vssd1 vssd1 vccd1 vccd1 _15836_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2332 _15518_/X vssd1 vssd1 vccd1 vccd1 _18437_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08947_ hold29/X hold667/X _08991_/S vssd1 vssd1 vccd1 vccd1 _08948_/B sky130_fd_sc_hd__mux2_1
Xhold3088 _15202_/X vssd1 vssd1 vccd1 vccd1 _18383_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2343 _15871_/Q vssd1 vssd1 vccd1 vccd1 hold2343/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3099 _18304_/Q vssd1 vssd1 vccd1 vccd1 hold3099/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2354 _14542_/X vssd1 vssd1 vccd1 vccd1 _18067_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1620 _17971_/Q vssd1 vssd1 vccd1 vccd1 hold1620/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2365 _15565_/Q vssd1 vssd1 vccd1 vccd1 hold2365/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2376 _18202_/Q vssd1 vssd1 vccd1 vccd1 hold2376/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1631 _07880_/X vssd1 vssd1 vccd1 vccd1 _15585_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2387 _08487_/X vssd1 vssd1 vccd1 vccd1 _15872_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1642 _09167_/X vssd1 vssd1 vccd1 vccd1 _16196_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1653 _14631_/X vssd1 vssd1 vccd1 vccd1 _18108_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08878_ hold71/X hold772/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08879_/B sky130_fd_sc_hd__mux2_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2398 _15743_/Q vssd1 vssd1 vccd1 vccd1 hold2398/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1664 _15610_/Q vssd1 vssd1 vccd1 vccd1 hold1664/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1675 _14307_/X vssd1 vssd1 vccd1 vccd1 _17953_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1686 _15654_/Q vssd1 vssd1 vccd1 vccd1 hold1686/X sky130_fd_sc_hd__dlygate4sd3_1
X_07829_ hold330/X hold355/X vssd1 vssd1 vccd1 vccd1 _07829_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_169_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1697 _09330_/X vssd1 vssd1 vccd1 vccd1 _16275_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10840_ hold5398/X _11789_/B _10839_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _10840_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_233_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10771_ hold4616/X _11153_/B _10770_/X _14552_/C1 vssd1 vssd1 vccd1 vccd1 _10771_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12510_ _14556_/A _12510_/B vssd1 vssd1 vccd1 vccd1 _12510_/Y sky130_fd_sc_hd__nor2_1
X_13490_ hold1450/X hold5325/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13491_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_165_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12441_ hold320/X hold866/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12442_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_136_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_212_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15160_ hold2211/X _15167_/B _15159_/X _15160_/C1 vssd1 vssd1 vccd1 vccd1 _15160_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12372_ hold3505/X _12273_/A _12371_/X vssd1 vssd1 vccd1 vccd1 _12372_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11323_ hold5500/X _12335_/B _11322_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _11323_/X
+ sky130_fd_sc_hd__o211a_1
X_14111_ hold1596/X _14148_/B _14110_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _14111_/X
+ sky130_fd_sc_hd__o211a_1
X_15091_ _15145_/A _15119_/B vssd1 vssd1 vccd1 vccd1 _15091_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11254_ hold5293/X _11732_/B _11253_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _11254_/X
+ sky130_fd_sc_hd__o211a_1
X_14042_ _14543_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14042_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10205_ hold2681/X _16559_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10206_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11185_ _11218_/A _11185_/B vssd1 vssd1 vccd1 vccd1 _11185_/Y sky130_fd_sc_hd__nor2_1
XTAP_6441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4290 _17106_/Q vssd1 vssd1 vccd1 vccd1 hold4290/X sky130_fd_sc_hd__dlygate4sd3_1
X_17801_ _17894_/CLK _17801_/D vssd1 vssd1 vccd1 vccd1 _17801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10136_ hold2115/X hold3515/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10137_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_238_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_235_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15993_ _18400_/CLK _15993_/D vssd1 vssd1 vccd1 vccd1 hold870/A sky130_fd_sc_hd__dfxtp_1
XTAP_5751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17732_ _17732_/CLK _17732_/D vssd1 vssd1 vccd1 vccd1 _17732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10067_ _10067_/A _10067_/B _10067_/C vssd1 vssd1 vccd1 vccd1 _10067_/X sky130_fd_sc_hd__and3_1
X_14944_ _15213_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14944_/X sky130_fd_sc_hd__or2_1
XTAP_5784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17663_ _17729_/CLK _17663_/D vssd1 vssd1 vccd1 vccd1 _17663_/Q sky130_fd_sc_hd__dfxtp_1
X_14875_ hold2207/X hold332/X _14874_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14875_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16614_ _18172_/CLK _16614_/D vssd1 vssd1 vccd1 vccd1 _16614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13826_ _17729_/Q _13862_/B _13862_/C vssd1 vssd1 vccd1 vccd1 _13826_/X sky130_fd_sc_hd__and3_1
X_17594_ _17626_/CLK _17594_/D vssd1 vssd1 vccd1 vccd1 _17594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_245_wb_clk_i clkbuf_6_57_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18156_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16545_ _18232_/CLK _16545_/D vssd1 vssd1 vccd1 vccd1 _16545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13757_ hold1307/X _17706_/Q _13874_/C vssd1 vssd1 vccd1 vccd1 _13758_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_156_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10969_ hold4821/X _11162_/B _10968_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _10969_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12708_ _12786_/A _12708_/B vssd1 vssd1 vccd1 vccd1 _17412_/D sky130_fd_sc_hd__and2_1
X_16476_ _18389_/CLK _16476_/D vssd1 vssd1 vccd1 vccd1 _16476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13688_ hold1538/X hold5337/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13689_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_73_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18215_ _18215_/CLK _18215_/D vssd1 vssd1 vccd1 vccd1 _18215_/Q sky130_fd_sc_hd__dfxtp_1
X_15427_ _16095_/Q _09392_/B _09392_/C hold346/X vssd1 vssd1 vccd1 vccd1 _15427_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12639_ _12849_/A _12639_/B vssd1 vssd1 vccd1 vccd1 _17389_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18146_ _18146_/CLK _18146_/D vssd1 vssd1 vccd1 vccd1 _18146_/Q sky130_fd_sc_hd__dfxtp_1
X_15358_ hold455/X _09386_/A _15441_/A2 hold701/X vssd1 vssd1 vccd1 vccd1 _15358_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_198_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5908 _18411_/Q vssd1 vssd1 vccd1 vccd1 hold5908/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold205 hold205/A vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5919 _18402_/Q vssd1 vssd1 vccd1 vccd1 hold5919/X sky130_fd_sc_hd__dlygate4sd3_1
X_14309_ hold2969/X _14333_/A2 _14308_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _14309_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18077_ _18265_/CLK _18077_/D vssd1 vssd1 vccd1 vccd1 _18077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15289_ hold205/X _15485_/A2 _15488_/A2 hold292/X _15288_/X vssd1 vssd1 vccd1 vccd1
+ _15292_/C sky130_fd_sc_hd__a221o_1
Xhold216 hold216/A vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 hold227/A vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold238 hold481/X vssd1 vssd1 vccd1 vccd1 hold482/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold249 input8/X vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__buf_1
X_17028_ _17908_/CLK _17028_/D vssd1 vssd1 vccd1 vccd1 _17028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout707 _09047_/A vssd1 vssd1 vccd1 vccd1 _15374_/A sky130_fd_sc_hd__clkbuf_4
X_09850_ hold3880/X _11204_/B _09849_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _09850_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout718 _12412_/A vssd1 vssd1 vccd1 vccd1 _15314_/A sky130_fd_sc_hd__clkbuf_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout729 _09003_/A vssd1 vssd1 vccd1 vccd1 _12420_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_237_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ hold131/X hold431/X _08801_/S vssd1 vssd1 vccd1 vccd1 hold432/A sky130_fd_sc_hd__mux2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ hold3773/X _10067_/B _09780_/X _15228_/C1 vssd1 vssd1 vccd1 vccd1 _09781_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _15491_/A hold758/X vssd1 vssd1 vccd1 vccd1 _15986_/D sky130_fd_sc_hd__and2_1
XFILLER_0_217_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08663_ _17519_/Q hold937/X vssd1 vssd1 vccd1 vccd1 _12380_/B sky130_fd_sc_hd__or2_1
XFILLER_0_240_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08594_ hold278/X hold490/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold491/A sky130_fd_sc_hd__mux2_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09215_ hold2754/X _09214_/B _09214_/Y _12837_/A vssd1 vssd1 vccd1 vccd1 _09215_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09146_ _15529_/A _09156_/B vssd1 vssd1 vccd1 vccd1 _09146_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09077_ hold2382/X _09106_/B _09076_/X _12987_/A vssd1 vssd1 vccd1 vccd1 _09077_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08028_ hold2338/X _08029_/B _08027_/Y _08137_/A vssd1 vssd1 vccd1 vccd1 _08028_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_49_wb_clk_i clkbuf_6_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17820_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_163_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold750 hold750/A vssd1 vssd1 vccd1 vccd1 hold750/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold761 hold761/A vssd1 vssd1 vccd1 vccd1 hold761/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 hold772/A vssd1 vssd1 vccd1 vccd1 hold772/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 hold783/A vssd1 vssd1 vccd1 vccd1 hold783/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 hold794/A vssd1 vssd1 vccd1 vccd1 hold794/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_229_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_228_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09979_ hold3597/X _10046_/B _09978_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09979_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2140 _14289_/X vssd1 vssd1 vccd1 vccd1 _17944_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2151 _17959_/Q vssd1 vssd1 vccd1 vccd1 hold2151/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2162 _14779_/X vssd1 vssd1 vccd1 vccd1 _18180_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2173 _15659_/Q vssd1 vssd1 vccd1 vccd1 hold2173/X sky130_fd_sc_hd__dlygate4sd3_1
X_12990_ _15244_/A _12990_/B vssd1 vssd1 vccd1 vccd1 _17506_/D sky130_fd_sc_hd__and2_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2184 _14291_/X vssd1 vssd1 vccd1 vccd1 _17945_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2195 _18049_/Q vssd1 vssd1 vccd1 vccd1 hold2195/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1450 _15802_/Q vssd1 vssd1 vccd1 vccd1 hold1450/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1461 _18175_/Q vssd1 vssd1 vccd1 vccd1 hold1461/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1472 _08281_/X vssd1 vssd1 vccd1 vccd1 _15775_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11941_ hold5345/X _12329_/B _11940_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11941_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_231_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1483 _18296_/Q vssd1 vssd1 vccd1 vccd1 hold1483/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1494 _09421_/X vssd1 vssd1 vccd1 vccd1 _16296_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _15215_/A _14664_/B vssd1 vssd1 vccd1 vccd1 _14660_/Y sky130_fd_sc_hd__nand2_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ hold5799/X _12350_/B _11871_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _11872_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_6_37_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_37_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _13719_/A _13611_/B vssd1 vssd1 vccd1 vccd1 _13611_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ hold1583/X _16765_/Q _11660_/S vssd1 vssd1 vccd1 vccd1 _10824_/B sky130_fd_sc_hd__mux2_1
X_14591_ hold2282/X _14610_/B _14590_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14591_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16330_ _18371_/CLK _16330_/D vssd1 vssd1 vccd1 vccd1 _16330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13542_ _13734_/A _13542_/B vssd1 vssd1 vccd1 vccd1 _13542_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10754_ hold2183/X _16742_/Q _11723_/C vssd1 vssd1 vccd1 vccd1 _10755_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_211_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16261_ _17378_/CLK _16261_/D vssd1 vssd1 vccd1 vccd1 _16261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13473_ _13752_/A _13473_/B vssd1 vssd1 vccd1 vccd1 _13473_/X sky130_fd_sc_hd__or2_1
X_10685_ hold2635/X hold4309/X _11654_/S vssd1 vssd1 vccd1 vccd1 _10686_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18000_ _18059_/CLK _18000_/D vssd1 vssd1 vccd1 vccd1 _18000_/Q sky130_fd_sc_hd__dfxtp_1
X_15212_ hold6077/X _15219_/B hold377/X _15212_/C1 vssd1 vssd1 vccd1 vccd1 hold378/A
+ sky130_fd_sc_hd__o211a_1
X_12424_ _15324_/A _12424_/B vssd1 vssd1 vccd1 vccd1 _17305_/D sky130_fd_sc_hd__and2_1
XFILLER_0_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16192_ _17881_/CLK _16192_/D vssd1 vssd1 vccd1 vccd1 _16192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15143_ _15197_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15143_/X sky130_fd_sc_hd__or2_1
XFILLER_0_152_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12355_ _13819_/A _12355_/B vssd1 vssd1 vccd1 vccd1 _12355_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_168_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11306_ _17774_/Q _16926_/Q _11783_/C vssd1 vssd1 vccd1 vccd1 _11307_/B sky130_fd_sc_hd__mux2_1
X_15074_ hold338/X _15182_/B vssd1 vssd1 vccd1 vccd1 _15119_/B sky130_fd_sc_hd__or2_4
XFILLER_0_132_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12286_ hold5068/X _12317_/B _12285_/X _14211_/C1 vssd1 vssd1 vccd1 vccd1 _12286_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11237_ hold2223/X hold3704/X _11717_/C vssd1 vssd1 vccd1 vccd1 _11238_/B sky130_fd_sc_hd__mux2_1
X_14025_ hold1911/X _14038_/B _14024_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _14025_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11168_ _16880_/Q _11744_/B _11168_/C vssd1 vssd1 vccd1 vccd1 _11168_/X sky130_fd_sc_hd__and3_1
XTAP_6260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10119_ _10563_/A _10119_/B vssd1 vssd1 vccd1 vccd1 _10119_/X sky130_fd_sc_hd__or2_1
XTAP_5570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15976_ _17295_/CLK _15976_/D vssd1 vssd1 vccd1 vccd1 hold799/A sky130_fd_sc_hd__dfxtp_1
X_11099_ hold1616/X _16857_/Q _11210_/C vssd1 vssd1 vccd1 vccd1 _11100_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_234_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17715_ _17747_/CLK _17715_/D vssd1 vssd1 vccd1 vccd1 _17715_/Q sky130_fd_sc_hd__dfxtp_1
X_14927_ hold6054/X _14946_/B _14926_/X _15048_/A vssd1 vssd1 vccd1 vccd1 _14927_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_426_wb_clk_i clkbuf_6_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17590_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17646_ _17678_/CLK _17646_/D vssd1 vssd1 vccd1 vccd1 _17646_/Q sky130_fd_sc_hd__dfxtp_1
X_14858_ _15197_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14858_/X sky130_fd_sc_hd__or2_1
XFILLER_0_216_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13809_ hold5723/X _13719_/A _13808_/X vssd1 vssd1 vccd1 vccd1 _13809_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_212_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17577_ _17737_/CLK _17577_/D vssd1 vssd1 vccd1 vccd1 _17577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14789_ _14789_/A _14843_/B vssd1 vssd1 vccd1 vccd1 _14830_/B sky130_fd_sc_hd__or2_4
XFILLER_0_86_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16528_ _18106_/CLK _16528_/D vssd1 vssd1 vccd1 vccd1 _16528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16459_ _17535_/CLK _16459_/D vssd1 vssd1 vccd1 vccd1 _16459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09000_ hold226/X hold264/X _09056_/S vssd1 vssd1 vccd1 vccd1 hold265/A sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18129_ _18129_/CLK _18129_/D vssd1 vssd1 vccd1 vccd1 _18129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5705 _17113_/Q vssd1 vssd1 vccd1 vccd1 hold5705/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5716 _12352_/Y vssd1 vssd1 vccd1 vccd1 _17274_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5727 _13815_/Y vssd1 vssd1 vccd1 vccd1 _13816_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5738 _12265_/X vssd1 vssd1 vccd1 vccd1 _17245_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5749 _17172_/Q vssd1 vssd1 vccd1 vccd1 hold5749/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09902_ hold2819/X hold4650/X _11162_/C vssd1 vssd1 vccd1 vccd1 _09903_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout504 _11183_/C vssd1 vssd1 vccd1 vccd1 _11216_/C sky130_fd_sc_hd__buf_6
XFILLER_0_111_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout515 _09499_/Y vssd1 vssd1 vccd1 vccd1 _10385_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout526 _09285_/Y vssd1 vssd1 vccd1 vccd1 _09323_/B sky130_fd_sc_hd__buf_4
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09833_ hold1833/X _16435_/Q _10031_/C vssd1 vssd1 vccd1 vccd1 _09834_/B sky130_fd_sc_hd__mux2_1
Xfanout537 _09066_/Y vssd1 vssd1 vccd1 vccd1 _09102_/B sky130_fd_sc_hd__buf_4
Xfanout548 hold114/X vssd1 vssd1 vccd1 vccd1 hold115/A sky130_fd_sc_hd__buf_6
XFILLER_0_67_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout559 hold107/X vssd1 vssd1 vccd1 vccd1 hold108/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_226_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09764_ hold3171/X hold3562/X _10040_/C vssd1 vssd1 vccd1 vccd1 _09765_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08715_ hold438/X hold812/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08716_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_167_wb_clk_i clkbuf_6_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18271_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_174_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09695_ hold2596/X hold3572/X _10025_/C vssd1 vssd1 vccd1 vccd1 _09696_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08646_ _12416_/A hold488/X vssd1 vssd1 vccd1 vccd1 _15945_/D sky130_fd_sc_hd__and2_1
XFILLER_0_83_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08577_ _15274_/A _08577_/B vssd1 vssd1 vccd1 vccd1 _15912_/D sky130_fd_sc_hd__and2_1
XFILLER_0_7_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10470_ _10470_/A _10470_/B vssd1 vssd1 vccd1 vccd1 _10470_/X sky130_fd_sc_hd__or2_1
XFILLER_0_91_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09129_ hold1246/X _09177_/A2 _09128_/X _12855_/A vssd1 vssd1 vccd1 vccd1 _09129_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12140_ hold1574/X _17204_/Q _12332_/C vssd1 vssd1 vccd1 vccd1 _12141_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12071_ hold2310/X _17181_/Q _12332_/C vssd1 vssd1 vccd1 vccd1 _12072_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold580 hold580/A vssd1 vssd1 vccd1 vccd1 hold580/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold591 hold591/A vssd1 vssd1 vccd1 vccd1 hold591/X sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ _11088_/A _11022_/B vssd1 vssd1 vccd1 vccd1 _11022_/X sky130_fd_sc_hd__or2_1
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15830_ _17721_/CLK _15830_/D vssd1 vssd1 vccd1 vccd1 _15830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _17739_/CLK _15761_/D vssd1 vssd1 vccd1 vccd1 _15761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12973_ hold2830/X hold3787/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12973_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_232_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _17500_/CLK _17500_/D vssd1 vssd1 vccd1 vccd1 _17500_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1280 _08097_/X vssd1 vssd1 vccd1 vccd1 _15688_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14712_ _15213_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14712_/X sky130_fd_sc_hd__or2_1
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1291 _15747_/Q vssd1 vssd1 vccd1 vccd1 hold1291/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ hold1293/X _17132_/Q _13721_/S vssd1 vssd1 vccd1 vccd1 _11925_/B sky130_fd_sc_hd__mux2_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _17260_/CLK _15692_/D vssd1 vssd1 vccd1 vccd1 _15692_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _17754_/CLK _17431_/D vssd1 vssd1 vccd1 vccd1 _17431_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ hold1041/X _14664_/B _14642_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _14643_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ hold2902/X hold4433/X _12335_/C vssd1 vssd1 vccd1 vccd1 _11856_/B sky130_fd_sc_hd__mux2_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10806_ _11121_/A _10806_/B vssd1 vssd1 vccd1 vccd1 _10806_/X sky130_fd_sc_hd__or2_1
X_17362_ _17516_/CLK _17362_/D vssd1 vssd1 vccd1 vccd1 _17362_/Q sky130_fd_sc_hd__dfxtp_1
X_14574_ hold927/X _14622_/B vssd1 vssd1 vccd1 vccd1 _14574_/X sky130_fd_sc_hd__or2_1
X_11786_ _17086_/Q _11786_/B _12329_/C vssd1 vssd1 vccd1 vccd1 _11786_/X sky130_fd_sc_hd__and3_1
XFILLER_0_83_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16313_ _16323_/CLK _16313_/D vssd1 vssd1 vccd1 vccd1 _16313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13525_ hold4709/X _13811_/B _13524_/X _08363_/A vssd1 vssd1 vccd1 vccd1 _13525_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17293_ _17293_/CLK _17293_/D vssd1 vssd1 vccd1 vccd1 hold810/A sky130_fd_sc_hd__dfxtp_1
X_10737_ _11121_/A _10737_/B vssd1 vssd1 vccd1 vccd1 _10737_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16244_ _17425_/CLK _16244_/D vssd1 vssd1 vccd1 vccd1 hold572/A sky130_fd_sc_hd__dfxtp_1
X_13456_ hold5231/X _13856_/B _13455_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13456_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10668_ _11049_/A _10668_/B vssd1 vssd1 vccd1 vccd1 _10668_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12407_ hold169/X _17297_/Q _12443_/S vssd1 vssd1 vccd1 vccd1 hold170/A sky130_fd_sc_hd__mux2_1
XFILLER_0_144_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16175_ _17750_/CLK _16175_/D vssd1 vssd1 vccd1 vccd1 _16175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10599_ hold4340/X _10563_/A _10598_/X vssd1 vssd1 vccd1 vccd1 _10600_/B sky130_fd_sc_hd__a21oi_1
X_13387_ hold5249/X _12356_/B _13386_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _13387_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput107 hold4201/X vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_12
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15126_ hold1648/X hold340/X _15125_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _15126_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput118 hold5916/X vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_12
Xoutput129 hold5920/X vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_12
XFILLER_0_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12338_ _12338_/A _12350_/B _13463_/S vssd1 vssd1 vccd1 vccd1 _12338_/X sky130_fd_sc_hd__and3_1
XFILLER_0_105_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15057_ hold220/X hold788/X _15071_/S vssd1 vssd1 vccd1 vccd1 hold789/A sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12269_ hold2439/X _17247_/Q _12371_/C vssd1 vssd1 vccd1 vccd1 _12270_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2909 _14301_/X vssd1 vssd1 vccd1 vccd1 _17950_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14008_ _14850_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14008_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_260_wb_clk_i clkbuf_6_58_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18066_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15959_ _17338_/CLK _15959_/D vssd1 vssd1 vccd1 vccd1 hold732/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08500_ _14732_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08500_/X sky130_fd_sc_hd__or2_1
X_09480_ _09483_/B _09483_/C vssd1 vssd1 vccd1 vccd1 _09482_/B sky130_fd_sc_hd__and2_1
XFILLER_0_210_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08431_ _15219_/A _08433_/B vssd1 vssd1 vccd1 vccd1 _08431_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17629_ _17661_/CLK _17629_/D vssd1 vssd1 vccd1 vccd1 _17629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08362_ _15531_/A hold1172/X hold115/X vssd1 vssd1 vccd1 vccd1 _08363_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08293_ _14457_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08293_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5502 _17606_/Q vssd1 vssd1 vccd1 vccd1 hold5502/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5513 _17643_/Q vssd1 vssd1 vccd1 vccd1 hold5513/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5524 _10978_/X vssd1 vssd1 vccd1 vccd1 _16816_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5535 _16792_/Q vssd1 vssd1 vccd1 vccd1 hold5535/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4801 _16400_/Q vssd1 vssd1 vccd1 vccd1 hold4801/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5546 _13789_/X vssd1 vssd1 vccd1 vccd1 _17716_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5557 _17673_/Q vssd1 vssd1 vccd1 vccd1 hold5557/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4812 _12112_/X vssd1 vssd1 vccd1 vccd1 _17194_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4823 _17697_/Q vssd1 vssd1 vccd1 vccd1 hold4823/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5568 _11620_/X vssd1 vssd1 vccd1 vccd1 _17030_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4834 _09604_/X vssd1 vssd1 vccd1 vccd1 _16358_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5579 _17702_/Q vssd1 vssd1 vccd1 vccd1 hold5579/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4845 _16814_/Q vssd1 vssd1 vccd1 vccd1 hold4845/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4856 _12226_/X vssd1 vssd1 vccd1 vccd1 _17232_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4867 _17635_/Q vssd1 vssd1 vccd1 vccd1 hold4867/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout301 _11061_/A vssd1 vssd1 vccd1 vccd1 _11049_/A sky130_fd_sc_hd__buf_4
Xfanout312 _10986_/A vssd1 vssd1 vccd1 vccd1 _11109_/A sky130_fd_sc_hd__buf_4
Xhold4878 _11263_/X vssd1 vssd1 vccd1 vccd1 _16911_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout323 wire337/X vssd1 vssd1 vccd1 vccd1 _10539_/A sky130_fd_sc_hd__clkbuf_4
Xhold4889 _16875_/Q vssd1 vssd1 vccd1 vccd1 hold4889/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout334 _10542_/A vssd1 vssd1 vccd1 vccd1 _10536_/A sky130_fd_sc_hd__buf_4
XFILLER_0_22_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_348_wb_clk_i clkbuf_6_42_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17639_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout345 _09368_/Y vssd1 vssd1 vccd1 vccd1 _15489_/A sky130_fd_sc_hd__clkbuf_8
Xfanout356 _08657_/S vssd1 vssd1 vccd1 vccd1 _08661_/S sky130_fd_sc_hd__buf_8
XFILLER_0_226_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09816_ _09948_/A _09816_/B vssd1 vssd1 vccd1 vccd1 _09816_/X sky130_fd_sc_hd__or2_1
Xfanout367 _15127_/Y vssd1 vssd1 vccd1 vccd1 _15167_/B sky130_fd_sc_hd__buf_8
Xfanout378 _14912_/Y vssd1 vssd1 vccd1 vccd1 _14952_/B sky130_fd_sc_hd__buf_8
Xfanout389 _14730_/B vssd1 vssd1 vccd1 vccd1 _14732_/B sky130_fd_sc_hd__buf_6
XFILLER_0_241_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09747_ _09957_/A _09747_/B vssd1 vssd1 vccd1 vccd1 _09747_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09678_ _10482_/A _09678_/B vssd1 vssd1 vccd1 vccd1 _09678_/X sky130_fd_sc_hd__or2_1
XFILLER_0_213_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08629_ hold180/X hold525/X _08657_/S vssd1 vssd1 vccd1 vccd1 hold526/A sky130_fd_sc_hd__mux2_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11640_ _11649_/A _11640_/B vssd1 vssd1 vccd1 vccd1 _11640_/X sky130_fd_sc_hd__or2_1
XFILLER_0_194_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11571_ _11661_/A _11571_/B vssd1 vssd1 vccd1 vccd1 _11571_/X sky130_fd_sc_hd__or2_1
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13310_ _13310_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13310_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_64_wb_clk_i clkbuf_6_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17750_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10522_ hold5424/X _11213_/B _10521_/X _14342_/A vssd1 vssd1 vccd1 vccd1 _10522_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14290_ _14970_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14290_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13241_ _13241_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13241_/X sky130_fd_sc_hd__and2_1
X_10453_ hold4626/X _10646_/B _10452_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10453_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10384_ hold4009/X _11186_/B _10383_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10384_/X
+ sky130_fd_sc_hd__o211a_1
X_13172_ hold3483/X _13171_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13172_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12123_ _12219_/A _12123_/B vssd1 vssd1 vccd1 vccd1 _12123_/X sky130_fd_sc_hd__or2_1
XFILLER_0_241_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17980_ _18042_/CLK _17980_/D vssd1 vssd1 vccd1 vccd1 _17980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12054_ _12273_/A _12054_/B vssd1 vssd1 vccd1 vccd1 _12054_/X sky130_fd_sc_hd__or2_1
X_16931_ _17779_/CLK _16931_/D vssd1 vssd1 vccd1 vccd1 _16931_/Q sky130_fd_sc_hd__dfxtp_1
X_11005_ hold5209/X _11195_/B _11004_/X _14462_/C1 vssd1 vssd1 vccd1 vccd1 _11005_/X
+ sky130_fd_sc_hd__o211a_1
X_16862_ _18065_/CLK _16862_/D vssd1 vssd1 vccd1 vccd1 _16862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15813_ _17628_/CLK _15813_/D vssd1 vssd1 vccd1 vccd1 _15813_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout890 _15085_/A vssd1 vssd1 vccd1 vccd1 _15193_/A sky130_fd_sc_hd__buf_8
XFILLER_0_232_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16793_ _18028_/CLK _16793_/D vssd1 vssd1 vccd1 vccd1 _16793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15744_ _17747_/CLK _15744_/D vssd1 vssd1 vccd1 vccd1 _15744_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12956_ hold4151/X _12955_/X _12986_/S vssd1 vssd1 vccd1 vccd1 _12957_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _18463_/A vssd1 vssd1 vccd1 vccd1 _18463_/X sky130_fd_sc_hd__buf_1
XFILLER_0_213_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11907_ _13797_/A _11907_/B vssd1 vssd1 vccd1 vccd1 _11907_/X sky130_fd_sc_hd__or2_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15675_ _17771_/CLK _15675_/D vssd1 vssd1 vccd1 vccd1 _15675_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12887_ hold3352/X _12886_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12888_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_158_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17414_ _17430_/CLK _17414_/D vssd1 vssd1 vccd1 vccd1 _17414_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14626_ _14627_/A _15182_/B vssd1 vssd1 vccd1 vccd1 _14626_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_28_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18394_ _18394_/CLK hold486/X vssd1 vssd1 vccd1 vccd1 _18394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11838_ _12219_/A _11838_/B vssd1 vssd1 vccd1 vccd1 _11838_/X sky130_fd_sc_hd__or2_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _17345_/CLK hold57/X vssd1 vssd1 vccd1 vccd1 _17345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _15492_/A _14573_/B vssd1 vssd1 vccd1 vccd1 _14557_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_126_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11769_ hold4353/X _11694_/A _11768_/X vssd1 vssd1 vccd1 vccd1 _11769_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13508_ hold2615/X hold4785/X _13817_/C vssd1 vssd1 vccd1 vccd1 _13509_/B sky130_fd_sc_hd__mux2_1
X_17276_ _17614_/CLK _17276_/D vssd1 vssd1 vccd1 vccd1 _17276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14488_ hold2573/X _14487_/B _14487_/Y _14356_/A vssd1 vssd1 vccd1 vccd1 _14488_/X
+ sky130_fd_sc_hd__o211a_1
X_16227_ _18458_/CLK _16227_/D vssd1 vssd1 vccd1 vccd1 _16227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13439_ hold2741/X hold4630/X _13862_/C vssd1 vssd1 vccd1 vccd1 _13440_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_141_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16158_ _17513_/CLK _16158_/D vssd1 vssd1 vccd1 vccd1 _16158_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4108 _12530_/X vssd1 vssd1 vccd1 vccd1 _12531_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4119 _17030_/Q vssd1 vssd1 vccd1 vccd1 hold4119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15109_ _15543_/A hold340/X vssd1 vssd1 vccd1 vccd1 _15109_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_228_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3407 _10605_/Y vssd1 vssd1 vccd1 vccd1 _10606_/B sky130_fd_sc_hd__dlygate4sd3_1
X_16089_ _18417_/CLK _16089_/D vssd1 vssd1 vccd1 vccd1 hold754/A sky130_fd_sc_hd__dfxtp_1
X_08980_ _15314_/A _08980_/B vssd1 vssd1 vccd1 vccd1 _16107_/D sky130_fd_sc_hd__and2_1
XFILLER_0_227_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3418 _16349_/Q vssd1 vssd1 vccd1 vccd1 _13262_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3429 _10569_/Y vssd1 vssd1 vccd1 vccd1 _10570_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_441_wb_clk_i clkbuf_6_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17720_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07931_ hold3027/X _07924_/B _07930_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _07931_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2706 _08059_/X vssd1 vssd1 vccd1 vccd1 _15669_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2717 _08469_/X vssd1 vssd1 vccd1 vccd1 _15863_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2728 _14851_/X vssd1 vssd1 vccd1 vccd1 _18214_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2739 _18112_/Q vssd1 vssd1 vccd1 vccd1 hold2739/X sky130_fd_sc_hd__dlygate4sd3_1
X_07862_ hold1865/X _07865_/B _07861_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _07862_/X
+ sky130_fd_sc_hd__o211a_1
X_09601_ hold3572/X _10025_/B _09600_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09601_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07793_ hold5978/X _07788_/A hold1119/X _14556_/A vssd1 vssd1 vccd1 vccd1 _07794_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_09532_ hold5825/X _10022_/B _09531_/X _15202_/C1 vssd1 vssd1 vccd1 vccd1 _09532_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09463_ _09463_/A _09463_/B _09463_/C _09463_/D vssd1 vssd1 vccd1 vccd1 _09472_/D
+ sky130_fd_sc_hd__and4_1
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08414_ hold2741/X _08442_/A2 _08413_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _08414_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09394_ hold5963/A _15490_/B1 _09393_/X _15481_/A1 vssd1 vssd1 vccd1 vccd1 _09394_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_231_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08345_ _08347_/A _08345_/B vssd1 vssd1 vccd1 vccd1 _15804_/D sky130_fd_sc_hd__and2_1
XFILLER_0_191_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08276_ _15555_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08276_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6000 _16531_/Q vssd1 vssd1 vccd1 vccd1 hold6000/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6011 _17540_/Q vssd1 vssd1 vccd1 vccd1 hold6011/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6022 _17753_/Q vssd1 vssd1 vccd1 vccd1 hold6022/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6033 _17528_/Q vssd1 vssd1 vccd1 vccd1 hold6033/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6044 data_in[23] vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6055 _17888_/Q vssd1 vssd1 vccd1 vccd1 hold6055/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5310 _11503_/X vssd1 vssd1 vccd1 vccd1 _16991_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5321 _17044_/Q vssd1 vssd1 vccd1 vccd1 hold5321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6066 _18268_/Q vssd1 vssd1 vccd1 vccd1 hold6066/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6077 _18388_/Q vssd1 vssd1 vccd1 vccd1 hold6077/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5332 _11896_/X vssd1 vssd1 vccd1 vccd1 _17122_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold6088 data_in[20] vssd1 vssd1 vccd1 vccd1 hold120/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5343 _16825_/Q vssd1 vssd1 vccd1 vccd1 hold5343/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6099 _18423_/Q vssd1 vssd1 vccd1 vccd1 hold6099/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5354 _10834_/X vssd1 vssd1 vccd1 vccd1 _16768_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4620 _16641_/Q vssd1 vssd1 vccd1 vccd1 hold4620/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5365 _10846_/X vssd1 vssd1 vccd1 vccd1 _16772_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4631 _13345_/X vssd1 vssd1 vccd1 vccd1 _17568_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5376 _17004_/Q vssd1 vssd1 vccd1 vccd1 hold5376/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4642 _17633_/Q vssd1 vssd1 vccd1 vccd1 hold4642/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5387 _13666_/X vssd1 vssd1 vccd1 vccd1 _17675_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4653 _09904_/X vssd1 vssd1 vccd1 vccd1 _16458_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5398 _16802_/Q vssd1 vssd1 vccd1 vccd1 hold5398/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4664 _17602_/Q vssd1 vssd1 vccd1 vccd1 hold4664/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3930 hold6132/X vssd1 vssd1 vccd1 vccd1 hold3930/X sky130_fd_sc_hd__clkbuf_2
Xhold4675 _11721_/Y vssd1 vssd1 vccd1 vccd1 _11722_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3941 _10492_/X vssd1 vssd1 vccd1 vccd1 _16654_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_182_wb_clk_i clkbuf_6_51_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18393_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4686 _13534_/X vssd1 vssd1 vccd1 vccd1 _17631_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3952 _17688_/Q vssd1 vssd1 vccd1 vccd1 hold3952/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4697 _17596_/Q vssd1 vssd1 vccd1 vccd1 hold4697/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3963 _13723_/X vssd1 vssd1 vccd1 vccd1 _17694_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_111_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17344_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold3974 _16661_/Q vssd1 vssd1 vccd1 vccd1 hold3974/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout153 _12905_/S vssd1 vssd1 vccd1 vccd1 _12920_/S sky130_fd_sc_hd__buf_6
Xhold3985 _16777_/Q vssd1 vssd1 vccd1 vccd1 hold3985/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3996 _10201_/X vssd1 vssd1 vccd1 vccd1 _16557_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout164 _13817_/B vssd1 vssd1 vccd1 vccd1 _12308_/B sky130_fd_sc_hd__clkbuf_8
Xfanout175 _11723_/B vssd1 vssd1 vccd1 vccd1 _11726_/B sky130_fd_sc_hd__clkbuf_8
Xfanout186 _13868_/B vssd1 vssd1 vccd1 vccd1 _13847_/B sky130_fd_sc_hd__clkbuf_8
Xfanout197 fanout210/X vssd1 vssd1 vccd1 vccd1 _12365_/B sky130_fd_sc_hd__buf_4
XFILLER_0_226_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12810_ _12810_/A _12810_/B vssd1 vssd1 vccd1 vccd1 _17446_/D sky130_fd_sc_hd__and2_1
XFILLER_0_69_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13790_ hold2671/X _17717_/Q _13880_/C vssd1 vssd1 vccd1 vccd1 _13791_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_96_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _12750_/A _12741_/B vssd1 vssd1 vccd1 vccd1 _17423_/D sky130_fd_sc_hd__and2_1
XFILLER_0_201_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _07805_/A _15477_/A2 _09392_/A _16075_/Q vssd1 vssd1 vccd1 vccd1 _15460_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12672_ _12873_/A _12672_/B vssd1 vssd1 vccd1 vccd1 _17400_/D sky130_fd_sc_hd__and2_1
XFILLER_0_166_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14411_ _15199_/A _14443_/B vssd1 vssd1 vccd1 vccd1 _14411_/X sky130_fd_sc_hd__or2_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ hold4177/X _12299_/B _11622_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _11623_/X
+ sky130_fd_sc_hd__o211a_1
X_15391_ _16303_/Q _15477_/A2 _15487_/B1 hold667/X _15390_/X vssd1 vssd1 vccd1 vccd1
+ _15392_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_167_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17130_ _17194_/CLK _17130_/D vssd1 vssd1 vccd1 vccd1 _17130_/Q sky130_fd_sc_hd__dfxtp_1
X_14342_ _14342_/A _14342_/B vssd1 vssd1 vccd1 vccd1 _17970_/D sky130_fd_sc_hd__and2_1
XFILLER_0_37_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11554_ hold4040/X _11741_/B _11553_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11554_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10505_ hold1925/X hold3805/X _10595_/C vssd1 vssd1 vccd1 vccd1 _10506_/B sky130_fd_sc_hd__mux2_1
X_17061_ _18427_/CLK _17061_/D vssd1 vssd1 vccd1 vccd1 _17061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14273_ hold2435/X _14272_/B _14272_/Y _14528_/C1 vssd1 vssd1 vccd1 vccd1 _14273_/X
+ sky130_fd_sc_hd__o211a_1
X_11485_ hold4149/X _11771_/B _11484_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _11485_/X
+ sky130_fd_sc_hd__o211a_1
X_16012_ _18419_/CLK _16012_/D vssd1 vssd1 vccd1 vccd1 _16012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13224_ _13217_/X _13223_/X _13296_/B1 vssd1 vssd1 vccd1 vccd1 _17546_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_21_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10436_ hold2928/X hold4628/X _11213_/C vssd1 vssd1 vccd1 vccd1 _10437_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_221_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13155_ _13154_/X _16912_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13155_/X sky130_fd_sc_hd__mux2_1
X_10367_ hold2867/X _16613_/Q _10601_/C vssd1 vssd1 vccd1 vccd1 _10368_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ hold4797/X _13811_/B _12105_/X _08363_/A vssd1 vssd1 vccd1 vccd1 _12106_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13086_ _13086_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13086_/X sky130_fd_sc_hd__or2_1
X_10298_ hold2021/X _16590_/Q _10604_/C vssd1 vssd1 vccd1 vccd1 _10299_/B sky130_fd_sc_hd__mux2_1
X_17963_ _17997_/CLK _17963_/D vssd1 vssd1 vccd1 vccd1 _17963_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12037_ hold5430/X _12329_/B _12036_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _12037_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16914_ _17859_/CLK _16914_/D vssd1 vssd1 vccd1 vccd1 _16914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17894_ _17894_/CLK _17894_/D vssd1 vssd1 vccd1 vccd1 _17894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16845_ _18048_/CLK _16845_/D vssd1 vssd1 vccd1 vccd1 _16845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_233_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_233_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16776_ _18043_/CLK _16776_/D vssd1 vssd1 vccd1 vccd1 _16776_/Q sky130_fd_sc_hd__dfxtp_1
X_13988_ _14543_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13988_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15727_ _17730_/CLK _15727_/D vssd1 vssd1 vccd1 vccd1 _15727_/Q sky130_fd_sc_hd__dfxtp_1
X_12939_ _12948_/A _12939_/B vssd1 vssd1 vccd1 vccd1 _17489_/D sky130_fd_sc_hd__and2_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_238_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15658_ _17202_/CLK _15658_/D vssd1 vssd1 vccd1 vccd1 _15658_/Q sky130_fd_sc_hd__dfxtp_1
X_18446_ _18447_/CLK _18446_/D vssd1 vssd1 vccd1 vccd1 _18446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14609_ hold2300/X _14612_/B _14608_/Y _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14609_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18377_ _18377_/CLK _18377_/D vssd1 vssd1 vccd1 vccd1 _18377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15589_ _17269_/CLK _15589_/D vssd1 vssd1 vccd1 vccd1 _15589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08130_ _14529_/A hold1411/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08130_/X sky130_fd_sc_hd__mux2_1
X_17328_ _17328_/CLK hold78/X vssd1 vssd1 vccd1 vccd1 _17328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08061_ hold1277/X _08097_/A2 _08060_/X _12103_/C1 vssd1 vssd1 vccd1 vccd1 _08061_/X
+ sky130_fd_sc_hd__o211a_1
X_17259_ _17259_/CLK _17259_/D vssd1 vssd1 vccd1 vccd1 _17259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3204 _16345_/Q vssd1 vssd1 vccd1 vccd1 _13230_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3215 _09919_/X vssd1 vssd1 vccd1 vccd1 _16463_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3226 _17429_/Q vssd1 vssd1 vccd1 vccd1 hold3226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3237 _16379_/Q vssd1 vssd1 vccd1 vccd1 hold3237/X sky130_fd_sc_hd__dlygate4sd3_1
X_08963_ hold172/X hold688/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08964_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3248 _10099_/X vssd1 vssd1 vccd1 vccd1 _16523_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2503 _15687_/Q vssd1 vssd1 vccd1 vccd1 hold2503/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3259 _16615_/Q vssd1 vssd1 vccd1 vccd1 hold3259/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2514 _17917_/Q vssd1 vssd1 vccd1 vccd1 hold2514/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2525 _15694_/Q vssd1 vssd1 vccd1 vccd1 hold2525/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2536 _18318_/Q vssd1 vssd1 vccd1 vccd1 hold2536/X sky130_fd_sc_hd__dlygate4sd3_1
X_07914_ _15537_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07914_/X sky130_fd_sc_hd__or2_1
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1802 _14887_/X vssd1 vssd1 vccd1 vccd1 _18232_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2547 _14548_/X vssd1 vssd1 vccd1 vccd1 _18070_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08894_ hold77/X hold531/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08895_/B sky130_fd_sc_hd__mux2_1
Xhold1813 _18426_/Q vssd1 vssd1 vccd1 vccd1 hold1813/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2558 _09219_/X vssd1 vssd1 vccd1 vccd1 _16221_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2569 _18367_/Q vssd1 vssd1 vccd1 vccd1 hold2569/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1824 _09211_/X vssd1 vssd1 vccd1 vccd1 _16217_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1835 _18244_/Q vssd1 vssd1 vccd1 vccd1 hold1835/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1846 _14819_/X vssd1 vssd1 vccd1 vccd1 _18199_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07845_ _14517_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07845_/X sky130_fd_sc_hd__or2_1
Xhold1857 _18380_/Q vssd1 vssd1 vccd1 vccd1 hold1857/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1868 _14490_/X vssd1 vssd1 vccd1 vccd1 _18042_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1879 _16322_/Q vssd1 vssd1 vccd1 vccd1 _09483_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_224_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09515_ hold2390/X _13102_/A _10004_/C vssd1 vssd1 vccd1 vccd1 _09516_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _09444_/X _09446_/B _09478_/B vssd1 vssd1 vccd1 vccd1 _16308_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_91_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09377_ hold5931/A _09342_/B _09342_/Y _09376_/X _15314_/A vssd1 vssd1 vccd1 vccd1
+ _09377_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08328_ hold1332/X _08336_/A2 _08327_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _08328_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08259_ hold1538/X _08262_/B _08258_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _08259_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_363_wb_clk_i clkbuf_6_35_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17743_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11270_ hold971/X hold4312/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11271_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5140 _16978_/Q vssd1 vssd1 vccd1 vccd1 hold5140/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10221_ _10413_/A _10221_/B vssd1 vssd1 vccd1 vccd1 _10221_/X sky130_fd_sc_hd__or2_1
Xhold5151 _13489_/X vssd1 vssd1 vccd1 vccd1 _17616_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5162 _11584_/X vssd1 vssd1 vccd1 vccd1 _17018_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5173 _16883_/Q vssd1 vssd1 vccd1 vccd1 hold5173/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5184 _11383_/X vssd1 vssd1 vccd1 vccd1 _16951_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4450 _11787_/Y vssd1 vssd1 vccd1 vccd1 _11788_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5195 _17042_/Q vssd1 vssd1 vccd1 vccd1 hold5195/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10152_ _10536_/A _10152_/B vssd1 vssd1 vccd1 vccd1 _10152_/X sky130_fd_sc_hd__or2_1
Xhold4461 _16572_/Q vssd1 vssd1 vccd1 vccd1 hold4461/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4472 _12306_/Y vssd1 vssd1 vccd1 vccd1 _12307_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4483 _10360_/X vssd1 vssd1 vccd1 vccd1 _16610_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4494 _10252_/X vssd1 vssd1 vccd1 vccd1 _16574_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3760 _12953_/X vssd1 vssd1 vccd1 vccd1 _12954_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10083_ _10563_/A _10083_/B vssd1 vssd1 vccd1 vccd1 _10083_/X sky130_fd_sc_hd__or2_1
X_14960_ _14960_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14960_/X sky130_fd_sc_hd__or2_1
Xhold3771 _16840_/Q vssd1 vssd1 vccd1 vccd1 hold3771/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3782 _10315_/X vssd1 vssd1 vccd1 vccd1 _16595_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3793 _17410_/Q vssd1 vssd1 vccd1 vccd1 hold3793/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13911_ _13911_/A _13911_/B vssd1 vssd1 vccd1 vccd1 _17763_/D sky130_fd_sc_hd__and2_1
XTAP_5977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14891_ hold2869/X hold332/X _14890_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _14891_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16630_ _18154_/CLK _16630_/D vssd1 vssd1 vccd1 vccd1 _16630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13842_ hold4498/X _13752_/A _13841_/X vssd1 vssd1 vccd1 vccd1 _13842_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_215_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16561_ _18099_/CLK _16561_/D vssd1 vssd1 vccd1 vccd1 _16561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13773_ _13773_/A _13773_/B vssd1 vssd1 vccd1 vccd1 _13773_/X sky130_fd_sc_hd__or2_1
X_10985_ hold2171/X _16819_/Q _10985_/S vssd1 vssd1 vccd1 vccd1 _10986_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18300_ _18390_/CLK _18300_/D vssd1 vssd1 vccd1 vccd1 _18300_/Q sky130_fd_sc_hd__dfxtp_1
X_15512_ hold1155/X _15560_/A2 _15511_/X _12864_/A vssd1 vssd1 vccd1 vccd1 _15512_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12724_ hold1069/X _17419_/Q _12766_/S vssd1 vssd1 vccd1 vccd1 _12724_/X sky130_fd_sc_hd__mux2_1
X_16492_ _18242_/CLK _16492_/D vssd1 vssd1 vccd1 vccd1 _16492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18231_ _18231_/CLK hold333/X vssd1 vssd1 vccd1 vccd1 _18231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15443_ _15481_/A1 _15435_/X _15442_/X _15481_/B1 hold5965/A vssd1 vssd1 vccd1 vccd1
+ _15443_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_195_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12655_ hold2179/X _17396_/Q _12850_/S vssd1 vssd1 vccd1 vccd1 _12655_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18162_ _18162_/CLK _18162_/D vssd1 vssd1 vccd1 vccd1 _18162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11606_ hold1718/X _17026_/Q _11774_/C vssd1 vssd1 vccd1 vccd1 _11607_/B sky130_fd_sc_hd__mux2_1
X_15374_ _15374_/A _15374_/B vssd1 vssd1 vccd1 vccd1 _18413_/D sky130_fd_sc_hd__and2_1
XFILLER_0_183_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12586_ hold2944/X _17373_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _12586_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17113_ _17608_/CLK _17113_/D vssd1 vssd1 vccd1 vccd1 _17113_/Q sky130_fd_sc_hd__dfxtp_1
X_14325_ hold2429/X _14326_/B _14324_/Y _14390_/A vssd1 vssd1 vccd1 vccd1 _14325_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18093_ _18125_/CLK _18093_/D vssd1 vssd1 vccd1 vccd1 _18093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11537_ hold2520/X _17003_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _11538_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_184_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold409 hold409/A vssd1 vssd1 vccd1 vccd1 hold409/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17044_ _17892_/CLK _17044_/D vssd1 vssd1 vccd1 vccd1 _17044_/Q sky130_fd_sc_hd__dfxtp_1
X_14256_ _14596_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14256_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11468_ hold1660/X _16980_/Q _11660_/S vssd1 vssd1 vccd1 vccd1 _11469_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13207_ _13311_/A1 _13205_/X _13206_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13207_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10419_ _10515_/A _10419_/B vssd1 vssd1 vccd1 vccd1 _10419_/X sky130_fd_sc_hd__or2_1
X_14187_ hold1534/X _14202_/B _14186_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14187_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_1326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11399_ hold2023/X hold5561/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11400_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _17568_/Q _17102_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13138_/X sky130_fd_sc_hd__mux2_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13069_ _13068_/X hold3930/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13069_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17946_ _18010_/CLK _17946_/D vssd1 vssd1 vccd1 vccd1 _17946_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1109 _15150_/X vssd1 vssd1 vccd1 vccd1 _18358_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17877_ _17877_/CLK _17877_/D vssd1 vssd1 vccd1 vccd1 _17877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16828_ _18031_/CLK _16828_/D vssd1 vssd1 vccd1 vccd1 _16828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_215_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16759_ _18024_/CLK _16759_/D vssd1 vssd1 vccd1 vccd1 _16759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09300_ hold2834/X _09325_/B _09299_/X _12984_/A vssd1 vssd1 vccd1 vccd1 _09300_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_232_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09231_ hold1614/X _09218_/B _09230_/X _12843_/A vssd1 vssd1 vccd1 vccd1 _09231_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18429_ _18429_/CLK _18429_/D vssd1 vssd1 vccd1 vccd1 _18429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09162_ _15545_/A _09164_/B vssd1 vssd1 vccd1 vccd1 _09162_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_111_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08113_ _13927_/A _08113_/B vssd1 vssd1 vccd1 vccd1 _15695_/D sky130_fd_sc_hd__and2_1
XFILLER_0_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09093_ hold2719/X _09102_/B _09092_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _09093_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08044_ hold1358/X _08033_/B _08043_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _08044_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold910 hold910/A vssd1 vssd1 vccd1 vccd1 hold910/X sky130_fd_sc_hd__buf_6
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold921 hold921/A vssd1 vssd1 vccd1 vccd1 hold921/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold932 hold932/A vssd1 vssd1 vccd1 vccd1 hold932/X sky130_fd_sc_hd__buf_6
XFILLER_0_226_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold943 hold974/X vssd1 vssd1 vccd1 vccd1 hold975/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 hold954/A vssd1 vssd1 vccd1 vccd1 hold954/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold965 la_data_in[9] vssd1 vssd1 vccd1 vccd1 hold965/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3001 _09187_/X vssd1 vssd1 vccd1 vccd1 _16205_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 input63/X vssd1 vssd1 vccd1 vccd1 hold976/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold987 hold987/A vssd1 vssd1 vccd1 vccd1 hold987/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3012 _17849_/Q vssd1 vssd1 vccd1 vccd1 hold3012/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 hold998/A vssd1 vssd1 vccd1 vccd1 hold998/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3023 _18019_/Q vssd1 vssd1 vccd1 vccd1 hold3023/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3034 _14587_/X vssd1 vssd1 vccd1 vccd1 _18087_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ _09995_/A _10004_/B _10004_/C vssd1 vssd1 vccd1 vccd1 _09995_/X sky130_fd_sc_hd__and3_1
XTAP_5207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2300 _18098_/Q vssd1 vssd1 vccd1 vccd1 hold2300/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3045 _18162_/Q vssd1 vssd1 vccd1 vccd1 hold3045/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3056 _09304_/X vssd1 vssd1 vccd1 vccd1 _16262_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2311 _07949_/X vssd1 vssd1 vccd1 vccd1 _15617_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2322 _15728_/Q vssd1 vssd1 vccd1 vccd1 hold2322/X sky130_fd_sc_hd__dlygate4sd3_1
X_08946_ _12410_/A _08946_/B vssd1 vssd1 vccd1 vccd1 _16090_/D sky130_fd_sc_hd__and2_1
Xhold3067 _17978_/Q vssd1 vssd1 vccd1 vccd1 hold3067/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2333 _15883_/Q vssd1 vssd1 vccd1 vccd1 hold2333/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3078 _15758_/Q vssd1 vssd1 vccd1 vccd1 hold3078/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2344 _08485_/X vssd1 vssd1 vccd1 vccd1 _15871_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3089 _18441_/Q vssd1 vssd1 vccd1 vccd1 hold3089/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1610 _14973_/X vssd1 vssd1 vccd1 vccd1 _18272_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2355 _15886_/Q vssd1 vssd1 vccd1 vccd1 hold2355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1621 _18310_/Q vssd1 vssd1 vccd1 vccd1 hold1621/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2366 _07840_/X vssd1 vssd1 vccd1 vccd1 _15565_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1632 _15804_/Q vssd1 vssd1 vccd1 vccd1 hold1632/X sky130_fd_sc_hd__dlygate4sd3_1
X_08877_ _15274_/A hold875/X vssd1 vssd1 vccd1 vccd1 _16056_/D sky130_fd_sc_hd__and2_1
Xhold2377 _14825_/X vssd1 vssd1 vccd1 vccd1 _18202_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2388 _15832_/Q vssd1 vssd1 vccd1 vccd1 hold2388/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1643 _18458_/Q vssd1 vssd1 vccd1 vccd1 hold1643/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2399 _08214_/X vssd1 vssd1 vccd1 vccd1 _15743_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1654 _16228_/Q vssd1 vssd1 vccd1 vccd1 hold1654/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1665 _07933_/X vssd1 vssd1 vccd1 vccd1 _15610_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07828_ _14556_/A hold353/A _14555_/C vssd1 vssd1 vccd1 vccd1 hold354/A sky130_fd_sc_hd__or3_1
Xhold1676 _17801_/Q vssd1 vssd1 vccd1 vccd1 hold1676/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1687 _08026_/X vssd1 vssd1 vccd1 vccd1 _15654_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_6_27_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_27_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
Xhold1698 _17886_/Q vssd1 vssd1 vccd1 vccd1 hold1698/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10770_ _11136_/A _10770_/B vssd1 vssd1 vccd1 vccd1 _10770_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09429_ _07785_/Y hold733/X _15274_/A _09428_/X vssd1 vssd1 vccd1 vccd1 hold734/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12440_ _12440_/A hold696/X vssd1 vssd1 vccd1 vccd1 _17313_/D sky130_fd_sc_hd__and2_1
XFILLER_0_192_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12371_ _17281_/Q _12374_/B _12371_/C vssd1 vssd1 vccd1 vccd1 _12371_/X sky130_fd_sc_hd__and3_1
XFILLER_0_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14110_ _14395_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14110_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11322_ _12240_/A _11322_/B vssd1 vssd1 vccd1 vccd1 _11322_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15090_ hold1110/X hold341/X _15089_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _15090_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14041_ hold2324/X _14040_/B _14040_/Y _13933_/A vssd1 vssd1 vccd1 vccd1 _14041_/X
+ sky130_fd_sc_hd__o211a_1
X_11253_ _11637_/A _11253_/B vssd1 vssd1 vccd1 vccd1 _11253_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10204_ hold3558/X _10646_/B _10203_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _10204_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11184_ hold3490/X _11121_/A _11183_/X vssd1 vssd1 vccd1 vccd1 _11184_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4280 _11227_/Y vssd1 vssd1 vccd1 vccd1 _16899_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17800_ _17874_/CLK _17800_/D vssd1 vssd1 vccd1 vccd1 _17800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10135_ hold3328/X _10637_/B _10134_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10135_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4291 _12327_/Y vssd1 vssd1 vccd1 vccd1 _12328_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15992_ _17318_/CLK _15992_/D vssd1 vssd1 vccd1 vccd1 hold544/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3590 _16729_/Q vssd1 vssd1 vccd1 vccd1 hold3590/X sky130_fd_sc_hd__dlygate4sd3_1
X_14943_ hold645/X _14946_/B _14942_/X _15070_/A vssd1 vssd1 vccd1 vccd1 hold646/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10066_ _10603_/A _10066_/B vssd1 vssd1 vccd1 vccd1 _16512_/D sky130_fd_sc_hd__nor2_1
X_17731_ _17731_/CLK _17731_/D vssd1 vssd1 vccd1 vccd1 _17731_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14874_ _15213_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14874_/X sky130_fd_sc_hd__or2_1
X_17662_ _17726_/CLK _17662_/D vssd1 vssd1 vccd1 vccd1 _17662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16613_ _18177_/CLK _16613_/D vssd1 vssd1 vccd1 vccd1 _16613_/Q sky130_fd_sc_hd__dfxtp_1
X_13825_ _13864_/A _13825_/B vssd1 vssd1 vccd1 vccd1 _13825_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_203_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17593_ _17721_/CLK _17593_/D vssd1 vssd1 vccd1 vccd1 _17593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16544_ _18192_/CLK _16544_/D vssd1 vssd1 vccd1 vccd1 _16544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13756_ hold5581/X _13880_/B _13755_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13756_/X
+ sky130_fd_sc_hd__o211a_1
X_10968_ _11067_/A _10968_/B vssd1 vssd1 vccd1 vccd1 _10968_/X sky130_fd_sc_hd__or2_1
XFILLER_0_58_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12707_ hold3722/X _12706_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12707_/X sky130_fd_sc_hd__mux2_1
X_16475_ _18388_/CLK _16475_/D vssd1 vssd1 vccd1 vccd1 _16475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13687_ hold5555/X _13880_/B _13686_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13687_/X
+ sky130_fd_sc_hd__o211a_1
X_10899_ _11091_/A _10899_/B vssd1 vssd1 vccd1 vccd1 _10899_/X sky130_fd_sc_hd__or2_1
XFILLER_0_116_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15426_ _17318_/Q _09357_/A _09392_/A hold532/X vssd1 vssd1 vccd1 vccd1 _15426_/X
+ sky130_fd_sc_hd__a22o_1
X_18214_ _18214_/CLK _18214_/D vssd1 vssd1 vccd1 vccd1 _18214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_285_wb_clk_i clkbuf_6_48_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18321_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12638_ hold3370/X _12637_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12638_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_127_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15357_ hold396/X _15487_/A2 _09386_/D hold815/X _15356_/X vssd1 vssd1 vccd1 vccd1
+ _15362_/B sky130_fd_sc_hd__a221o_1
X_18145_ _18262_/CLK _18145_/D vssd1 vssd1 vccd1 vccd1 _18145_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_214_wb_clk_i clkbuf_6_60_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18205_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12569_ hold4142/X _12568_/X _12986_/S vssd1 vssd1 vccd1 vccd1 _12570_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_124_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5909 _09490_/B vssd1 vssd1 vccd1 vccd1 hold5909/X sky130_fd_sc_hd__dlygate4sd3_1
X_14308_ _14988_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14308_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18076_ _18393_/CLK hold912/X vssd1 vssd1 vccd1 vccd1 _18076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15288_ hold165/X _15484_/A2 _09392_/D _17289_/Q vssd1 vssd1 vccd1 vccd1 _15288_/X
+ sky130_fd_sc_hd__a22o_1
Xhold206 hold206/A vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 la_data_in[18] vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 hold381/X vssd1 vssd1 vccd1 vccd1 hold382/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17027_ _17904_/CLK _17027_/D vssd1 vssd1 vccd1 vccd1 _17027_/Q sky130_fd_sc_hd__dfxtp_1
X_14239_ hold1939/X _14268_/B _14238_/X _14372_/A vssd1 vssd1 vccd1 vccd1 _14239_/X
+ sky130_fd_sc_hd__o211a_1
Xhold239 hold483/X vssd1 vssd1 vccd1 vccd1 hold484/A sky130_fd_sc_hd__buf_6
XFILLER_0_111_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_229_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout708 fanout739/X vssd1 vssd1 vccd1 vccd1 _09047_/A sky130_fd_sc_hd__clkbuf_4
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout719 _09907_/C1 vssd1 vssd1 vccd1 vccd1 _12412_/A sky130_fd_sc_hd__buf_4
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08800_ _12440_/A hold804/X vssd1 vssd1 vccd1 vccd1 _16019_/D sky130_fd_sc_hd__and2_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _09978_/A _09780_/B vssd1 vssd1 vccd1 vccd1 _09780_/X sky130_fd_sc_hd__or2_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ hold226/X hold757/X _08779_/S vssd1 vssd1 vccd1 vccd1 hold758/A sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _17929_/CLK _17929_/D vssd1 vssd1 vccd1 vccd1 _17929_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_234_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08662_ _15274_/A hold862/X vssd1 vssd1 vccd1 vccd1 _15953_/D sky130_fd_sc_hd__and2_1
XFILLER_0_234_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08593_ _15314_/A _08593_/B vssd1 vssd1 vccd1 vccd1 _15920_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09214_ _15543_/A _09214_/B vssd1 vssd1 vccd1 vccd1 _09214_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_162_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09145_ hold1338/X _09177_/A2 _09144_/X _12888_/A vssd1 vssd1 vccd1 vccd1 _09145_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_228_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09076_ _15517_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09076_/X sky130_fd_sc_hd__or2_1
XFILLER_0_115_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08027_ _15541_/A _08029_/B vssd1 vssd1 vccd1 vccd1 _08027_/Y sky130_fd_sc_hd__nand2_1
Xhold740 hold740/A vssd1 vssd1 vccd1 vccd1 hold740/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 hold751/A vssd1 vssd1 vccd1 vccd1 hold751/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 hold762/A vssd1 vssd1 vccd1 vccd1 hold762/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold773 hold773/A vssd1 vssd1 vccd1 vccd1 hold773/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold784 hold784/A vssd1 vssd1 vccd1 vccd1 hold784/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 hold795/A vssd1 vssd1 vccd1 vccd1 hold795/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_1292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_89_wb_clk_i clkbuf_6_17_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17288_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09978_ _09978_/A _09978_/B vssd1 vssd1 vccd1 vccd1 _09978_/X sky130_fd_sc_hd__or2_1
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2130 _14510_/X vssd1 vssd1 vccd1 vccd1 _18051_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2141 _18102_/Q vssd1 vssd1 vccd1 vccd1 hold2141/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_wb_clk_i clkbuf_6_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17462_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08929_ _15324_/A hold568/X vssd1 vssd1 vccd1 vccd1 _16082_/D sky130_fd_sc_hd__and2_1
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2152 _14319_/X vssd1 vssd1 vccd1 vccd1 _17959_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2163 _17912_/Q vssd1 vssd1 vccd1 vccd1 hold2163/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2174 _08036_/X vssd1 vssd1 vccd1 vccd1 _15659_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2185 _18271_/Q vssd1 vssd1 vccd1 vccd1 hold2185/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1440 _17794_/Q vssd1 vssd1 vccd1 vccd1 hold1440/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1451 _15718_/Q vssd1 vssd1 vccd1 vccd1 hold1451/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2196 _14506_/X vssd1 vssd1 vccd1 vccd1 _18049_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ _12234_/A _11940_/B vssd1 vssd1 vccd1 vccd1 _11940_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1462 _14769_/X vssd1 vssd1 vccd1 vccd1 _18175_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1473 _16256_/Q vssd1 vssd1 vccd1 vccd1 hold1473/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1484 _17900_/Q vssd1 vssd1 vccd1 vccd1 hold1484/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1495 _18196_/Q vssd1 vssd1 vccd1 vccd1 hold1495/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _12255_/A _11871_/B vssd1 vssd1 vccd1 vccd1 _11871_/X sky130_fd_sc_hd__or2_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ hold1585/X hold5787/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13611_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10822_ hold4819/X _11204_/B _10821_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _10822_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _15199_/A _14622_/B vssd1 vssd1 vccd1 vccd1 _14590_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13541_ hold613/X _17634_/Q _13829_/C vssd1 vssd1 vccd1 vccd1 _13542_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10753_ hold4995/X _11153_/B _10752_/X _14354_/A vssd1 vssd1 vccd1 vccd1 _10753_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16260_ _17516_/CLK _16260_/D vssd1 vssd1 vccd1 vccd1 _16260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13472_ hold1227/X _17611_/Q _13841_/C vssd1 vssd1 vccd1 vccd1 _13473_/B sky130_fd_sc_hd__mux2_1
X_10684_ hold5243/X _11171_/B _10683_/X _14372_/A vssd1 vssd1 vccd1 vccd1 _10684_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15211_ hold630/A _15233_/B vssd1 vssd1 vccd1 vccd1 hold377/A sky130_fd_sc_hd__or2_1
XFILLER_0_164_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12423_ hold373/X hold410/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12424_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16191_ _17881_/CLK _16191_/D vssd1 vssd1 vccd1 vccd1 _16191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15142_ hold1903/X _15165_/B _15141_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _15142_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12354_ hold4273/X _13314_/A _12353_/X vssd1 vssd1 vccd1 vccd1 _12354_/Y sky130_fd_sc_hd__a21oi_1
X_11305_ hold5561/X _12329_/B _11304_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _11305_/X
+ sky130_fd_sc_hd__o211a_1
X_15073_ hold338/X _15182_/B vssd1 vssd1 vccd1 vccd1 hold339/A sky130_fd_sc_hd__nor2_1
XFILLER_0_26_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12285_ _12285_/A _12285_/B vssd1 vssd1 vccd1 vccd1 _12285_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14024_ _14596_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14024_/X sky130_fd_sc_hd__or2_1
XFILLER_0_142_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11236_ hold5624/X _12305_/B _11235_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11236_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11167_ _12301_/A _11167_/B vssd1 vssd1 vccd1 vccd1 _11167_/Y sky130_fd_sc_hd__nor2_1
XTAP_6261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10118_ hold1012/X _16530_/Q _10634_/C vssd1 vssd1 vccd1 vccd1 _10119_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_235_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15975_ _16086_/CLK _15975_/D vssd1 vssd1 vccd1 vccd1 hold465/A sky130_fd_sc_hd__dfxtp_1
X_11098_ hold5000/X _11195_/B _11097_/X _14526_/C1 vssd1 vssd1 vccd1 vccd1 _11098_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_216_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17714_ _17746_/CLK _17714_/D vssd1 vssd1 vccd1 vccd1 _17714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10049_ _16507_/Q _10049_/B _10049_/C vssd1 vssd1 vccd1 vccd1 _10049_/X sky130_fd_sc_hd__and3_1
X_14926_ _15195_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14926_/X sky130_fd_sc_hd__or2_1
XFILLER_0_175_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_216_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17645_ _17709_/CLK _17645_/D vssd1 vssd1 vccd1 vccd1 _17645_/Q sky130_fd_sc_hd__dfxtp_1
X_14857_ hold1925/X _14880_/B _14856_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14857_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13808_ _17723_/Q _13808_/B _13814_/C vssd1 vssd1 vccd1 vccd1 _13808_/X sky130_fd_sc_hd__and3_1
XFILLER_0_147_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14788_ _14789_/A _14843_/B vssd1 vssd1 vccd1 vccd1 _14788_/Y sky130_fd_sc_hd__nor2_2
X_17576_ _17576_/CLK _17576_/D vssd1 vssd1 vccd1 vccd1 _17576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_212_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16527_ _18213_/CLK _16527_/D vssd1 vssd1 vccd1 vccd1 _16527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13739_ hold1123/X _17700_/Q _13871_/C vssd1 vssd1 vccd1 vccd1 _13740_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16458_ _18371_/CLK _16458_/D vssd1 vssd1 vccd1 vccd1 _16458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15409_ hold529/X _15485_/A2 _15488_/A2 hold624/X _15408_/X vssd1 vssd1 vccd1 vccd1
+ _15412_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_6_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16389_ _18334_/CLK _16389_/D vssd1 vssd1 vccd1 vccd1 _16389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18128_ _18212_/CLK _18128_/D vssd1 vssd1 vccd1 vccd1 _18128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5706 _12348_/Y vssd1 vssd1 vccd1 vccd1 _12349_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5717 _17118_/Q vssd1 vssd1 vccd1 vccd1 hold5717/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5728 _13816_/Y vssd1 vssd1 vccd1 vccd1 _17725_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5739 _17615_/Q vssd1 vssd1 vccd1 vccd1 hold5739/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18059_ _18059_/CLK _18059_/D vssd1 vssd1 vccd1 vccd1 _18059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09901_ _09995_/A _10028_/B _09900_/X _08954_/A vssd1 vssd1 vccd1 vccd1 _09901_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout505 _10538_/S vssd1 vssd1 vccd1 vccd1 _11183_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_226_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout516 _10649_/C vssd1 vssd1 vccd1 vccd1 _10625_/C sky130_fd_sc_hd__clkbuf_8
X_09832_ hold4849/X _11171_/B _09831_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _09832_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout527 hold271/X vssd1 vssd1 vccd1 vccd1 _09283_/S sky130_fd_sc_hd__buf_6
XFILLER_0_67_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout538 _08868_/X vssd1 vssd1 vccd1 vccd1 _12501_/A3 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout549 hold114/X vssd1 vssd1 vccd1 vccd1 _08390_/S sky130_fd_sc_hd__clkbuf_8
X_09763_ hold3993/X _10049_/B _09762_/X _15146_/C1 vssd1 vssd1 vccd1 vccd1 _09763_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08714_ _12438_/A _08714_/B vssd1 vssd1 vccd1 vccd1 _15978_/D sky130_fd_sc_hd__and2_1
XFILLER_0_198_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09694_ hold4042/X _09992_/B _09693_/X _15202_/C1 vssd1 vssd1 vccd1 vccd1 _09694_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08645_ hold92/X hold487/X _08657_/S vssd1 vssd1 vccd1 vccd1 hold488/A sky130_fd_sc_hd__mux2_1
XFILLER_0_222_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08576_ hold53/X hold666/X _08592_/S vssd1 vssd1 vccd1 vccd1 _08577_/B sky130_fd_sc_hd__mux2_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_136_wb_clk_i clkbuf_6_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17347_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_194_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09128_ _15511_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09128_/X sky130_fd_sc_hd__or2_1
XFILLER_0_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09059_ _12420_/A hold546/X vssd1 vssd1 vccd1 vccd1 _16146_/D sky130_fd_sc_hd__and2_1
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12070_ hold4749/X _12356_/B _12069_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _12070_/X
+ sky130_fd_sc_hd__o211a_1
Xhold570 hold570/A vssd1 vssd1 vccd1 vccd1 hold570/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_241_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold581 hold581/A vssd1 vssd1 vccd1 vccd1 hold581/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold592 hold592/A vssd1 vssd1 vccd1 vccd1 hold592/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11021_ hold2666/X _16831_/Q _11183_/C vssd1 vssd1 vccd1 vccd1 _11022_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ _17744_/CLK _15760_/D vssd1 vssd1 vccd1 vccd1 _15760_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _12978_/A _12972_/B vssd1 vssd1 vccd1 vccd1 _17500_/D sky130_fd_sc_hd__and2_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_232_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1270 _09235_/X vssd1 vssd1 vccd1 vccd1 _09236_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ hold2049/X _14718_/B _14710_/X _14853_/C1 vssd1 vssd1 vccd1 vccd1 _14711_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1281 _17977_/Q vssd1 vssd1 vccd1 vccd1 hold1281/X sky130_fd_sc_hd__dlygate4sd3_1
X_11923_ hold5612/X _12305_/B _11922_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _11923_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_231_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1292 _08222_/X vssd1 vssd1 vccd1 vccd1 _15747_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15691_ _17878_/CLK _15691_/D vssd1 vssd1 vccd1 vccd1 _15691_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _15197_/A _14672_/B vssd1 vssd1 vccd1 vccd1 _14642_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ _17430_/CLK _17430_/D vssd1 vssd1 vccd1 vccd1 _17430_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11854_ hold5757/X _12332_/B _11853_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _11854_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10805_ hold2429/X hold3960/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10806_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14573_ hold307/X _14573_/B vssd1 vssd1 vccd1 vccd1 _14622_/B sky130_fd_sc_hd__nand2_8
X_17361_ _17517_/CLK _17361_/D vssd1 vssd1 vccd1 vccd1 _17361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11785_ _12331_/A _11785_/B vssd1 vssd1 vccd1 vccd1 _11785_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16312_ _18408_/CLK _16312_/D vssd1 vssd1 vccd1 vccd1 _16312_/Q sky130_fd_sc_hd__dfxtp_1
X_13524_ _13716_/A _13524_/B vssd1 vssd1 vccd1 vccd1 _13524_/X sky130_fd_sc_hd__or2_1
X_17292_ _17301_/CLK _17292_/D vssd1 vssd1 vccd1 vccd1 hold839/A sky130_fd_sc_hd__dfxtp_1
X_10736_ hold1402/X hold4356/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10737_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16243_ _17426_/CLK _16243_/D vssd1 vssd1 vccd1 vccd1 _16243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13455_ _13773_/A _13455_/B vssd1 vssd1 vccd1 vccd1 _13455_/X sky130_fd_sc_hd__or2_1
X_10667_ hold1746/X hold4328/X _11153_/C vssd1 vssd1 vccd1 vccd1 _10668_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12406_ _15364_/A hold702/X vssd1 vssd1 vccd1 vccd1 _17296_/D sky130_fd_sc_hd__and2_1
XFILLER_0_207_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16174_ _18400_/CLK _16174_/D vssd1 vssd1 vccd1 vccd1 _16174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13386_ _13482_/A _13386_/B vssd1 vssd1 vccd1 vccd1 _13386_/X sky130_fd_sc_hd__or2_1
XFILLER_0_51_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10598_ _10598_/A _10598_/B _11186_/C vssd1 vssd1 vccd1 vccd1 _10598_/X sky130_fd_sc_hd__and3_1
XFILLER_0_24_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15125_ _15233_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15125_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput108 hold5929/X vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_12
X_12337_ _12337_/A _12337_/B vssd1 vssd1 vccd1 vccd1 _12337_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_121_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput119 hold5965/X vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_12
XFILLER_0_51_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15056_ _15056_/A hold655/X vssd1 vssd1 vccd1 vccd1 _18313_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12268_ hold5761/X _12362_/B _12267_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _12268_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14007_ hold2205/X _14040_/B _14006_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _14007_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11219_ _16897_/Q _11222_/B _11219_/C vssd1 vssd1 vccd1 vccd1 _11219_/X sky130_fd_sc_hd__and3_1
XFILLER_0_235_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12199_ hold4937/X _12293_/B _12198_/X _12199_/C1 vssd1 vssd1 vccd1 vccd1 _12199_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput90 _13265_/A vssd1 vssd1 vccd1 vccd1 output90/X sky130_fd_sc_hd__buf_6
XFILLER_0_37_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15958_ _16129_/CLK _15958_/D vssd1 vssd1 vccd1 vccd1 _15958_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14909_ hold2390/X _14896_/Y _14908_/X _15042_/A vssd1 vssd1 vccd1 vccd1 _14909_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15889_ _17318_/CLK _15889_/D vssd1 vssd1 vccd1 vccd1 hold475/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_231_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08430_ hold2285/X _08433_/B _08429_/Y _08133_/A vssd1 vssd1 vccd1 vccd1 _08430_/X
+ sky130_fd_sc_hd__o211a_1
X_17628_ _17628_/CLK _17628_/D vssd1 vssd1 vccd1 vccd1 _17628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08361_ _08361_/A _08361_/B vssd1 vssd1 vccd1 vccd1 _15812_/D sky130_fd_sc_hd__and2_1
XFILLER_0_129_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17559_ _17719_/CLK _17559_/D vssd1 vssd1 vccd1 vccd1 _17559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08292_ hold2807/X _08336_/A2 _08291_/X _13729_/C1 vssd1 vssd1 vccd1 vccd1 _08292_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_229_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5503 _13363_/X vssd1 vssd1 vccd1 vccd1 _17574_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5514 _13474_/X vssd1 vssd1 vccd1 vccd1 _17611_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5525 _16937_/Q vssd1 vssd1 vccd1 vccd1 hold5525/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5536 _10810_/X vssd1 vssd1 vccd1 vccd1 _16760_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4802 _09634_/X vssd1 vssd1 vccd1 vccd1 _16368_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5547 _16902_/Q vssd1 vssd1 vccd1 vccd1 hold5547/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5558 _13564_/X vssd1 vssd1 vccd1 vccd1 _17641_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4813 _17628_/Q vssd1 vssd1 vccd1 vccd1 hold4813/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5569 _16842_/Q vssd1 vssd1 vccd1 vccd1 hold5569/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4824 _13636_/X vssd1 vssd1 vccd1 vccd1 _17665_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4835 _17130_/Q vssd1 vssd1 vccd1 vccd1 hold4835/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4846 _10876_/X vssd1 vssd1 vccd1 vccd1 _16782_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4857 _17187_/Q vssd1 vssd1 vccd1 vccd1 hold4857/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout302 _11106_/A vssd1 vssd1 vccd1 vccd1 _11010_/A sky130_fd_sc_hd__buf_4
XFILLER_0_121_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4868 _13450_/X vssd1 vssd1 vccd1 vccd1 _17603_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4879 _17622_/Q vssd1 vssd1 vccd1 vccd1 hold4879/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout313 _10986_/A vssd1 vssd1 vccd1 vccd1 _11091_/A sky130_fd_sc_hd__buf_4
XFILLER_0_121_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout324 _10560_/A vssd1 vssd1 vccd1 vccd1 _09978_/A sky130_fd_sc_hd__buf_4
Xfanout335 fanout335/A vssd1 vssd1 vccd1 vccd1 _10542_/A sky130_fd_sc_hd__buf_4
XFILLER_0_10_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout346 _09056_/S vssd1 vssd1 vccd1 vccd1 _09060_/S sky130_fd_sc_hd__buf_8
Xfanout357 _08623_/S vssd1 vssd1 vccd1 vccd1 _08657_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_226_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09815_ hold1624/X _16429_/Q _10025_/C vssd1 vssd1 vccd1 vccd1 _09816_/B sky130_fd_sc_hd__mux2_1
Xfanout368 _15127_/Y vssd1 vssd1 vccd1 vccd1 _15165_/B sky130_fd_sc_hd__clkbuf_8
Xfanout379 _14912_/Y vssd1 vssd1 vccd1 vccd1 _14946_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_213_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09746_ hold2751/X _16406_/Q _10040_/C vssd1 vssd1 vccd1 vccd1 _09747_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_388_wb_clk_i clkbuf_6_35_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17204_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_213_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09677_ hold1483/X _16383_/Q _10385_/S vssd1 vssd1 vccd1 vccd1 _09678_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_317_wb_clk_i clkbuf_6_47_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18070_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08628_ _15364_/A hold607/X vssd1 vssd1 vccd1 vccd1 _15936_/D sky130_fd_sc_hd__and2_1
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08559_ _12426_/A hold505/X vssd1 vssd1 vccd1 vccd1 _15903_/D sky130_fd_sc_hd__and2_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11570_ hold3049/X hold4947/X _11660_/S vssd1 vssd1 vccd1 vccd1 _11571_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_9_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10521_ _11103_/A _10521_/B vssd1 vssd1 vccd1 vccd1 _10521_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13240_ _13233_/X _13239_/X _13296_/B1 vssd1 vssd1 vccd1 vccd1 _17548_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_208_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10452_ _10551_/A _10452_/B vssd1 vssd1 vccd1 vccd1 _10452_/X sky130_fd_sc_hd__or2_1
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13171_ _13170_/X hold5999/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13171_/X sky130_fd_sc_hd__mux2_1
X_10383_ _10986_/A _10383_/B vssd1 vssd1 vccd1 vccd1 _10383_/X sky130_fd_sc_hd__or2_1
X_12122_ hold1344/X hold4061/X _12323_/C vssd1 vssd1 vccd1 vccd1 _12123_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_33_wb_clk_i clkbuf_6_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18432_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_206_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_236_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12053_ hold1358/X _17175_/Q _12371_/C vssd1 vssd1 vccd1 vccd1 _12054_/B sky130_fd_sc_hd__mux2_1
X_16930_ _17905_/CLK _16930_/D vssd1 vssd1 vccd1 vccd1 _16930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11004_ _11661_/A _11004_/B vssd1 vssd1 vccd1 vccd1 _11004_/X sky130_fd_sc_hd__or2_1
X_16861_ _17973_/CLK _16861_/D vssd1 vssd1 vccd1 vccd1 _16861_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout880 _15145_/A vssd1 vssd1 vccd1 vccd1 hold2105/A sky130_fd_sc_hd__buf_6
XFILLER_0_205_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout891 hold423/X vssd1 vssd1 vccd1 vccd1 _15085_/A sky130_fd_sc_hd__buf_12
X_15812_ _17689_/CLK _15812_/D vssd1 vssd1 vccd1 vccd1 _15812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16792_ _18059_/CLK _16792_/D vssd1 vssd1 vccd1 vccd1 _16792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12955_ hold2769/X hold3239/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12955_/X sky130_fd_sc_hd__mux2_1
X_15743_ _17746_/CLK _15743_/D vssd1 vssd1 vccd1 vccd1 _15743_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11906_ hold1716/X _17126_/Q _13796_/S vssd1 vssd1 vccd1 vccd1 _11907_/B sky130_fd_sc_hd__mux2_1
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18462_ _18462_/CLK _18462_/D vssd1 vssd1 vccd1 vccd1 _18462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15674_ _17262_/CLK _15674_/D vssd1 vssd1 vccd1 vccd1 _15674_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ hold2193/X hold3147/X _12916_/S vssd1 vssd1 vccd1 vccd1 _12886_/X sky130_fd_sc_hd__mux2_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _17754_/CLK _17413_/D vssd1 vssd1 vccd1 vccd1 _17413_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14625_ hold959/X _14612_/B _14624_/X _15218_/C1 vssd1 vssd1 vccd1 vccd1 hold960/A
+ sky130_fd_sc_hd__o211a_1
X_11837_ hold2428/X hold4315/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11838_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18393_ _18393_/CLK _18393_/D vssd1 vssd1 vccd1 vccd1 _18393_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _17344_/CLK hold9/X vssd1 vssd1 vccd1 vccd1 _17344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14556_ _14556_/A hold353/A hold361/A vssd1 vssd1 vccd1 vccd1 _14843_/B sky130_fd_sc_hd__or3_4
XFILLER_0_138_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11768_ _17080_/Q _11789_/B _11789_/C vssd1 vssd1 vccd1 vccd1 _11768_/X sky130_fd_sc_hd__and3_1
XFILLER_0_16_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10719_ _11127_/A _10719_/B vssd1 vssd1 vccd1 vccd1 _10719_/X sky130_fd_sc_hd__or2_1
X_13507_ hold3909/X _13795_/A2 _13506_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13507_/X
+ sky130_fd_sc_hd__o211a_1
X_14487_ _15547_/A _14487_/B vssd1 vssd1 vccd1 vccd1 _14487_/Y sky130_fd_sc_hd__nand2_1
X_17275_ _17741_/CLK _17275_/D vssd1 vssd1 vccd1 vccd1 _17275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11699_ hold1231/X hold4953/X _12173_/S vssd1 vssd1 vccd1 vccd1 _11700_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13438_ hold4758/X _13829_/B _13437_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13438_/X
+ sky130_fd_sc_hd__o211a_1
X_16226_ _18458_/CLK _16226_/D vssd1 vssd1 vccd1 vccd1 _16226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16157_ _17506_/CLK _16157_/D vssd1 vssd1 vccd1 vccd1 _16157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13369_ hold4077/X _13847_/B _13368_/X _13765_/C1 vssd1 vssd1 vccd1 vccd1 _13369_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4109 _16956_/Q vssd1 vssd1 vccd1 vccd1 hold4109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15108_ hold2752/X hold341/X _15107_/Y _15048_/A vssd1 vssd1 vccd1 vccd1 _15108_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16088_ _17337_/CLK _16088_/D vssd1 vssd1 vccd1 vccd1 _16088_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3408 _16346_/Q vssd1 vssd1 vccd1 vccd1 _13238_/A sky130_fd_sc_hd__buf_1
XFILLER_0_80_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_224_1295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3419 _10056_/Y vssd1 vssd1 vccd1 vccd1 _10057_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_107_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15039_ hold951/X hold1399/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15040_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07930_ _15553_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07930_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2707 _18001_/Q vssd1 vssd1 vccd1 vccd1 hold2707/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2718 _15805_/Q vssd1 vssd1 vccd1 vccd1 hold2718/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2729 _17940_/Q vssd1 vssd1 vccd1 vccd1 hold2729/X sky130_fd_sc_hd__dlygate4sd3_1
X_07861_ _15539_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07861_/X sky130_fd_sc_hd__or2_1
XFILLER_0_236_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09600_ _09912_/A _09600_/B vssd1 vssd1 vccd1 vccd1 _09600_/X sky130_fd_sc_hd__or2_1
XFILLER_0_177_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07792_ _07809_/B vssd1 vssd1 vccd1 vccd1 _09339_/B sky130_fd_sc_hd__inv_2
XFILLER_0_190_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09531_ _09981_/A _09531_/B vssd1 vssd1 vccd1 vccd1 _09531_/X sky130_fd_sc_hd__or2_1
XFILLER_0_155_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_1356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_410_wb_clk_i clkbuf_6_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17167_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_211_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09462_ _09461_/X _09478_/B _09462_/C vssd1 vssd1 vccd1 vccd1 _16314_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_17_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08413_ _14413_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08413_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09393_ _07805_/Y _09362_/A _09369_/D _09392_/X vssd1 vssd1 vccd1 vccd1 _09393_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08344_ hold911/X hold1632/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08345_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08275_ hold2589/X _08268_/B _08274_/X _12804_/A vssd1 vssd1 vccd1 vccd1 _08275_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6001 _16532_/Q vssd1 vssd1 vccd1 vccd1 hold6001/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6012 _17542_/Q vssd1 vssd1 vccd1 vccd1 hold6012/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6023 _17546_/Q vssd1 vssd1 vccd1 vccd1 hold6023/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6034 _17529_/Q vssd1 vssd1 vccd1 vccd1 hold6034/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6045 data_in[18] vssd1 vssd1 vccd1 vccd1 hold242/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5300 _11467_/X vssd1 vssd1 vccd1 vccd1 _16979_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold6056 _16211_/Q vssd1 vssd1 vccd1 vccd1 hold6056/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5311 _17087_/Q vssd1 vssd1 vccd1 vccd1 hold5311/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5322 _11566_/X vssd1 vssd1 vccd1 vccd1 _17012_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold6067 _16276_/Q vssd1 vssd1 vccd1 vccd1 hold6067/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6078 data_in[27] vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5333 _17055_/Q vssd1 vssd1 vccd1 vccd1 hold5333/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5344 _10909_/X vssd1 vssd1 vccd1 vccd1 _16793_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4610 _16499_/Q vssd1 vssd1 vccd1 vccd1 hold4610/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6089 _18413_/Q vssd1 vssd1 vccd1 vccd1 hold6089/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5355 _17672_/Q vssd1 vssd1 vccd1 vccd1 hold5355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4621 _10357_/X vssd1 vssd1 vccd1 vccd1 _16609_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5366 _16861_/Q vssd1 vssd1 vccd1 vccd1 hold5366/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4632 _16706_/Q vssd1 vssd1 vccd1 vccd1 hold4632/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5377 _11446_/X vssd1 vssd1 vccd1 vccd1 _16972_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5388 _16756_/Q vssd1 vssd1 vccd1 vccd1 hold5388/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4643 _13444_/X vssd1 vssd1 vccd1 vccd1 _17601_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4654 _17160_/Q vssd1 vssd1 vccd1 vccd1 hold4654/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5399 _10840_/X vssd1 vssd1 vccd1 vccd1 _16770_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4665 _13351_/X vssd1 vssd1 vccd1 vccd1 _17570_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3920 _11125_/X vssd1 vssd1 vccd1 vccd1 _16865_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4676 _17558_/Q vssd1 vssd1 vccd1 vccd1 hold4676/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3931 _17265_/Q vssd1 vssd1 vccd1 vccd1 _12323_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4687 _16409_/Q vssd1 vssd1 vccd1 vccd1 hold4687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3942 _16885_/Q vssd1 vssd1 vccd1 vccd1 hold3942/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3953 _13609_/X vssd1 vssd1 vccd1 vccd1 _17656_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4698 _13333_/X vssd1 vssd1 vccd1 vccd1 _17564_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3964 _17409_/Q vssd1 vssd1 vccd1 vccd1 hold3964/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3975 _10417_/X vssd1 vssd1 vccd1 vccd1 _16629_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout154 _12905_/S vssd1 vssd1 vccd1 vccd1 _12923_/S sky130_fd_sc_hd__buf_6
Xhold3986 _10765_/X vssd1 vssd1 vccd1 vccd1 _16745_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout165 _12217_/A2 vssd1 vssd1 vccd1 vccd1 _13817_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_227_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3997 _16597_/Q vssd1 vssd1 vccd1 vccd1 hold3997/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout176 _11723_/B vssd1 vssd1 vccd1 vccd1 _11732_/B sky130_fd_sc_hd__buf_4
XFILLER_0_22_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout187 fanout210/X vssd1 vssd1 vccd1 vccd1 _13868_/B sky130_fd_sc_hd__clkbuf_4
Xfanout198 _11786_/B vssd1 vssd1 vccd1 vccd1 _12329_/B sky130_fd_sc_hd__buf_4
XFILLER_0_96_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09729_ _11010_/A _09729_/B vssd1 vssd1 vccd1 vccd1 _09729_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_151_wb_clk_i clkbuf_6_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18242_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12740_ hold3177/X _12739_/X _12749_/S vssd1 vssd1 vccd1 vccd1 _12741_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ hold3122/X _12670_/X _12851_/S vssd1 vssd1 vccd1 vccd1 _12671_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ hold994/X _14446_/A2 _14409_/X _14344_/A vssd1 vssd1 vccd1 vccd1 hold995/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _11622_/A _11622_/B vssd1 vssd1 vccd1 vccd1 _11622_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15390_ hold625/X _15448_/A2 _15446_/B1 hold728/X vssd1 vssd1 vccd1 vccd1 _15390_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14341_ hold927/X hold2008/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14342_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_147_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11553_ _11553_/A _11553_/B vssd1 vssd1 vccd1 vccd1 _11553_/X sky130_fd_sc_hd__or2_1
XFILLER_0_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10504_ _10598_/A _10070_/B _10503_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10504_/X
+ sky130_fd_sc_hd__o211a_1
X_17060_ _17908_/CLK _17060_/D vssd1 vssd1 vccd1 vccd1 _17060_/Q sky130_fd_sc_hd__dfxtp_1
X_14272_ _15221_/A _14272_/B vssd1 vssd1 vccd1 vccd1 _14272_/Y sky130_fd_sc_hd__nand2_1
X_11484_ _12243_/A _11484_/B vssd1 vssd1 vccd1 vccd1 _11484_/X sky130_fd_sc_hd__or2_1
X_16011_ _18418_/CLK _16011_/D vssd1 vssd1 vccd1 vccd1 hold458/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13223_ _13311_/A1 _13221_/X _13222_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13223_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_21_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10435_ hold3251/X _10625_/B _10434_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _10435_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13154_ _17570_/Q _17104_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13154_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_221_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10366_ hold3882/X _10070_/B _10365_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _10366_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _13716_/A _12105_/B vssd1 vssd1 vccd1 vccd1 _12105_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _13084_/X hold3417/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13085_/X sky130_fd_sc_hd__mux2_1
X_17962_ _18126_/CLK _17962_/D vssd1 vssd1 vccd1 vccd1 _17962_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10297_ hold4024/X _10619_/B _10296_/X _14853_/C1 vssd1 vssd1 vccd1 vccd1 _10297_/X
+ sky130_fd_sc_hd__o211a_1
X_12036_ _12234_/A _12036_/B vssd1 vssd1 vccd1 vccd1 _12036_/X sky130_fd_sc_hd__or2_1
X_16913_ _17838_/CLK _16913_/D vssd1 vssd1 vccd1 vccd1 _16913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_239_wb_clk_i clkbuf_6_60_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18129_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17893_ _17895_/CLK _17893_/D vssd1 vssd1 vccd1 vccd1 _17893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_217_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16844_ _17983_/CLK _16844_/D vssd1 vssd1 vccd1 vccd1 _16844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16775_ _18010_/CLK _16775_/D vssd1 vssd1 vccd1 vccd1 _16775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13987_ hold2363/X _13986_/B _13986_/Y _13941_/A vssd1 vssd1 vccd1 vccd1 _13987_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15726_ _17697_/CLK _15726_/D vssd1 vssd1 vccd1 vccd1 _15726_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ hold4535/X _12937_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12939_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_137_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18445_ _18445_/CLK _18445_/D vssd1 vssd1 vccd1 vccd1 _18445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15657_ _17902_/CLK _15657_/D vssd1 vssd1 vccd1 vccd1 _15657_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ hold3300/X _12868_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12870_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_145_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14608_ _15163_/A _14612_/B vssd1 vssd1 vccd1 vccd1 _14608_/Y sky130_fd_sc_hd__nand2_1
X_18376_ _18376_/CLK _18376_/D vssd1 vssd1 vccd1 vccd1 _18376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15588_ _17204_/CLK _15588_/D vssd1 vssd1 vccd1 vccd1 _15588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17327_ _17331_/CLK hold3/X vssd1 vssd1 vccd1 vccd1 _17327_/Q sky130_fd_sc_hd__dfxtp_1
X_14539_ _15165_/A _14541_/B vssd1 vssd1 vccd1 vccd1 _14539_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08060_ _15519_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08060_/X sky130_fd_sc_hd__or2_1
XFILLER_0_154_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17258_ _18445_/CLK _17258_/D vssd1 vssd1 vccd1 vccd1 _17258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16209_ _17440_/CLK hold987/X vssd1 vssd1 vccd1 vccd1 hold986/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17189_ _17221_/CLK _17189_/D vssd1 vssd1 vccd1 vccd1 _17189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3205 _10044_/Y vssd1 vssd1 vccd1 vccd1 _10045_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3216 _16415_/Q vssd1 vssd1 vccd1 vccd1 hold3216/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08962_ _12426_/A hold589/X vssd1 vssd1 vccd1 vccd1 _16098_/D sky130_fd_sc_hd__and2_1
Xhold3227 _12758_/X vssd1 vssd1 vccd1 vccd1 _12759_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3238 _09571_/X vssd1 vssd1 vccd1 vccd1 _16347_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3249 _16489_/Q vssd1 vssd1 vccd1 vccd1 _09995_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2504 _08095_/X vssd1 vssd1 vccd1 vccd1 _15687_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2515 _14231_/X vssd1 vssd1 vccd1 vccd1 _17917_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07913_ hold1825/X _07918_/B _07912_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _07913_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2526 _17824_/Q vssd1 vssd1 vccd1 vccd1 hold2526/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08893_ _15314_/A hold731/X vssd1 vssd1 vccd1 vccd1 _16064_/D sky130_fd_sc_hd__and2_1
Xhold2537 _15593_/Q vssd1 vssd1 vccd1 vccd1 hold2537/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2548 _18280_/Q vssd1 vssd1 vccd1 vccd1 hold2548/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1803 _18399_/Q vssd1 vssd1 vccd1 vccd1 hold1803/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2559 _15793_/Q vssd1 vssd1 vccd1 vccd1 hold2559/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1814 _15493_/X vssd1 vssd1 vccd1 vccd1 _15494_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1825 _15600_/Q vssd1 vssd1 vccd1 vccd1 hold1825/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1836 _14915_/X vssd1 vssd1 vccd1 vccd1 _18244_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07844_ hold2426/X _07869_/B _07843_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _07844_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1847 _18376_/Q vssd1 vssd1 vccd1 vccd1 hold1847/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1858 _15196_/X vssd1 vssd1 vccd1 vccd1 _18380_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1869 _18387_/Q vssd1 vssd1 vccd1 vccd1 hold1869/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_6_17_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_17_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_190_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09514_ hold4677/X _09992_/B _09513_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _09514_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_231_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09445_ _09447_/C _09447_/D _09447_/B vssd1 vssd1 vccd1 vccd1 _09446_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_148_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09376_ hold813/X _15483_/B _09375_/X _07809_/B vssd1 vssd1 vccd1 vccd1 _09376_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08327_ _14330_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08327_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08258_ _14477_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08258_/X sky130_fd_sc_hd__or2_1
XFILLER_0_144_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08189_ _14517_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08189_/X sky130_fd_sc_hd__or2_1
Xhold5130 _11935_/X vssd1 vssd1 vccd1 vccd1 _17135_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10220_ hold2019/X _16564_/Q _10646_/C vssd1 vssd1 vccd1 vccd1 _10221_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5141 _11368_/X vssd1 vssd1 vccd1 vccd1 _16946_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5152 _16887_/Q vssd1 vssd1 vccd1 vccd1 hold5152/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5163 _16516_/Q vssd1 vssd1 vccd1 vccd1 hold5163/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5174 _11083_/X vssd1 vssd1 vccd1 vccd1 _16851_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5185 _16504_/Q vssd1 vssd1 vccd1 vccd1 hold5185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4440 _12325_/Y vssd1 vssd1 vccd1 vccd1 _17265_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10151_ hold2594/X hold3463/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10152_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_6_56_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_56_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
Xhold4451 _11788_/Y vssd1 vssd1 vccd1 vccd1 _17086_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5196 _11560_/X vssd1 vssd1 vccd1 vccd1 _17010_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4462 _10150_/X vssd1 vssd1 vccd1 vccd1 _16540_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4473 _12307_/Y vssd1 vssd1 vccd1 vccd1 _17259_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4484 _16364_/Q vssd1 vssd1 vccd1 vccd1 hold4484/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3750 _16361_/Q vssd1 vssd1 vccd1 vccd1 hold3750/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_234_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4495 _17577_/Q vssd1 vssd1 vccd1 vccd1 hold4495/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3761 _16666_/Q vssd1 vssd1 vccd1 vccd1 hold3761/X sky130_fd_sc_hd__dlygate4sd3_1
X_10082_ _18076_/Q _16518_/Q _10634_/C vssd1 vssd1 vccd1 vccd1 _10083_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_332_wb_clk_i clkbuf_6_41_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17144_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3772 _10954_/X vssd1 vssd1 vccd1 vccd1 _16808_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3783 _17416_/Q vssd1 vssd1 vccd1 vccd1 hold3783/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3794 _12701_/X vssd1 vssd1 vccd1 vccd1 _12702_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13910_ _15145_/A hold2256/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13911_/B sky130_fd_sc_hd__mux2_1
XTAP_5978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14890_ _15229_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14890_/X sky130_fd_sc_hd__or2_1
XTAP_5989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13841_ _17734_/Q _13847_/B _13841_/C vssd1 vssd1 vccd1 vccd1 _13841_/X sky130_fd_sc_hd__and3_1
XFILLER_0_57_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_230_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16560_ _18150_/CLK _16560_/D vssd1 vssd1 vccd1 vccd1 _16560_/Q sky130_fd_sc_hd__dfxtp_1
X_13772_ hold2749/X hold5396/X _13865_/C vssd1 vssd1 vccd1 vccd1 _13773_/B sky130_fd_sc_hd__mux2_1
X_10984_ hold5119/X _11210_/B _10983_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _10984_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15511_ _15511_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15511_/X sky130_fd_sc_hd__or2_1
XFILLER_0_214_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12723_ _12810_/A _12723_/B vssd1 vssd1 vccd1 vccd1 _17417_/D sky130_fd_sc_hd__and2_1
X_16491_ _17535_/CLK _16491_/D vssd1 vssd1 vccd1 vccd1 _16491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18230_ _18231_/CLK _18230_/D vssd1 vssd1 vccd1 vccd1 _18230_/Q sky130_fd_sc_hd__dfxtp_1
X_15442_ _15480_/A _15442_/B _15442_/C _15442_/D vssd1 vssd1 vccd1 vccd1 _15442_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_167_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12654_ _12873_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _17394_/D sky130_fd_sc_hd__and2_1
XFILLER_0_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11605_ hold4953/X _11798_/B _11604_/X _14143_/C1 vssd1 vssd1 vccd1 vccd1 _11605_/X
+ sky130_fd_sc_hd__o211a_1
X_18161_ _18212_/CLK _18161_/D vssd1 vssd1 vccd1 vccd1 _18161_/Q sky130_fd_sc_hd__dfxtp_1
X_15373_ _15490_/A1 _15365_/X _15372_/X _15490_/B1 _18413_/Q vssd1 vssd1 vccd1 vccd1
+ _15373_/X sky130_fd_sc_hd__a32o_1
X_12585_ _12894_/A _12585_/B vssd1 vssd1 vccd1 vccd1 _17371_/D sky130_fd_sc_hd__and2_1
XFILLER_0_108_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17112_ _17144_/CLK _17112_/D vssd1 vssd1 vccd1 vccd1 _17112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14324_ _15165_/A _14326_/B vssd1 vssd1 vccd1 vccd1 _14324_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11536_ hold5440/X _11726_/B _11535_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _11536_/X
+ sky130_fd_sc_hd__o211a_1
X_18092_ _18124_/CLK _18092_/D vssd1 vssd1 vccd1 vccd1 _18092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14255_ hold2794/X _14272_/B _14254_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14255_/X
+ sky130_fd_sc_hd__o211a_1
X_17043_ _17891_/CLK _17043_/D vssd1 vssd1 vccd1 vccd1 _17043_/Q sky130_fd_sc_hd__dfxtp_1
X_11467_ hold5299/X _11753_/B _11466_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11467_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13206_ _13206_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13206_/X sky130_fd_sc_hd__or2_1
XFILLER_0_238_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10418_ hold2920/X _16630_/Q _10628_/C vssd1 vssd1 vccd1 vccd1 _10419_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_0_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14186_ _14596_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14186_/X sky130_fd_sc_hd__or2_1
X_11398_ hold4101/X _11741_/B _11397_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _11398_/X
+ sky130_fd_sc_hd__o211a_1
X_13137_ _13137_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13137_/X sky130_fd_sc_hd__and2_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10349_ hold1839/X _16607_/Q _10595_/C vssd1 vssd1 vccd1 vccd1 _10350_/B sky130_fd_sc_hd__mux2_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ hold4634/X _13067_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13068_/X sky130_fd_sc_hd__mux2_2
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _17949_/CLK _17945_/D vssd1 vssd1 vccd1 vccd1 _17945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_224_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12019_ hold5543/X _12305_/B _12018_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _12019_/X
+ sky130_fd_sc_hd__o211a_1
X_17876_ _17908_/CLK _17876_/D vssd1 vssd1 vccd1 vccd1 _17876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_219_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_219_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16827_ _18030_/CLK _16827_/D vssd1 vssd1 vccd1 vccd1 _16827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16758_ _18023_/CLK _16758_/D vssd1 vssd1 vccd1 vccd1 _16758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15709_ _17202_/CLK _15709_/D vssd1 vssd1 vccd1 vccd1 _15709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16689_ _18087_/CLK _16689_/D vssd1 vssd1 vccd1 vccd1 _16689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09230_ _15559_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09230_/X sky130_fd_sc_hd__or2_1
XFILLER_0_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18428_ _18428_/CLK _18428_/D vssd1 vssd1 vccd1 vccd1 _18428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09161_ hold2562/X _09164_/B _09160_/Y _12906_/A vssd1 vssd1 vccd1 vccd1 _09161_/X
+ sky130_fd_sc_hd__o211a_1
X_18359_ _18395_/CLK _18359_/D vssd1 vssd1 vccd1 vccd1 _18359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08112_ _15517_/A hold2428/X hold108/X vssd1 vssd1 vccd1 vccd1 _08113_/B sky130_fd_sc_hd__mux2_1
X_09092_ _15099_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _09092_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08043_ _15557_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08043_/X sky130_fd_sc_hd__or2_1
XFILLER_0_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold900 hold900/A vssd1 vssd1 vccd1 vccd1 hold900/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 hold911/A vssd1 vssd1 vccd1 vccd1 hold911/X sky130_fd_sc_hd__buf_12
Xhold922 hold922/A vssd1 vssd1 vccd1 vccd1 hold922/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold933 hold933/A vssd1 vssd1 vccd1 vccd1 hold933/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold944 hold976/X vssd1 vssd1 vccd1 vccd1 hold944/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold955 hold955/A vssd1 vssd1 vccd1 vccd1 hold955/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 hold966/A vssd1 vssd1 vccd1 vccd1 input68/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_229_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold977 hold977/A vssd1 vssd1 vccd1 vccd1 hold977/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3002 _18028_/Q vssd1 vssd1 vccd1 vccd1 hold3002/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3013 _14089_/X vssd1 vssd1 vccd1 vccd1 _17849_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ _11158_/A _09994_/B vssd1 vssd1 vccd1 vccd1 _16488_/D sky130_fd_sc_hd__nor2_1
Xhold988 hold988/A vssd1 vssd1 vccd1 vccd1 hold988/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3024 _14442_/X vssd1 vssd1 vccd1 vccd1 _18019_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 hold999/A vssd1 vssd1 vccd1 vccd1 hold999/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3035 _17907_/Q vssd1 vssd1 vccd1 vccd1 hold3035/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2301 _14609_/X vssd1 vssd1 vccd1 vccd1 _18098_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3046 _14743_/X vssd1 vssd1 vccd1 vccd1 _18162_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3057 _16184_/Q vssd1 vssd1 vccd1 vccd1 hold3057/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2312 _17798_/Q vssd1 vssd1 vccd1 vccd1 hold2312/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08945_ hold147/X hold796/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08946_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2323 _08184_/X vssd1 vssd1 vccd1 vccd1 _15728_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3068 _17865_/Q vssd1 vssd1 vccd1 vccd1 hold3068/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2334 _08512_/X vssd1 vssd1 vccd1 vccd1 _15883_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3079 _08247_/X vssd1 vssd1 vccd1 vccd1 _15758_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1600 _15639_/Q vssd1 vssd1 vccd1 vccd1 hold1600/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2345 _18326_/Q vssd1 vssd1 vccd1 vccd1 hold2345/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2356 _08518_/X vssd1 vssd1 vccd1 vccd1 _15886_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1611 _17898_/Q vssd1 vssd1 vccd1 vccd1 hold1611/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08876_ hold684/X hold874/X _08930_/S vssd1 vssd1 vccd1 vccd1 hold875/A sky130_fd_sc_hd__mux2_1
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2367 _15858_/Q vssd1 vssd1 vccd1 vccd1 hold2367/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1622 _16176_/Q vssd1 vssd1 vccd1 vccd1 hold1622/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2378 _17517_/Q vssd1 vssd1 vccd1 vccd1 hold2378/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1633 _15726_/Q vssd1 vssd1 vccd1 vccd1 hold1633/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2389 _08404_/X vssd1 vssd1 vccd1 vccd1 _15832_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1644 _15560_/X vssd1 vssd1 vccd1 vccd1 _18458_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1655 _09233_/X vssd1 vssd1 vccd1 vccd1 _09234_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07827_ hold444/A hold405/A hold337/A hold509/A vssd1 vssd1 vccd1 vccd1 hold330/A
+ sky130_fd_sc_hd__or4b_2
Xhold1666 _16216_/Q vssd1 vssd1 vccd1 vccd1 hold1666/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1677 _13989_/X vssd1 vssd1 vccd1 vccd1 _17801_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1688 _18024_/Q vssd1 vssd1 vccd1 vccd1 hold1688/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1699 _14167_/X vssd1 vssd1 vccd1 vccd1 _17886_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09428_ hold704/X _16300_/Q vssd1 vssd1 vccd1 vccd1 _09428_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09359_ hold97/X _15165_/A _09359_/C vssd1 vssd1 vccd1 vccd1 _09366_/C sky130_fd_sc_hd__or3_2
XFILLER_0_192_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12370_ _13888_/A _12370_/B vssd1 vssd1 vccd1 vccd1 _12370_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_209_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11321_ hold1613/X hold4506/X _12335_/C vssd1 vssd1 vccd1 vccd1 _11322_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_160_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14040_ _15221_/A _14040_/B vssd1 vssd1 vccd1 vccd1 _14040_/Y sky130_fd_sc_hd__nand2_1
X_11252_ hold2055/X hold4419/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11253_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10203_ _10413_/A _10203_/B vssd1 vssd1 vccd1 vccd1 _10203_/X sky130_fd_sc_hd__or2_1
XFILLER_0_197_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11183_ _16885_/Q _11225_/B _11183_/C vssd1 vssd1 vccd1 vccd1 _11183_/X sky130_fd_sc_hd__and3_1
XTAP_6421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4270 _17564_/Q vssd1 vssd1 vccd1 vccd1 hold4270/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10134_ _10542_/A _10134_/B vssd1 vssd1 vccd1 vccd1 _10134_/X sky130_fd_sc_hd__or2_1
XTAP_6443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4281 _16717_/Q vssd1 vssd1 vccd1 vccd1 hold4281/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4292 _12328_/Y vssd1 vssd1 vccd1 vccd1 _17266_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15991_ _17325_/CLK _15991_/D vssd1 vssd1 vccd1 vccd1 hold593/A sky130_fd_sc_hd__dfxtp_1
XTAP_5720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_237_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3580 _16493_/Q vssd1 vssd1 vccd1 vccd1 hold3580/X sky130_fd_sc_hd__dlygate4sd3_1
X_17730_ _17730_/CLK _17730_/D vssd1 vssd1 vccd1 vccd1 _17730_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14942_ hold630/X hold407/X vssd1 vssd1 vccd1 vccd1 _14942_/X sky130_fd_sc_hd__or2_1
XTAP_5753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10065_ _13286_/A _10476_/A _10064_/X vssd1 vssd1 vccd1 vccd1 _10065_/Y sky130_fd_sc_hd__a21oi_1
Xhold3591 _11196_/Y vssd1 vssd1 vccd1 vccd1 _11197_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17661_ _17661_/CLK _17661_/D vssd1 vssd1 vccd1 vccd1 _17661_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2890 _17758_/Q vssd1 vssd1 vccd1 vccd1 hold2890/X sky130_fd_sc_hd__dlygate4sd3_1
X_14873_ hold1714/X _14880_/B _14872_/X _14893_/C1 vssd1 vssd1 vccd1 vccd1 _14873_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16612_ _18222_/CLK _16612_/D vssd1 vssd1 vccd1 vccd1 _16612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13824_ hold4262/X _13794_/A _13823_/X vssd1 vssd1 vccd1 vccd1 _13825_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_216_1356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17592_ _17624_/CLK _17592_/D vssd1 vssd1 vccd1 vccd1 _17592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16543_ _18229_/CLK _16543_/D vssd1 vssd1 vccd1 vccd1 _16543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10967_ hold1964/X _16813_/Q _11162_/C vssd1 vssd1 vccd1 vccd1 _10968_/B sky130_fd_sc_hd__mux2_1
X_13755_ _13791_/A _13755_/B vssd1 vssd1 vccd1 vccd1 _13755_/X sky130_fd_sc_hd__or2_1
XFILLER_0_58_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12706_ hold917/X _17413_/Q _12766_/S vssd1 vssd1 vccd1 vccd1 _12706_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16474_ _18387_/CLK _16474_/D vssd1 vssd1 vccd1 vccd1 _16474_/Q sky130_fd_sc_hd__dfxtp_1
X_10898_ hold2713/X _16790_/Q _11186_/C vssd1 vssd1 vccd1 vccd1 _10899_/B sky130_fd_sc_hd__mux2_1
X_13686_ _13791_/A _13686_/B vssd1 vssd1 vccd1 vccd1 _13686_/X sky130_fd_sc_hd__or2_1
XFILLER_0_167_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18213_ _18213_/CLK _18213_/D vssd1 vssd1 vccd1 vccd1 _18213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15425_ _15425_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15425_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12637_ hold3089/X _17390_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12637_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_143_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18144_ _18176_/CLK _18144_/D vssd1 vssd1 vccd1 vccd1 _18144_/Q sky130_fd_sc_hd__dfxtp_1
X_15356_ _17339_/Q _15486_/B1 _09362_/D hold686/X vssd1 vssd1 vccd1 vccd1 _15356_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12568_ hold1400/X hold3220/X _12925_/S vssd1 vssd1 vccd1 vccd1 _12568_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14307_ hold1674/X _14333_/A2 _14306_/X _14372_/A vssd1 vssd1 vccd1 vccd1 _14307_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11519_ hold2771/X _16997_/Q _11717_/C vssd1 vssd1 vccd1 vccd1 _11520_/B sky130_fd_sc_hd__mux2_1
X_18075_ _18393_/CLK hold916/X vssd1 vssd1 vccd1 vccd1 _18075_/Q sky130_fd_sc_hd__dfxtp_1
X_12499_ hold35/X _12509_/A2 _12501_/A3 _12498_/X _09061_/A vssd1 vssd1 vccd1 vccd1
+ hold36/A sky130_fd_sc_hd__o311a_1
X_15287_ hold156/X _15487_/A2 _15484_/B1 hold94/X _15286_/X vssd1 vssd1 vccd1 vccd1
+ _15292_/B sky130_fd_sc_hd__a221o_1
Xhold207 hold207/A vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_184_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold218 hold218/A vssd1 vssd1 vccd1 vccd1 input46/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 hold383/X vssd1 vssd1 vccd1 vccd1 hold384/A sky130_fd_sc_hd__buf_6
X_17026_ _17905_/CLK _17026_/D vssd1 vssd1 vccd1 vccd1 _17026_/Q sky130_fd_sc_hd__dfxtp_1
X_14238_ _14972_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14238_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_254_wb_clk_i clkbuf_6_58_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17960_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14169_ hold1962/X _14198_/B _14168_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _14169_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout709 _12394_/A vssd1 vssd1 vccd1 vccd1 _15324_/A sky130_fd_sc_hd__clkbuf_4
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08730_ _08730_/A _08934_/A vssd1 vssd1 vccd1 vccd1 _08735_/S sky130_fd_sc_hd__or2_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _17960_/CLK _17928_/D vssd1 vssd1 vccd1 vccd1 _17928_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08661_ hold278/X hold861/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold862/A sky130_fd_sc_hd__mux2_1
XFILLER_0_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17859_ _17859_/CLK _17859_/D vssd1 vssd1 vccd1 vccd1 _17859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08592_ hold320/X hold872/X _08592_/S vssd1 vssd1 vccd1 vccd1 _08593_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_88_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09213_ hold2954/X _09214_/B _09212_/Y _12822_/A vssd1 vssd1 vccd1 vccd1 _09213_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09144_ hold951/X _09156_/B vssd1 vssd1 vccd1 vccd1 _09144_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09075_ hold2916/X _09106_/B _09074_/X _12948_/A vssd1 vssd1 vccd1 vccd1 _09075_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08026_ hold1686/X _08029_/B _08025_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _08026_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold730 hold730/A vssd1 vssd1 vccd1 vccd1 hold730/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 hold741/A vssd1 vssd1 vccd1 vccd1 hold741/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold752 hold752/A vssd1 vssd1 vccd1 vccd1 hold752/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 hold763/A vssd1 vssd1 vccd1 vccd1 hold763/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold774 hold774/A vssd1 vssd1 vccd1 vccd1 hold774/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 hold785/A vssd1 vssd1 vccd1 vccd1 hold785/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold796 hold796/A vssd1 vssd1 vccd1 vccd1 hold796/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09977_ hold2675/X _16483_/Q _10067_/C vssd1 vssd1 vccd1 vccd1 _09978_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_200_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2120 _14219_/X vssd1 vssd1 vccd1 vccd1 _17911_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2131 _17796_/Q vssd1 vssd1 vccd1 vccd1 hold2131/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2142 _14617_/X vssd1 vssd1 vccd1 vccd1 _18102_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08928_ hold495/X hold567/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold568/A sky130_fd_sc_hd__mux2_1
Xhold2153 _18224_/Q vssd1 vssd1 vccd1 vccd1 hold2153/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2164 _14221_/X vssd1 vssd1 vccd1 vccd1 _17912_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2175 _17947_/Q vssd1 vssd1 vccd1 vccd1 hold2175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1430 _15864_/Q vssd1 vssd1 vccd1 vccd1 hold1430/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2186 _14971_/X vssd1 vssd1 vccd1 vccd1 _18271_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1441 _13975_/X vssd1 vssd1 vccd1 vccd1 _17794_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1452 _08160_/X vssd1 vssd1 vccd1 vccd1 _08161_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2197 _15679_/Q vssd1 vssd1 vccd1 vccd1 hold2197/X sky130_fd_sc_hd__dlygate4sd3_1
X_08859_ _15434_/A hold262/X vssd1 vssd1 vccd1 vccd1 _16048_/D sky130_fd_sc_hd__and2_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1463 hold1540/X vssd1 vssd1 vccd1 vccd1 hold1541/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1474 _09292_/X vssd1 vssd1 vccd1 vccd1 _16256_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1485 _14195_/X vssd1 vssd1 vccd1 vccd1 _17900_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1496 _14813_/X vssd1 vssd1 vccd1 vccd1 _18196_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_58_wb_clk_i clkbuf_6_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18072_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _15706_/Q hold5714/X _13463_/S vssd1 vssd1 vccd1 vccd1 _11871_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10821_ _11109_/A _10821_/B vssd1 vssd1 vccd1 vccd1 _10821_/X sky130_fd_sc_hd__or2_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10752_ _11136_/A _10752_/B vssd1 vssd1 vccd1 vccd1 _10752_/X sky130_fd_sc_hd__or2_1
X_13540_ hold4731/X _13829_/B _13539_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13540_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13471_ hold5452/X _13874_/B _13470_/X _13684_/C1 vssd1 vssd1 vccd1 vccd1 _13471_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10683_ _11010_/A _10683_/B vssd1 vssd1 vccd1 vccd1 _10683_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12422_ _15434_/A _12422_/B vssd1 vssd1 vccd1 vccd1 _17304_/D sky130_fd_sc_hd__and2_1
X_15210_ hold1869/X _15221_/B _15209_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _15210_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16190_ _17881_/CLK _16190_/D vssd1 vssd1 vccd1 vccd1 _16190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15141_ _15195_/A _15157_/B vssd1 vssd1 vccd1 vccd1 _15141_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12353_ _17275_/Q _12353_/B _13409_/S vssd1 vssd1 vccd1 vccd1 _12353_/X sky130_fd_sc_hd__and3_1
XFILLER_0_90_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11304_ _12234_/A _11304_/B vssd1 vssd1 vccd1 vccd1 _11304_/X sky130_fd_sc_hd__or2_1
X_15072_ _15072_/A _15072_/B vssd1 vssd1 vccd1 vccd1 _18321_/D sky130_fd_sc_hd__and2_1
XFILLER_0_121_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12284_ hold1356/X _17252_/Q _12317_/C vssd1 vssd1 vccd1 vccd1 _12285_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14023_ hold2964/X _14038_/B _14022_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _14023_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11235_ _12093_/A _11235_/B vssd1 vssd1 vccd1 vccd1 _11235_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11166_ hold4309/X _11655_/A _11165_/X vssd1 vssd1 vccd1 vccd1 _11166_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10117_ hold3816/X _10619_/B _10116_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10117_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15974_ _17293_/CLK _15974_/D vssd1 vssd1 vccd1 vccd1 hold471/A sky130_fd_sc_hd__dfxtp_1
XTAP_5550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11097_ _11661_/A _11097_/B vssd1 vssd1 vccd1 vccd1 _11097_/X sky130_fd_sc_hd__or2_1
XTAP_5561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17713_ _17745_/CLK _17713_/D vssd1 vssd1 vccd1 vccd1 _17713_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10048_ _10603_/A _10048_/B vssd1 vssd1 vccd1 vccd1 _10048_/Y sky130_fd_sc_hd__nor2_1
X_14925_ hold2977/X _14952_/B _14924_/X _15202_/C1 vssd1 vssd1 vccd1 vccd1 _14925_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17644_ _17748_/CLK _17644_/D vssd1 vssd1 vccd1 vccd1 _17644_/Q sky130_fd_sc_hd__dfxtp_1
X_14856_ _15195_/A _14892_/B vssd1 vssd1 vccd1 vccd1 _14856_/X sky130_fd_sc_hd__or2_1
XFILLER_0_202_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13807_ _13819_/A _13807_/B vssd1 vssd1 vccd1 vccd1 _13807_/Y sky130_fd_sc_hd__nor2_1
X_17575_ _17735_/CLK _17575_/D vssd1 vssd1 vccd1 vccd1 _17575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14787_ hold1692/X _14774_/B _14786_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14787_/X
+ sky130_fd_sc_hd__o211a_1
X_11999_ hold2445/X hold4699/X _13796_/S vssd1 vssd1 vccd1 vccd1 _12000_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_202_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16526_ _18188_/CLK _16526_/D vssd1 vssd1 vccd1 vccd1 _16526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13738_ _13832_/A _13862_/B _13737_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _17699_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16457_ _18370_/CLK _16457_/D vssd1 vssd1 vccd1 vccd1 _16457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13669_ hold5496/X _13883_/B _13668_/X _13765_/C1 vssd1 vssd1 vccd1 vccd1 _13669_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15408_ hold743/X _15484_/A2 _09392_/D hold540/X vssd1 vssd1 vccd1 vccd1 _15408_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_182_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16388_ _18375_/CLK _16388_/D vssd1 vssd1 vccd1 vccd1 _16388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_435_wb_clk_i clkbuf_6_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17726_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18127_ _18215_/CLK _18127_/D vssd1 vssd1 vccd1 vccd1 _18127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15339_ hold465/X _09365_/B _15488_/A2 hold386/X _15338_/X vssd1 vssd1 vccd1 vccd1
+ _15342_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5707 _12349_/Y vssd1 vssd1 vccd1 vccd1 _17273_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5718 _12363_/Y vssd1 vssd1 vccd1 vccd1 _12364_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5729 _16336_/Q vssd1 vssd1 vccd1 vccd1 _13158_/A sky130_fd_sc_hd__dlygate4sd3_1
X_18058_ _18058_/CLK _18058_/D vssd1 vssd1 vccd1 vccd1 _18058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09900_ _09933_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09900_/X sky130_fd_sc_hd__or2_1
X_17009_ _17890_/CLK _17009_/D vssd1 vssd1 vccd1 vccd1 _17009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout506 _10604_/C vssd1 vssd1 vccd1 vccd1 _10628_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout517 _10649_/C vssd1 vssd1 vccd1 vccd1 _10640_/C sky130_fd_sc_hd__clkbuf_8
X_09831_ _11010_/A _09831_/B vssd1 vssd1 vccd1 vccd1 _09831_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout528 hold270/X vssd1 vssd1 vccd1 vccd1 hold271/A sky130_fd_sc_hd__clkbuf_1
Xfanout539 _08868_/X vssd1 vssd1 vccd1 vccd1 _12445_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_225_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09762_ _09954_/A _09762_/B vssd1 vssd1 vccd1 vccd1 _09762_/X sky130_fd_sc_hd__or2_1
XFILLER_0_225_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08713_ hold143/X hold174/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08714_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_207_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09693_ _11106_/A _09693_/B vssd1 vssd1 vccd1 vccd1 _09693_/X sky130_fd_sc_hd__or2_1
XFILLER_0_241_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08644_ _15314_/A _08644_/B vssd1 vssd1 vccd1 vccd1 _15944_/D sky130_fd_sc_hd__and2_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_234_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08575_ _15324_/A hold374/X vssd1 vssd1 vccd1 vccd1 _15911_/D sky130_fd_sc_hd__and2_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_176_wb_clk_i clkbuf_6_49_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18379_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_106_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09127_ hold1622/X _09177_/A2 _09126_/X _12855_/A vssd1 vssd1 vccd1 vccd1 _09127_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_105_wb_clk_i clkbuf_6_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17328_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_161_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09058_ hold495/X hold545/X _09060_/S vssd1 vssd1 vccd1 vccd1 hold546/A sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08009_ hold933/X _08045_/B vssd1 vssd1 vccd1 vccd1 _08009_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold560 hold560/A vssd1 vssd1 vccd1 vccd1 hold560/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold571 hold571/A vssd1 vssd1 vccd1 vccd1 hold571/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 hold582/A vssd1 vssd1 vccd1 vccd1 hold582/X sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ hold5339/X _11753_/B _11019_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11020_/X
+ sky130_fd_sc_hd__o211a_1
Xhold593 hold593/A vssd1 vssd1 vccd1 vccd1 hold593/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_217_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ hold3222/X _12970_/X _12971_/S vssd1 vssd1 vccd1 vccd1 _12971_/X sky130_fd_sc_hd__mux2_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1260 _16156_/Q vssd1 vssd1 vccd1 vccd1 hold1260/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ _15103_/A _14730_/B vssd1 vssd1 vccd1 vccd1 _14710_/X sky130_fd_sc_hd__or2_1
Xhold1271 _18092_/Q vssd1 vssd1 vccd1 vccd1 hold1271/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1282 _14355_/X vssd1 vssd1 vccd1 vccd1 _14356_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _12093_/A _11922_/B vssd1 vssd1 vccd1 vccd1 _11922_/X sky130_fd_sc_hd__or2_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15690_ _17209_/CLK hold956/X vssd1 vssd1 vccd1 vccd1 hold955/A sky130_fd_sc_hd__dfxtp_1
Xhold1293 _15672_/Q vssd1 vssd1 vccd1 vccd1 hold1293/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ hold2721/X _14664_/B _14640_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _14641_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_197_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _12255_/A _11853_/B vssd1 vssd1 vccd1 vccd1 _11853_/X sky130_fd_sc_hd__or2_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ hold4949/X _11186_/B _10803_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _10804_/X
+ sky130_fd_sc_hd__o211a_1
X_17360_ _17360_/CLK _17360_/D vssd1 vssd1 vccd1 vccd1 _17360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14572_ hold307/X _14573_/B vssd1 vssd1 vccd1 vccd1 _14572_/X sky130_fd_sc_hd__and2_2
X_11784_ hold3788/X _11667_/A _11783_/X vssd1 vssd1 vccd1 vccd1 _11784_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16311_ _18404_/CLK _16311_/D vssd1 vssd1 vccd1 vccd1 _16311_/Q sky130_fd_sc_hd__dfxtp_1
X_13523_ hold1172/X _17628_/Q _13811_/C vssd1 vssd1 vccd1 vccd1 _13524_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_165_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17291_ _17291_/CLK _17291_/D vssd1 vssd1 vccd1 vccd1 hold888/A sky130_fd_sc_hd__dfxtp_1
X_10735_ hold5372/X _11213_/B _10734_/X _14342_/A vssd1 vssd1 vccd1 vccd1 _10735_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16242_ _17690_/CLK _16242_/D vssd1 vssd1 vccd1 vccd1 _16242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10666_ hold3828/X _11144_/B _10665_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _10666_/X
+ sky130_fd_sc_hd__o211a_1
X_13454_ hold1704/X _17605_/Q _13871_/C vssd1 vssd1 vccd1 vccd1 _13455_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12405_ hold77/X hold701/X _12405_/S vssd1 vssd1 vccd1 vccd1 hold702/A sky130_fd_sc_hd__mux2_1
X_16173_ _18400_/CLK _16173_/D vssd1 vssd1 vccd1 vccd1 _16173_/Q sky130_fd_sc_hd__dfxtp_1
X_13385_ hold2343/X hold4442/X _13481_/S vssd1 vssd1 vccd1 vccd1 _13386_/B sky130_fd_sc_hd__mux2_1
X_10597_ _10651_/A _10597_/B vssd1 vssd1 vccd1 vccd1 _16689_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15124_ hold6061/X hold341/X _15123_/X _15066_/A vssd1 vssd1 vccd1 vccd1 hold342/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput109 hold4185/X vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_12
X_12336_ hold4433/X _12240_/A _12335_/X vssd1 vssd1 vccd1 vccd1 _12336_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_239_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15055_ hold597/X hold654/X _15071_/S vssd1 vssd1 vccd1 vccd1 hold655/A sky130_fd_sc_hd__mux2_1
X_12267_ _12267_/A _12267_/B vssd1 vssd1 vccd1 vccd1 _12267_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11218_ _11218_/A _11218_/B vssd1 vssd1 vccd1 vccd1 _11218_/Y sky130_fd_sc_hd__nor2_1
X_14006_ hold911/X _14042_/B vssd1 vssd1 vccd1 vccd1 _14006_/X sky130_fd_sc_hd__or2_1
XFILLER_0_208_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12198_ _12198_/A _12198_/B vssd1 vssd1 vccd1 vccd1 _12198_/X sky130_fd_sc_hd__or2_1
Xoutput80 _13193_/A vssd1 vssd1 vccd1 vccd1 output80/X sky130_fd_sc_hd__buf_6
Xoutput91 _13273_/A vssd1 vssd1 vccd1 vccd1 output91/X sky130_fd_sc_hd__buf_6
XFILLER_0_177_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11149_ _11158_/A _11149_/B vssd1 vssd1 vccd1 vccd1 _16873_/D sky130_fd_sc_hd__nor2_1
XTAP_6070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15957_ _16124_/CLK _15957_/D vssd1 vssd1 vccd1 vccd1 hold718/A sky130_fd_sc_hd__dfxtp_1
XTAP_5380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14908_ _15193_/A _14910_/B vssd1 vssd1 vccd1 vccd1 _14908_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15888_ _17318_/CLK _15888_/D vssd1 vssd1 vccd1 vccd1 hold813/A sky130_fd_sc_hd__dfxtp_1
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_1251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17627_ _17689_/CLK _17627_/D vssd1 vssd1 vccd1 vccd1 _17627_/Q sky130_fd_sc_hd__dfxtp_1
X_14839_ hold1750/X _14826_/B _14838_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14839_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08360_ _15529_/A hold2541/X hold115/X vssd1 vssd1 vccd1 vccd1 _08361_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17558_ _17686_/CLK _17558_/D vssd1 vssd1 vccd1 vccd1 _17558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_wb_clk_i clkbuf_6_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18457_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16509_ _18390_/CLK _16509_/D vssd1 vssd1 vccd1 vccd1 _16509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08291_ _14850_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08291_/X sky130_fd_sc_hd__or2_1
X_17489_ _17492_/CLK _17489_/D vssd1 vssd1 vccd1 vccd1 _17489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5504 _17682_/Q vssd1 vssd1 vccd1 vccd1 hold5504/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5515 _16836_/Q vssd1 vssd1 vccd1 vccd1 hold5515/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5526 _11245_/X vssd1 vssd1 vccd1 vccd1 _16905_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5537 _16945_/Q vssd1 vssd1 vccd1 vccd1 hold5537/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4803 _17222_/Q vssd1 vssd1 vccd1 vccd1 hold4803/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5548 _11716_/X vssd1 vssd1 vccd1 vccd1 _17062_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4814 _13429_/X vssd1 vssd1 vccd1 vccd1 _17596_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5559 _17131_/Q vssd1 vssd1 vccd1 vccd1 hold5559/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4825 _17223_/Q vssd1 vssd1 vccd1 vccd1 hold4825/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4836 _11824_/X vssd1 vssd1 vccd1 vccd1 _17098_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4847 _16358_/Q vssd1 vssd1 vccd1 vccd1 hold4847/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4858 _11995_/X vssd1 vssd1 vccd1 vccd1 _17155_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout303 _11106_/A vssd1 vssd1 vccd1 vccd1 _11067_/A sky130_fd_sc_hd__buf_4
Xhold4869 _16878_/Q vssd1 vssd1 vccd1 vccd1 hold4869/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout314 _10539_/A vssd1 vssd1 vccd1 vccd1 _10986_/A sky130_fd_sc_hd__clkbuf_4
Xfanout325 _10560_/A vssd1 vssd1 vccd1 vccd1 _10476_/A sky130_fd_sc_hd__buf_4
XFILLER_0_160_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout347 _09062_/S vssd1 vssd1 vccd1 vccd1 _09056_/S sky130_fd_sc_hd__buf_8
X_09814_ hold4768/X _10028_/B _09813_/X _15042_/A vssd1 vssd1 vccd1 vccd1 _09814_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout358 _08594_/S vssd1 vssd1 vccd1 vccd1 _08592_/S sky130_fd_sc_hd__buf_8
XFILLER_0_185_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout369 _15119_/B vssd1 vssd1 vccd1 vccd1 _15125_/B sky130_fd_sc_hd__buf_6
XFILLER_0_199_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_236_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09745_ hold4829/X _10031_/B _09744_/X _15146_/C1 vssd1 vssd1 vccd1 vccd1 _09745_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09676_ hold3228/X _10052_/B _09675_/X _15019_/C1 vssd1 vssd1 vccd1 vccd1 _09676_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ hold172/X _15936_/Q _08657_/S vssd1 vssd1 vccd1 vccd1 hold607/A sky130_fd_sc_hd__mux2_1
XFILLER_0_222_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08558_ hold169/X hold504/X _08592_/S vssd1 vssd1 vccd1 vccd1 hold505/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_357_wb_clk_i clkbuf_6_41_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17250_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_212_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08489_ hold2394/X _08488_/B _08488_/Y _13777_/C1 vssd1 vssd1 vccd1 vccd1 _08489_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10520_ hold1980/X hold5420/X _11213_/C vssd1 vssd1 vccd1 vccd1 _10521_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_162_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10451_ hold1845/X hold4620/X _10646_/C vssd1 vssd1 vccd1 vccd1 _10452_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_116_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13170_ _17572_/Q _17106_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13170_/X sky130_fd_sc_hd__mux2_1
X_10382_ hold2416/X _16618_/Q _10985_/S vssd1 vssd1 vccd1 vccd1 _10383_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12121_ hold5123/X _12217_/A2 _12120_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _12121_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12052_ hold5050/X _11771_/B _12051_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _12052_/X
+ sky130_fd_sc_hd__o211a_1
Xhold390 hold390/A vssd1 vssd1 vccd1 vccd1 hold390/X sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ hold3002/X _16825_/Q _11660_/S vssd1 vssd1 vccd1 vccd1 _11004_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_217_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_73_wb_clk_i clkbuf_6_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18010_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16860_ _18031_/CLK _16860_/D vssd1 vssd1 vccd1 vccd1 _16860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout870 _15219_/A vssd1 vssd1 vccd1 vccd1 _15165_/A sky130_fd_sc_hd__buf_12
X_15811_ _17426_/CLK _15811_/D vssd1 vssd1 vccd1 vccd1 _15811_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout881 hold2103/X vssd1 vssd1 vccd1 vccd1 hold2104/A sky130_fd_sc_hd__buf_6
X_16791_ _18056_/CLK _16791_/D vssd1 vssd1 vccd1 vccd1 _16791_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout892 hold945/X vssd1 vssd1 vccd1 vccd1 _15517_/A sky130_fd_sc_hd__buf_12
XFILLER_0_189_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15742_ _17745_/CLK _15742_/D vssd1 vssd1 vccd1 vccd1 _15742_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _12984_/A _12954_/B vssd1 vssd1 vccd1 vccd1 _17494_/D sky130_fd_sc_hd__and2_1
XFILLER_0_77_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1090 _14859_/X vssd1 vssd1 vccd1 vccd1 _18218_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _18461_/CLK _18461_/D vssd1 vssd1 vccd1 vccd1 _18461_/Q sky130_fd_sc_hd__dfxtp_2
X_11905_ hold4699/X _12308_/B _11904_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _11905_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15673_ _17741_/CLK _15673_/D vssd1 vssd1 vccd1 vccd1 _15673_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _12888_/A _12885_/B vssd1 vssd1 vccd1 vccd1 _17471_/D sky130_fd_sc_hd__and2_1
XFILLER_0_200_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17412_ _17754_/CLK _17412_/D vssd1 vssd1 vccd1 vccd1 _17412_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14624_ _14732_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14624_/X sky130_fd_sc_hd__or2_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18392_ _18392_/CLK _18392_/D vssd1 vssd1 vccd1 vccd1 _18392_/Q sky130_fd_sc_hd__dfxtp_1
X_11836_ hold4646/X _12356_/B _11835_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _11836_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _17345_/CLK hold21/X vssd1 vssd1 vccd1 vccd1 _17343_/Q sky130_fd_sc_hd__dfxtp_1
X_14555_ _18461_/Q _14555_/B _14555_/C vssd1 vssd1 vccd1 vccd1 _14573_/B sky130_fd_sc_hd__and3_4
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _12337_/A _11767_/B vssd1 vssd1 vccd1 vccd1 _11767_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_166_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13506_ _13734_/A _13506_/B vssd1 vssd1 vccd1 vccd1 _13506_/X sky130_fd_sc_hd__or2_1
X_10718_ hold2088/X hold3517/X _11219_/C vssd1 vssd1 vccd1 vccd1 _10719_/B sky130_fd_sc_hd__mux2_1
X_17274_ _17576_/CLK _17274_/D vssd1 vssd1 vccd1 vccd1 _17274_/Q sky130_fd_sc_hd__dfxtp_1
X_14486_ hold2501/X _14487_/B _14485_/Y _14552_/C1 vssd1 vssd1 vccd1 vccd1 _14486_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11698_ hold5589/X _12335_/B _11697_/X _14143_/C1 vssd1 vssd1 vccd1 vccd1 _11698_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16225_ _17456_/CLK _16225_/D vssd1 vssd1 vccd1 vccd1 _16225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13437_ _13734_/A _13437_/B vssd1 vssd1 vccd1 vccd1 _13437_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10649_ _16707_/Q _10649_/B _10649_/C vssd1 vssd1 vccd1 vccd1 _10649_/X sky130_fd_sc_hd__and3_1
XFILLER_0_180_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16156_ _17493_/CLK _16156_/D vssd1 vssd1 vccd1 vccd1 _16156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13368_ _13581_/A _13368_/B vssd1 vssd1 vccd1 vccd1 _13368_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15107_ _15541_/A hold341/X vssd1 vssd1 vccd1 vccd1 _15107_/Y sky130_fd_sc_hd__nand2_1
X_12319_ _13864_/A _12319_/B vssd1 vssd1 vccd1 vccd1 _12319_/Y sky130_fd_sc_hd__nor2_1
X_16087_ _17299_/CLK _16087_/D vssd1 vssd1 vccd1 vccd1 hold663/A sky130_fd_sc_hd__dfxtp_1
X_13299_ _13298_/X _16930_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13299_/X sky130_fd_sc_hd__mux2_1
Xhold3409 _10047_/Y vssd1 vssd1 vccd1 vccd1 _10048_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15038_ _15482_/A _15038_/B vssd1 vssd1 vccd1 vccd1 _18304_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2708 _14406_/X vssd1 vssd1 vccd1 vccd1 _18001_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2719 _16161_/Q vssd1 vssd1 vccd1 vccd1 hold2719/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07860_ hold1740/X _07865_/B _07859_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _07860_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07791_ hold361/X vssd1 vssd1 vccd1 vccd1 _14555_/C sky130_fd_sc_hd__inv_2
X_16989_ _17891_/CLK _16989_/D vssd1 vssd1 vccd1 vccd1 _16989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_223_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09530_ hold3182/X _13142_/A _10022_/C vssd1 vssd1 vccd1 vccd1 _09531_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_190_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_231_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09461_ _09463_/B _09463_/C _09463_/D vssd1 vssd1 vccd1 vccd1 _09461_/X sky130_fd_sc_hd__and3_1
XFILLER_0_91_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08412_ hold3076/X _08442_/A2 _08411_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08412_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09392_ _09392_/A _09392_/B _09392_/C _09392_/D vssd1 vssd1 vccd1 vccd1 _09392_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_148_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_450_wb_clk_i clkbuf_6_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17689_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08343_ _08389_/A _08343_/B vssd1 vssd1 vccd1 vccd1 _15803_/D sky130_fd_sc_hd__and2_1
XFILLER_0_15_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08274_ _15553_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08274_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6002 _16910_/Q vssd1 vssd1 vccd1 vccd1 hold6002/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6013 _17550_/Q vssd1 vssd1 vccd1 vccd1 hold6013/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6024 _17543_/Q vssd1 vssd1 vccd1 vccd1 hold6024/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6035 _17527_/Q vssd1 vssd1 vccd1 vccd1 hold6035/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6046 data_in[21] vssd1 vssd1 vccd1 vccd1 hold370/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5301 _17276_/Q vssd1 vssd1 vccd1 vccd1 hold5301/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5312 _11695_/X vssd1 vssd1 vccd1 vccd1 _17055_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold6057 _17856_/Q vssd1 vssd1 vccd1 vccd1 hold6057/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6068 _18337_/Q vssd1 vssd1 vccd1 vccd1 hold6068/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5323 _17252_/Q vssd1 vssd1 vccd1 vccd1 hold5323/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6079 _18274_/Q vssd1 vssd1 vccd1 vccd1 hold6079/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5334 _11599_/X vssd1 vssd1 vccd1 vccd1 _17023_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4600 _16577_/Q vssd1 vssd1 vccd1 vccd1 hold4600/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5345 _17169_/Q vssd1 vssd1 vccd1 vccd1 hold5345/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4611 _09931_/X vssd1 vssd1 vccd1 vccd1 _16467_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5356 _13561_/X vssd1 vssd1 vccd1 vccd1 _17640_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4622 _16463_/Q vssd1 vssd1 vccd1 vccd1 hold4622/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5367 _11017_/X vssd1 vssd1 vccd1 vccd1 _16829_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4633 _10552_/X vssd1 vssd1 vccd1 vccd1 _16674_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_6_46_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_46_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
Xhold5378 _17712_/Q vssd1 vssd1 vccd1 vccd1 hold5378/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5389 _10702_/X vssd1 vssd1 vccd1 vccd1 _16724_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4644 _16912_/Q vssd1 vssd1 vccd1 vccd1 hold4644/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3910 _13507_/X vssd1 vssd1 vccd1 vccd1 _17622_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4655 _11914_/X vssd1 vssd1 vccd1 vccd1 _17128_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3921 _16637_/Q vssd1 vssd1 vccd1 vccd1 hold3921/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4666 _16747_/Q vssd1 vssd1 vccd1 vccd1 hold4666/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4677 _16360_/Q vssd1 vssd1 vccd1 vccd1 hold4677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3932 _12229_/X vssd1 vssd1 vccd1 vccd1 _17233_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3943 _11089_/X vssd1 vssd1 vccd1 vccd1 _16853_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4688 _09661_/X vssd1 vssd1 vccd1 vccd1 _16377_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3954 _16602_/Q vssd1 vssd1 vccd1 vccd1 hold3954/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4699 _17157_/Q vssd1 vssd1 vccd1 vccd1 hold4699/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3965 _17454_/Q vssd1 vssd1 vccd1 vccd1 hold3965/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3976 _17144_/Q vssd1 vssd1 vccd1 vccd1 hold3976/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3987 _16576_/Q vssd1 vssd1 vccd1 vccd1 hold3987/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout155 _12986_/S vssd1 vssd1 vccd1 vccd1 _12929_/S sky130_fd_sc_hd__buf_6
Xhold3998 _10225_/X vssd1 vssd1 vccd1 vccd1 _16565_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout166 _13795_/A2 vssd1 vssd1 vccd1 vccd1 _13829_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_195_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout177 fanout210/X vssd1 vssd1 vccd1 vccd1 _11723_/B sky130_fd_sc_hd__clkbuf_4
Xfanout188 _12332_/B vssd1 vssd1 vccd1 vccd1 _12362_/B sky130_fd_sc_hd__buf_4
XFILLER_0_199_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout199 _11786_/B vssd1 vssd1 vccd1 vccd1 _11771_/B sky130_fd_sc_hd__clkbuf_8
X_07989_ hold1354/X _07991_/A2 _07988_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _07989_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09728_ hold654/X hold4801/X _11171_/C vssd1 vssd1 vccd1 vccd1 _09729_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_241_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09659_ _18290_/Q hold3245/X _10031_/C vssd1 vssd1 vccd1 vccd1 _09660_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_179_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_191_wb_clk_i clkbuf_6_52_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18349_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ hold2437/X _17401_/Q _12871_/S vssd1 vssd1 vccd1 vccd1 _12670_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11621_ hold2056/X _17031_/Q _11717_/C vssd1 vssd1 vccd1 vccd1 _11622_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_120_wb_clk_i clkbuf_6_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16026_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_194_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14340_ hold113/X _14502_/B vssd1 vssd1 vccd1 vccd1 _14340_/X sky130_fd_sc_hd__or2_4
XFILLER_0_231_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11552_ _17856_/Q _17008_/Q _11741_/C vssd1 vssd1 vccd1 vccd1 _11553_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_231_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10503_ _10986_/A _10503_/B vssd1 vssd1 vccd1 vccd1 _10503_/X sky130_fd_sc_hd__or2_1
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11483_ hold2090/X _16985_/Q _11783_/C vssd1 vssd1 vccd1 vccd1 _11484_/B sky130_fd_sc_hd__mux2_1
X_14271_ hold1360/X _14272_/B _14270_/Y _14526_/C1 vssd1 vssd1 vccd1 vccd1 _14271_/X
+ sky130_fd_sc_hd__o211a_1
X_16010_ _18417_/CLK _16010_/D vssd1 vssd1 vccd1 vccd1 hold574/A sky130_fd_sc_hd__dfxtp_1
X_10434_ _10470_/A _10434_/B vssd1 vssd1 vccd1 vccd1 _10434_/X sky130_fd_sc_hd__or2_1
X_13222_ _13222_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13222_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13153_ _13153_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13153_/X sky130_fd_sc_hd__and2_1
XFILLER_0_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10365_ _11091_/A _10365_/B vssd1 vssd1 vccd1 vccd1 _10365_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ hold1752/X _17192_/Q _13811_/C vssd1 vssd1 vccd1 vccd1 _12105_/B sky130_fd_sc_hd__mux2_1
Xhold5890 output96/X vssd1 vssd1 vccd1 vccd1 data_out[31] sky130_fd_sc_hd__buf_12
X_13084_ hold3442/X _13083_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13084_/X sky130_fd_sc_hd__mux2_2
X_17961_ _18208_/CLK _17961_/D vssd1 vssd1 vccd1 vccd1 _17961_/Q sky130_fd_sc_hd__dfxtp_1
X_10296_ _10524_/A _10296_/B vssd1 vssd1 vccd1 vccd1 _10296_/X sky130_fd_sc_hd__or2_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_218_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12035_ hold2509/X hold5345/X _12329_/C vssd1 vssd1 vccd1 vccd1 _12036_/B sky130_fd_sc_hd__mux2_1
X_16912_ _17867_/CLK _16912_/D vssd1 vssd1 vccd1 vccd1 _16912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17892_ _17892_/CLK _17892_/D vssd1 vssd1 vccd1 vccd1 _17892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16843_ _17976_/CLK _16843_/D vssd1 vssd1 vccd1 vccd1 _16843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16774_ _18041_/CLK _16774_/D vssd1 vssd1 vccd1 vccd1 _16774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_279_wb_clk_i clkbuf_6_50_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18234_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13986_ _15221_/A _13986_/B vssd1 vssd1 vccd1 vccd1 _13986_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_232_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15725_ _17742_/CLK _15725_/D vssd1 vssd1 vccd1 vccd1 _15725_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12937_ hold2382/X hold4467/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12937_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_208_wb_clk_i clkbuf_6_55_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18390_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18444_ _18445_/CLK _18444_/D vssd1 vssd1 vccd1 vccd1 _18444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15656_ _17899_/CLK _15656_/D vssd1 vssd1 vccd1 vccd1 _15656_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12868_ hold1186/X hold3120/X _12916_/S vssd1 vssd1 vccd1 vccd1 _12868_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_200_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ hold2824/X _14610_/B _14606_/Y _14807_/C1 vssd1 vssd1 vccd1 vccd1 _14607_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18375_ _18375_/CLK _18375_/D vssd1 vssd1 vccd1 vccd1 _18375_/Q sky130_fd_sc_hd__dfxtp_1
X_11819_ hold1506/X hold4762/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11820_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_145_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15587_ _17204_/CLK _15587_/D vssd1 vssd1 vccd1 vccd1 _15587_/Q sky130_fd_sc_hd__dfxtp_1
X_12799_ hold2747/X _17444_/Q _12811_/S vssd1 vssd1 vccd1 vccd1 _12799_/X sky130_fd_sc_hd__mux2_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17326_ _17345_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 _17326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14538_ hold2314/X _14537_/B _14537_/Y _13911_/A vssd1 vssd1 vccd1 vccd1 _14538_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17257_ _18447_/CLK _17257_/D vssd1 vssd1 vccd1 vccd1 _17257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14469_ _15203_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14469_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16208_ _17440_/CLK _16208_/D vssd1 vssd1 vccd1 vccd1 _16208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17188_ _17910_/CLK _17188_/D vssd1 vssd1 vccd1 vccd1 _17188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16139_ _16139_/CLK _16139_/D vssd1 vssd1 vccd1 vccd1 hold759/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3206 _16535_/Q vssd1 vssd1 vccd1 vccd1 hold3206/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3217 _09679_/X vssd1 vssd1 vccd1 vccd1 _16383_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08961_ hold169/X hold588/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold589/A sky130_fd_sc_hd__mux2_1
Xhold3228 _16414_/Q vssd1 vssd1 vccd1 vccd1 hold3228/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3239 _17496_/Q vssd1 vssd1 vccd1 vccd1 hold3239/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2505 _17889_/Q vssd1 vssd1 vccd1 vccd1 hold2505/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2516 _18111_/Q vssd1 vssd1 vccd1 vccd1 hold2516/X sky130_fd_sc_hd__dlygate4sd3_1
X_07912_ _14529_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07912_/X sky130_fd_sc_hd__or2_1
XFILLER_0_227_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2527 _14037_/X vssd1 vssd1 vccd1 vccd1 _17824_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08892_ hold163/X hold730/X _08930_/S vssd1 vssd1 vccd1 vccd1 hold731/A sky130_fd_sc_hd__mux2_1
Xhold2538 _07899_/X vssd1 vssd1 vccd1 vccd1 _15593_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1804 _15234_/X vssd1 vssd1 vccd1 vccd1 _18399_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2549 _14989_/X vssd1 vssd1 vccd1 vccd1 _18280_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1815 _18134_/Q vssd1 vssd1 vccd1 vccd1 hold1815/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1826 _07913_/X vssd1 vssd1 vccd1 vccd1 _15600_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07843_ _15521_/A _07871_/B vssd1 vssd1 vccd1 vccd1 _07843_/X sky130_fd_sc_hd__or2_1
XFILLER_0_236_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1837 _15640_/Q vssd1 vssd1 vccd1 vccd1 hold1837/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1848 _15188_/X vssd1 vssd1 vccd1 vccd1 _18376_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1859 _17816_/Q vssd1 vssd1 vccd1 vccd1 hold1859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09513_ _09987_/A _09513_/B vssd1 vssd1 vccd1 vccd1 _09513_/X sky130_fd_sc_hd__or2_1
XFILLER_0_56_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09444_ _09447_/B _09447_/C _09447_/D vssd1 vssd1 vccd1 vccd1 _09444_/X sky130_fd_sc_hd__and3_1
XFILLER_0_182_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09375_ _15480_/A _09375_/B _09375_/C _09375_/D vssd1 vssd1 vccd1 vccd1 _09375_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_136_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08326_ hold1218/X _08336_/A2 _08325_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08326_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08257_ hold1795/X _08262_/B _08256_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _08257_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_201_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08188_ hold2942/X _08209_/B _08187_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08188_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5120 _10984_/X vssd1 vssd1 vccd1 vccd1 _16818_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5131 _16788_/Q vssd1 vssd1 vccd1 vccd1 hold5131/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5142 _16568_/Q vssd1 vssd1 vccd1 vccd1 hold5142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5153 _11095_/X vssd1 vssd1 vccd1 vccd1 _16855_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5164 _10558_/X vssd1 vssd1 vccd1 vccd1 _16676_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5175 _17250_/Q vssd1 vssd1 vccd1 vccd1 hold5175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4430 _16913_/Q vssd1 vssd1 vccd1 vccd1 hold4430/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10150_ hold4461/X _10628_/B _10149_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10150_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5186 _09946_/X vssd1 vssd1 vccd1 vccd1 _16472_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4441 _17492_/Q vssd1 vssd1 vccd1 vccd1 hold4441/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4452 _16662_/Q vssd1 vssd1 vccd1 vccd1 hold4452/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5197 _17067_/Q vssd1 vssd1 vccd1 vccd1 hold5197/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4463 _16396_/Q vssd1 vssd1 vccd1 vccd1 hold4463/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4474 _17351_/Q vssd1 vssd1 vccd1 vccd1 hold4474/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4485 _09526_/X vssd1 vssd1 vccd1 vccd1 _16332_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3740 _16550_/Q vssd1 vssd1 vccd1 vccd1 hold3740/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10081_ hold3874/X _10571_/B _10080_/X _15228_/C1 vssd1 vssd1 vccd1 vccd1 _10081_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3751 _09517_/X vssd1 vssd1 vccd1 vccd1 _16329_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4496 _13851_/Y vssd1 vssd1 vccd1 vccd1 _13852_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3762 _10432_/X vssd1 vssd1 vccd1 vccd1 _16634_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3773 _16449_/Q vssd1 vssd1 vccd1 vccd1 hold3773/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3784 _12719_/X vssd1 vssd1 vccd1 vccd1 _12720_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3795 _16643_/Q vssd1 vssd1 vccd1 vccd1 hold3795/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13840_ _13873_/A _13840_/B vssd1 vssd1 vccd1 vccd1 _13840_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_138_1352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_372_wb_clk_i clkbuf_6_32_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17732_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_230_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13771_ hold5402/X _13871_/B _13770_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13771_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_230_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10983_ _11100_/A _10983_/B vssd1 vssd1 vccd1 vccd1 _10983_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_301_wb_clk_i clkbuf_6_38_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17865_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_230_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15510_ hold1477/X _15560_/A2 _15509_/X _12864_/A vssd1 vssd1 vccd1 vccd1 _15510_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12722_ hold3807/X _12721_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12723_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_97_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16490_ _18371_/CLK _16490_/D vssd1 vssd1 vccd1 vccd1 _16490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15441_ hold349/X _15441_/A2 _09386_/D hold281/X _15436_/X vssd1 vssd1 vccd1 vccd1
+ _15442_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12653_ hold3146/X _12652_/X _12851_/S vssd1 vssd1 vccd1 vccd1 _12654_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18160_ _18180_/CLK _18160_/D vssd1 vssd1 vccd1 vccd1 _18160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11604_ _12174_/A _11604_/B vssd1 vssd1 vccd1 vccd1 _11604_/X sky130_fd_sc_hd__or2_1
X_15372_ _15489_/A _15372_/B _15372_/C _15372_/D vssd1 vssd1 vccd1 vccd1 _15372_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12584_ hold3365/X _12583_/X _12923_/S vssd1 vssd1 vccd1 vccd1 _12585_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_37_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17111_ _17281_/CLK _17111_/D vssd1 vssd1 vccd1 vccd1 _17111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14323_ hold2408/X _14326_/B _14322_/Y _14388_/A vssd1 vssd1 vccd1 vccd1 _14323_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18091_ _18099_/CLK _18091_/D vssd1 vssd1 vccd1 vccd1 _18091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11535_ _11631_/A _11535_/B vssd1 vssd1 vccd1 vccd1 _11535_/X sky130_fd_sc_hd__or2_1
XFILLER_0_108_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17042_ _17858_/CLK _17042_/D vssd1 vssd1 vccd1 vccd1 _17042_/Q sky130_fd_sc_hd__dfxtp_1
X_14254_ _14988_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14254_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11466_ _11658_/A _11466_/B vssd1 vssd1 vccd1 vccd1 _11466_/X sky130_fd_sc_hd__or2_1
XFILLER_0_145_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13205_ _13204_/X hold4238/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13205_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10417_ hold3974/X _10631_/B _10416_/X _14691_/C1 vssd1 vssd1 vccd1 vccd1 _10417_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11397_ _12219_/A _11397_/B vssd1 vssd1 vccd1 vccd1 _11397_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14185_ hold1273/X _14202_/B _14184_/X _14346_/A vssd1 vssd1 vccd1 vccd1 _14185_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_221_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13136_ _13129_/X _13135_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17535_/D sky130_fd_sc_hd__o21a_1
X_10348_ hold4525/X _10628_/B _10347_/X _10564_/C1 vssd1 vssd1 vccd1 vccd1 _10348_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10279_ hold3259/X _10589_/B _10278_/X _14893_/C1 vssd1 vssd1 vccd1 vccd1 _10279_/X
+ sky130_fd_sc_hd__o211a_1
X_17944_ _17976_/CLK _17944_/D vssd1 vssd1 vccd1 vccd1 _17944_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _13066_/X hold5653/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13067_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12018_ _12093_/A _12018_/B vssd1 vssd1 vccd1 vccd1 _12018_/X sky130_fd_sc_hd__or2_1
X_17875_ _17904_/CLK _17875_/D vssd1 vssd1 vccd1 vccd1 _17875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16826_ _18066_/CLK _16826_/D vssd1 vssd1 vccd1 vccd1 _16826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_1365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16757_ _17960_/CLK _16757_/D vssd1 vssd1 vccd1 vccd1 _16757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13969_ hold2532/X _13995_/A2 _13968_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _13969_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_232_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15708_ _17614_/CLK _15708_/D vssd1 vssd1 vccd1 vccd1 hold622/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16688_ _18150_/CLK _16688_/D vssd1 vssd1 vccd1 vccd1 _16688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15639_ _17247_/CLK _15639_/D vssd1 vssd1 vccd1 vccd1 _15639_/Q sky130_fd_sc_hd__dfxtp_1
X_18427_ _18427_/CLK _18427_/D vssd1 vssd1 vccd1 vccd1 _18427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09160_ _15543_/A _09164_/B vssd1 vssd1 vccd1 vccd1 _09160_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_111_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18358_ _18388_/CLK _18358_/D vssd1 vssd1 vccd1 vccd1 _18358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08111_ _08111_/A _08111_/B vssd1 vssd1 vccd1 vccd1 _15694_/D sky130_fd_sc_hd__and2_1
X_17309_ _17309_/CLK _17309_/D vssd1 vssd1 vccd1 vccd1 hold460/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09091_ hold1446/X _09102_/B _09090_/X _14358_/A vssd1 vssd1 vccd1 vccd1 _09091_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18289_ _18321_/CLK _18289_/D vssd1 vssd1 vccd1 vccd1 _18289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08042_ hold1352/X _08033_/B _08041_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _08042_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold901 hold901/A vssd1 vssd1 vccd1 vccd1 hold901/X sky130_fd_sc_hd__buf_2
Xhold912 hold912/A vssd1 vssd1 vccd1 vccd1 hold912/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 hold923/A vssd1 vssd1 vccd1 vccd1 hold923/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold934 hold934/A vssd1 vssd1 vccd1 vccd1 hold934/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 hold945/A vssd1 vssd1 vccd1 vccd1 hold945/X sky130_fd_sc_hd__buf_12
Xhold956 hold956/A vssd1 vssd1 vccd1 vccd1 hold956/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 input68/X vssd1 vssd1 vccd1 vccd1 hold967/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold978 hold978/A vssd1 vssd1 vccd1 vccd1 hold978/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3003 _14462_/X vssd1 vssd1 vccd1 vccd1 _18028_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ _13094_/A _09987_/A _09992_/X vssd1 vssd1 vccd1 vccd1 _09993_/Y sky130_fd_sc_hd__a21oi_1
Xhold989 hold989/A vssd1 vssd1 vccd1 vccd1 input50/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3014 _17901_/Q vssd1 vssd1 vccd1 vccd1 hold3014/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3025 _17784_/Q vssd1 vssd1 vccd1 vccd1 hold3025/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3036 _14209_/X vssd1 vssd1 vccd1 vccd1 _17907_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2302 _18150_/Q vssd1 vssd1 vccd1 vccd1 hold2302/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3047 _15681_/Q vssd1 vssd1 vccd1 vccd1 hold3047/X sky130_fd_sc_hd__dlygate4sd3_1
X_08944_ _12416_/A _08944_/B vssd1 vssd1 vccd1 vccd1 _16089_/D sky130_fd_sc_hd__and2_1
Xhold3058 _09143_/X vssd1 vssd1 vccd1 vccd1 _16184_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2313 _13983_/X vssd1 vssd1 vccd1 vccd1 _17798_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3069 _14123_/X vssd1 vssd1 vccd1 vccd1 _17865_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2324 _17826_/Q vssd1 vssd1 vccd1 vccd1 hold2324/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2335 _15884_/Q vssd1 vssd1 vccd1 vccd1 hold2335/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2346 _15084_/X vssd1 vssd1 vccd1 vccd1 _18326_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1601 _07996_/X vssd1 vssd1 vccd1 vccd1 _15639_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2357 _15794_/Q vssd1 vssd1 vccd1 vccd1 hold2357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1612 _14191_/X vssd1 vssd1 vccd1 vccd1 _17898_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08875_ _15324_/A hold188/X vssd1 vssd1 vccd1 vccd1 _16055_/D sky130_fd_sc_hd__and2_1
Xhold1623 _09127_/X vssd1 vssd1 vccd1 vccd1 _16176_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2368 _08459_/X vssd1 vssd1 vccd1 vccd1 _15858_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2379 _13018_/X vssd1 vssd1 vccd1 vccd1 _17517_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1634 _08180_/X vssd1 vssd1 vccd1 vccd1 _15726_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1645 _16151_/Q vssd1 vssd1 vccd1 vccd1 hold1645/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07826_ _07826_/A _13048_/A vssd1 vssd1 vccd1 vccd1 _07826_/X sky130_fd_sc_hd__and2_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1656 _17786_/Q vssd1 vssd1 vccd1 vccd1 hold1656/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1667 _09209_/X vssd1 vssd1 vccd1 vccd1 _16216_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1678 _15602_/Q vssd1 vssd1 vccd1 vccd1 hold1678/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1689 _14454_/X vssd1 vssd1 vccd1 vccd1 _18024_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09427_ _07804_/A hold739/X _15274_/A _09426_/X vssd1 vssd1 vccd1 vccd1 hold740/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_212_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09358_ _09366_/A _09363_/B _09361_/C vssd1 vssd1 vccd1 vccd1 _09358_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08309_ _15533_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08309_/X sky130_fd_sc_hd__or2_1
XFILLER_0_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09289_ _15511_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09289_/X sky130_fd_sc_hd__or2_1
X_11320_ hold5086/X _11798_/B _11319_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _11320_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11251_ hold4901/X _11732_/B _11250_/X _13895_/A vssd1 vssd1 vccd1 vccd1 _11251_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10202_ hold2723/X _16558_/Q _10604_/C vssd1 vssd1 vccd1 vccd1 _10203_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_219_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11182_ _12331_/A _11182_/B vssd1 vssd1 vccd1 vccd1 _11182_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4260 _11154_/Y vssd1 vssd1 vccd1 vccd1 _11155_/B sky130_fd_sc_hd__dlygate4sd3_1
X_10133_ hold2287/X hold3206/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10134_/B sky130_fd_sc_hd__mux2_1
XTAP_6433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4271 _13812_/Y vssd1 vssd1 vccd1 vccd1 _13813_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15990_ _16129_/CLK _15990_/D vssd1 vssd1 vccd1 vccd1 hold300/A sky130_fd_sc_hd__dfxtp_1
XTAP_5710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4282 _11160_/Y vssd1 vssd1 vccd1 vccd1 _11161_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4293 _17581_/Q vssd1 vssd1 vccd1 vccd1 hold4293/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3570 _17433_/Q vssd1 vssd1 vccd1 vccd1 hold3570/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3581 _09913_/X vssd1 vssd1 vccd1 vccd1 _16461_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10064_ _16512_/Q _10568_/B _10571_/C vssd1 vssd1 vccd1 vccd1 _10064_/X sky130_fd_sc_hd__and3_1
X_14941_ hold1988/X _14952_/B _14940_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _14941_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3592 _11197_/Y vssd1 vssd1 vccd1 vccd1 _16889_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2880 _14815_/X vssd1 vssd1 vccd1 vccd1 _18197_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17660_ _17724_/CLK _17660_/D vssd1 vssd1 vccd1 vccd1 _17660_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14872_ _15103_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14872_/X sky130_fd_sc_hd__or2_1
Xhold2891 _18142_/Q vssd1 vssd1 vccd1 vccd1 hold2891/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16611_ _18224_/CLK _16611_/D vssd1 vssd1 vccd1 vccd1 _16611_/Q sky130_fd_sc_hd__dfxtp_1
X_13823_ _13823_/A _13862_/B _13862_/C vssd1 vssd1 vccd1 vccd1 _13823_/X sky130_fd_sc_hd__and3_1
XFILLER_0_173_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17591_ _17719_/CLK _17591_/D vssd1 vssd1 vccd1 vccd1 _17591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16542_ _18210_/CLK _16542_/D vssd1 vssd1 vccd1 vccd1 _16542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13754_ hold2822/X _17705_/Q _13880_/C vssd1 vssd1 vccd1 vccd1 _13755_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10966_ hold3310/X _10013_/B _10965_/X _14552_/C1 vssd1 vssd1 vccd1 vccd1 _10966_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12705_ _12786_/A _12705_/B vssd1 vssd1 vccd1 vccd1 _17411_/D sky130_fd_sc_hd__and2_1
XFILLER_0_85_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16473_ _18386_/CLK _16473_/D vssd1 vssd1 vccd1 vccd1 _16473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13685_ hold1795/X hold5504/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13686_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10897_ hold3933/X _11225_/B _10896_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _10897_/X
+ sky130_fd_sc_hd__o211a_1
X_18212_ _18212_/CLK _18212_/D vssd1 vssd1 vccd1 vccd1 _18212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15424_ _15482_/A _15424_/B vssd1 vssd1 vccd1 vccd1 _18418_/D sky130_fd_sc_hd__and2_1
XFILLER_0_156_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12636_ _12843_/A _12636_/B vssd1 vssd1 vccd1 vccd1 _17388_/D sky130_fd_sc_hd__and2_1
XFILLER_0_182_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18143_ _18205_/CLK _18143_/D vssd1 vssd1 vccd1 vccd1 _18143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15355_ hold660/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15355_/X sky130_fd_sc_hd__or2_1
XFILLER_0_170_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12567_ _12984_/A _12567_/B vssd1 vssd1 vccd1 vccd1 _17365_/D sky130_fd_sc_hd__and2_1
XFILLER_0_54_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14306_ hold951/X _14338_/B vssd1 vssd1 vccd1 vccd1 _14306_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18074_ _18106_/CLK hold928/X vssd1 vssd1 vccd1 vccd1 _18074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11518_ hold5269/X _12317_/B _11517_/X _14211_/C1 vssd1 vssd1 vccd1 vccd1 _11518_/X
+ sky130_fd_sc_hd__o211a_1
X_15286_ _17332_/Q _15486_/B1 _15485_/B1 hold145/X vssd1 vssd1 vccd1 vccd1 _15286_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12498_ _17342_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12498_/X sky130_fd_sc_hd__or2_1
Xhold208 hold208/A vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold219 input46/X vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__buf_1
X_17025_ _17873_/CLK _17025_/D vssd1 vssd1 vccd1 vccd1 _17025_/Q sky130_fd_sc_hd__dfxtp_1
X_14237_ hold2199/X _14268_/B _14236_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _14237_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11449_ hold5593/X _11744_/B _11448_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _11449_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14168_ hold911/X _14214_/B vssd1 vssd1 vccd1 vccd1 _14168_/X sky130_fd_sc_hd__or2_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _13199_/A1 _13117_/X _13118_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13119_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_221_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_294_wb_clk_i clkbuf_6_39_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18028_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ hold2147/X _14107_/A2 _14098_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _14099_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17927_ _18028_/CLK _17927_/D vssd1 vssd1 vccd1 vccd1 _17927_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_223_wb_clk_i clkbuf_6_61_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18215_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_147_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08660_ _12412_/A _08660_/B vssd1 vssd1 vccd1 vccd1 _15952_/D sky130_fd_sc_hd__and2_1
X_17858_ _17858_/CLK _17858_/D vssd1 vssd1 vccd1 vccd1 _17858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16809_ _18461_/CLK _16809_/D vssd1 vssd1 vccd1 vccd1 _16809_/Q sky130_fd_sc_hd__dfxtp_1
X_08591_ _15344_/A hold600/X vssd1 vssd1 vccd1 vccd1 _15919_/D sky130_fd_sc_hd__and2_1
XFILLER_0_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17789_ _17853_/CLK _17789_/D vssd1 vssd1 vccd1 vccd1 _17789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09212_ _15541_/A _09214_/B vssd1 vssd1 vccd1 vccd1 _09212_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_45_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09143_ hold3057/X _09177_/A2 _09142_/X _12873_/A vssd1 vssd1 vccd1 vccd1 _09143_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09074_ _15515_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09074_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08025_ _15539_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08025_/X sky130_fd_sc_hd__or2_1
Xhold720 hold720/A vssd1 vssd1 vccd1 vccd1 hold720/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold731 hold731/A vssd1 vssd1 vccd1 vccd1 hold731/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 hold742/A vssd1 vssd1 vccd1 vccd1 hold742/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 hold753/A vssd1 vssd1 vccd1 vccd1 hold753/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold764 hold764/A vssd1 vssd1 vccd1 vccd1 hold764/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold775 hold775/A vssd1 vssd1 vccd1 vccd1 hold775/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 hold786/A vssd1 vssd1 vccd1 vccd1 hold786/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold797 hold797/A vssd1 vssd1 vccd1 vccd1 hold797/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09976_ hold3686/X _10070_/B _09975_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _09976_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_228_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2110 _14422_/X vssd1 vssd1 vccd1 vccd1 _18009_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2121 _17821_/Q vssd1 vssd1 vccd1 vccd1 hold2121/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2132 _13979_/X vssd1 vssd1 vccd1 vccd1 _17796_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08927_ _09047_/A hold517/X vssd1 vssd1 vccd1 vccd1 _16081_/D sky130_fd_sc_hd__and2_1
XFILLER_0_200_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2143 _18259_/Q vssd1 vssd1 vccd1 vccd1 hold2143/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2154 _14871_/X vssd1 vssd1 vccd1 vccd1 _18224_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2165 _17918_/Q vssd1 vssd1 vccd1 vccd1 hold2165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1420 _17942_/Q vssd1 vssd1 vccd1 vccd1 hold1420/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2176 _14295_/X vssd1 vssd1 vccd1 vccd1 _17947_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1431 _08471_/X vssd1 vssd1 vccd1 vccd1 _15864_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1442 _15875_/Q vssd1 vssd1 vccd1 vccd1 hold1442/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08858_ hold82/X hold261/X _08858_/S vssd1 vssd1 vccd1 vccd1 hold262/A sky130_fd_sc_hd__mux2_1
XFILLER_0_157_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2187 _18283_/Q vssd1 vssd1 vccd1 vccd1 hold2187/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1453 _18444_/Q vssd1 vssd1 vccd1 vccd1 hold1453/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2198 _08079_/X vssd1 vssd1 vccd1 vccd1 _15679_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1464 hold1542/X vssd1 vssd1 vccd1 vccd1 hold1464/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1475 _18373_/Q vssd1 vssd1 vccd1 vccd1 hold1475/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07809_ _18459_/Q _07809_/B vssd1 vssd1 vccd1 vccd1 _07809_/X sky130_fd_sc_hd__or2_1
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1486 _17776_/Q vssd1 vssd1 vccd1 vccd1 hold1486/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1497 _15877_/Q vssd1 vssd1 vccd1 vccd1 hold1497/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08789_ hold495/X hold565/X _08793_/S vssd1 vssd1 vccd1 vccd1 hold566/A sky130_fd_sc_hd__mux2_1
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10820_ hold2813/X _16764_/Q _11204_/C vssd1 vssd1 vccd1 vccd1 _10821_/B sky130_fd_sc_hd__mux2_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_98_wb_clk_i clkbuf_6_22_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17309_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_149_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10751_ hold2139/X hold4799/X _11153_/C vssd1 vssd1 vccd1 vccd1 _10752_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13470_ _13788_/A _13470_/B vssd1 vssd1 vccd1 vccd1 _13470_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_wb_clk_i clkbuf_6_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17374_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10682_ hold3180/X hold4284/X _11171_/C vssd1 vssd1 vccd1 vccd1 _10683_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12421_ hold5/X hold349/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12422_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_180_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_5_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_168_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15140_ hold2641/X _15167_/B _15139_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _15140_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12352_ _13873_/A _12352_/B vssd1 vssd1 vccd1 vccd1 _12352_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_35_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11303_ _17773_/Q hold3788/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11304_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_239_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15071_ _15233_/A hold1388/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15072_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12283_ hold5275/X _13886_/B _12282_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _12283_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14022_ _15529_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14022_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11234_ hold1710/X hold5547/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11235_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_219_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11165_ _11165_/A _11165_/B _11654_/S vssd1 vssd1 vccd1 vccd1 _11165_/X sky130_fd_sc_hd__and3_1
XTAP_6241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4090 _11413_/X vssd1 vssd1 vccd1 vccd1 _16961_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10116_ _10524_/A _10116_/B vssd1 vssd1 vccd1 vccd1 _10116_/X sky130_fd_sc_hd__or2_1
XTAP_6274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15973_ _17301_/CLK _15973_/D vssd1 vssd1 vccd1 vccd1 hold638/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11096_ hold1536/X _16856_/Q _11660_/S vssd1 vssd1 vccd1 vccd1 _11097_/B sky130_fd_sc_hd__mux2_1
XTAP_6285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_234_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_216_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10047_ _13238_/A _09978_/A _10046_/X vssd1 vssd1 vccd1 vccd1 _10047_/Y sky130_fd_sc_hd__a21oi_1
X_14924_ _15193_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14924_/X sky130_fd_sc_hd__or2_1
X_17712_ _17744_/CLK _17712_/D vssd1 vssd1 vccd1 vccd1 _17712_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_188_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14855_ hold1244/X hold332/X _14854_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14855_/X
+ sky130_fd_sc_hd__o211a_1
X_17643_ _17702_/CLK _17643_/D vssd1 vssd1 vccd1 vccd1 _17643_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13806_ hold5720/X _13719_/A _13805_/X vssd1 vssd1 vccd1 vccd1 _13806_/Y sky130_fd_sc_hd__a21oi_1
X_17574_ _17606_/CLK _17574_/D vssd1 vssd1 vccd1 vccd1 _17574_/Q sky130_fd_sc_hd__dfxtp_1
X_14786_ _15233_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14786_/X sky130_fd_sc_hd__or2_1
X_11998_ hold5601/X _12305_/B _11997_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _11998_/X
+ sky130_fd_sc_hd__o211a_1
X_16525_ _18115_/CLK _16525_/D vssd1 vssd1 vccd1 vccd1 _16525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13737_ _13737_/A _13737_/B vssd1 vssd1 vccd1 vccd1 _13737_/X sky130_fd_sc_hd__or2_1
X_10949_ hold1843/X _16807_/Q _11144_/C vssd1 vssd1 vccd1 vccd1 _10950_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16456_ _18373_/CLK _16456_/D vssd1 vssd1 vccd1 vccd1 _16456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13668_ _13788_/A _13668_/B vssd1 vssd1 vccd1 vccd1 _13668_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15407_ _17316_/Q _15487_/A2 _15484_/B1 hold454/X _15406_/X vssd1 vssd1 vccd1 vccd1
+ _15412_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_128_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12619_ _18435_/Q _17384_/Q _12850_/S vssd1 vssd1 vccd1 vccd1 _12619_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16387_ _18390_/CLK _16387_/D vssd1 vssd1 vccd1 vccd1 _16387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13599_ _13599_/A _13599_/B vssd1 vssd1 vccd1 vccd1 _13599_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18126_ _18126_/CLK _18126_/D vssd1 vssd1 vccd1 vccd1 _18126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15338_ hold528/X _15484_/A2 _15441_/A2 hold357/X vssd1 vssd1 vccd1 vccd1 _15338_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5708 _17117_/Q vssd1 vssd1 vccd1 vccd1 hold5708/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5719 _12364_/Y vssd1 vssd1 vccd1 vccd1 _17278_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18057_ _18057_/CLK _18057_/D vssd1 vssd1 vccd1 vccd1 _18057_/Q sky130_fd_sc_hd__dfxtp_1
X_15269_ hold832/X _09365_/B _09392_/C hold527/X _15268_/X vssd1 vssd1 vccd1 vccd1
+ _15272_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_112_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17008_ _17888_/CLK _17008_/D vssd1 vssd1 vccd1 vccd1 _17008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_404_wb_clk_i clkbuf_6_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17886_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout507 _10604_/C vssd1 vssd1 vccd1 vccd1 _10646_/C sky130_fd_sc_hd__clkbuf_8
X_09830_ hold1648/X hold4839/X _11171_/C vssd1 vssd1 vccd1 vccd1 _09831_/B sky130_fd_sc_hd__mux2_1
Xfanout518 _09499_/Y vssd1 vssd1 vccd1 vccd1 _10649_/C sky130_fd_sc_hd__clkbuf_8
Xfanout529 _09206_/B vssd1 vssd1 vccd1 vccd1 _09230_/B sky130_fd_sc_hd__buf_4
XFILLER_0_226_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09761_ hold2137/X hold3650/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09762_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08712_ _15364_/A hold534/X vssd1 vssd1 vccd1 vccd1 _15977_/D sky130_fd_sc_hd__and2_1
XFILLER_0_207_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_225_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09692_ hold2668/X _16388_/Q _11201_/C vssd1 vssd1 vccd1 vccd1 _09693_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_240_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08643_ hold53/X hold793/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08644_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_222_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08574_ hold373/X _15911_/Q _08594_/S vssd1 vssd1 vccd1 vccd1 hold374/A sky130_fd_sc_hd__mux2_1
XFILLER_0_179_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09126_ _15509_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09126_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09057_ _09057_/A hold125/X vssd1 vssd1 vccd1 vccd1 _16145_/D sky130_fd_sc_hd__and2_1
XFILLER_0_142_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08008_ hold2445/X _08029_/B _08007_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _08008_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_145_wb_clk_i clkbuf_6_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18334_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_198_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold550 hold550/A vssd1 vssd1 vccd1 vccd1 hold550/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 hold561/A vssd1 vssd1 vccd1 vccd1 hold561/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold572 hold572/A vssd1 vssd1 vccd1 vccd1 hold572/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold583 hold583/A vssd1 vssd1 vccd1 vccd1 hold583/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold594 la_data_in[17] vssd1 vssd1 vccd1 vccd1 hold594/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09959_ hold2852/X _16477_/Q _10601_/C vssd1 vssd1 vccd1 vccd1 _09960_/B sky130_fd_sc_hd__mux2_1
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ hold1931/X _17501_/Q _12970_/S vssd1 vssd1 vccd1 vccd1 _12970_/X sky130_fd_sc_hd__mux2_1
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1250 hold6110/X vssd1 vssd1 vccd1 vccd1 hold640/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1261 _09083_/X vssd1 vssd1 vccd1 vccd1 _16156_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ hold2811/X hold5559/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11922_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_213_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1272 _14597_/X vssd1 vssd1 vccd1 vccd1 _18092_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1283 _18236_/Q vssd1 vssd1 vccd1 vccd1 hold1283/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1294 _08065_/X vssd1 vssd1 vccd1 vccd1 _15672_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _14980_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14640_/X sky130_fd_sc_hd__or2_1
XFILLER_0_169_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ hold2582/X hold4248/X _13463_/S vssd1 vssd1 vccd1 vccd1 _11853_/B sky130_fd_sc_hd__mux2_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10803_ _11091_/A _10803_/B vssd1 vssd1 vccd1 vccd1 _10803_/X sky130_fd_sc_hd__or2_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14571_ _14980_/A _14557_/Y hold2239/X _15218_/C1 vssd1 vssd1 vccd1 vccd1 _14571_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11783_ _17085_/Q _11786_/B _11783_/C vssd1 vssd1 vccd1 vccd1 _11783_/X sky130_fd_sc_hd__and3_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16310_ _18404_/CLK _16310_/D vssd1 vssd1 vccd1 vccd1 _16310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13522_ hold4715/X _13814_/B _13521_/X _08361_/A vssd1 vssd1 vccd1 vccd1 _13522_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17290_ _18405_/CLK _17290_/D vssd1 vssd1 vccd1 vccd1 hold274/A sky130_fd_sc_hd__dfxtp_1
X_10734_ _11103_/A _10734_/B vssd1 vssd1 vccd1 vccd1 _10734_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16241_ _17661_/CLK _16241_/D vssd1 vssd1 vccd1 vccd1 _16241_/Q sky130_fd_sc_hd__dfxtp_1
X_13453_ hold5046/X _13856_/B _13452_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13453_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10665_ _11049_/A _10665_/B vssd1 vssd1 vccd1 vccd1 _10665_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12404_ _12412_/A hold750/X vssd1 vssd1 vccd1 vccd1 _17295_/D sky130_fd_sc_hd__and2_1
XFILLER_0_152_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16172_ _17509_/CLK _16172_/D vssd1 vssd1 vccd1 vccd1 _16172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13384_ hold5101/X _13862_/B _13383_/X _13729_/C1 vssd1 vssd1 vccd1 vccd1 _13384_/X
+ sky130_fd_sc_hd__o211a_1
X_10596_ hold3499/X _10524_/A _10595_/X vssd1 vssd1 vccd1 vccd1 _10596_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15123_ hold289/X _15125_/B vssd1 vssd1 vccd1 vccd1 _15123_/X sky130_fd_sc_hd__or2_1
XFILLER_0_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12335_ _17269_/Q _12335_/B _12335_/C vssd1 vssd1 vccd1 vccd1 _12335_/X sky130_fd_sc_hd__and3_1
XFILLER_0_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15054_ _15054_/A hold834/X vssd1 vssd1 vccd1 vccd1 _18312_/D sky130_fd_sc_hd__and2_1
XFILLER_0_142_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12266_ hold2318/X _17246_/Q _12362_/C vssd1 vssd1 vccd1 vccd1 _12267_/B sky130_fd_sc_hd__mux2_1
X_14005_ hold2209/X _14040_/B _14004_/X _14143_/C1 vssd1 vssd1 vccd1 vccd1 _14005_/X
+ sky130_fd_sc_hd__o211a_1
X_11217_ hold4356/X _11121_/A _11216_/X vssd1 vssd1 vccd1 vccd1 _11217_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_235_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12197_ hold1945/X hold4825/X _12293_/C vssd1 vssd1 vccd1 vccd1 _12198_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_208_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput81 _13201_/A vssd1 vssd1 vccd1 vccd1 output81/X sky130_fd_sc_hd__buf_6
Xoutput92 _13281_/A vssd1 vssd1 vccd1 vccd1 output92/X sky130_fd_sc_hd__buf_6
XTAP_6060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11148_ hold4328/X _11136_/A _11147_/X vssd1 vssd1 vccd1 vccd1 _11148_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15956_ _16124_/CLK _15956_/D vssd1 vssd1 vccd1 vccd1 hold189/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11079_ _11658_/A _11079_/B vssd1 vssd1 vccd1 vccd1 _11079_/X sky130_fd_sc_hd__or2_1
XFILLER_0_235_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14907_ hold1017/X _14896_/Y _14906_/X _15404_/A vssd1 vssd1 vccd1 vccd1 _14907_/X
+ sky130_fd_sc_hd__o211a_1
X_15887_ _17324_/CLK _15887_/D vssd1 vssd1 vccd1 vccd1 hold764/A sky130_fd_sc_hd__dfxtp_1
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17626_ _17626_/CLK _17626_/D vssd1 vssd1 vccd1 vccd1 _17626_/Q sky130_fd_sc_hd__dfxtp_1
X_14838_ _15231_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14838_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17557_ _18229_/CLK _17557_/D vssd1 vssd1 vccd1 vccd1 _17557_/Q sky130_fd_sc_hd__dfxtp_1
X_14769_ hold1461/X _14772_/B _14768_/Y _14769_/C1 vssd1 vssd1 vccd1 vccd1 _14769_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16508_ _18389_/CLK _16508_/D vssd1 vssd1 vccd1 vccd1 _16508_/Q sky130_fd_sc_hd__dfxtp_1
X_17488_ _17492_/CLK _17488_/D vssd1 vssd1 vccd1 vccd1 _17488_/Q sky130_fd_sc_hd__dfxtp_1
X_08290_ hold2971/X _08323_/B _08289_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _08290_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16439_ _18352_/CLK _16439_/D vssd1 vssd1 vccd1 vccd1 _16439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5505 _16972_/Q vssd1 vssd1 vccd1 vccd1 hold5505/X sky130_fd_sc_hd__dlygate4sd3_1
X_18109_ _18172_/CLK _18109_/D vssd1 vssd1 vccd1 vccd1 _18109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5516 _10942_/X vssd1 vssd1 vccd1 vccd1 _16804_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5527 _17713_/Q vssd1 vssd1 vccd1 vccd1 hold5527/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5538 _11269_/X vssd1 vssd1 vccd1 vccd1 _16913_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5549 _16794_/Q vssd1 vssd1 vccd1 vccd1 hold5549/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4804 _12100_/X vssd1 vssd1 vccd1 vccd1 _17190_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_36_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_36_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
Xhold4815 _17211_/Q vssd1 vssd1 vccd1 vccd1 hold4815/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4826 _12103_/X vssd1 vssd1 vccd1 vccd1 _17191_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4837 _16781_/Q vssd1 vssd1 vccd1 vccd1 hold4837/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4848 _09508_/X vssd1 vssd1 vccd1 vccd1 _16326_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4859 _17256_/Q vssd1 vssd1 vccd1 vccd1 hold4859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout304 _09987_/A vssd1 vssd1 vccd1 vccd1 _09981_/A sky130_fd_sc_hd__buf_4
Xfanout315 _10539_/A vssd1 vssd1 vccd1 vccd1 _09957_/A sky130_fd_sc_hd__buf_4
XFILLER_0_10_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout326 wire337/X vssd1 vssd1 vccd1 vccd1 _10560_/A sky130_fd_sc_hd__clkbuf_4
X_09813_ _09933_/A _09813_/B vssd1 vssd1 vccd1 vccd1 _09813_/X sky130_fd_sc_hd__or2_1
Xfanout348 _08934_/X vssd1 vssd1 vccd1 vccd1 _08991_/S sky130_fd_sc_hd__buf_8
Xfanout359 _08544_/S vssd1 vssd1 vccd1 vccd1 _08594_/S sky130_fd_sc_hd__buf_8
XFILLER_0_96_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09744_ _09948_/A _09744_/B vssd1 vssd1 vccd1 vccd1 _09744_/X sky130_fd_sc_hd__or2_1
XFILLER_0_185_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09675_ _09957_/A _09675_/B vssd1 vssd1 vccd1 vccd1 _09675_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08626_ _15364_/A hold586/X vssd1 vssd1 vccd1 vccd1 _15935_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08557_ _15324_/A _08557_/B vssd1 vssd1 vccd1 vccd1 _15902_/D sky130_fd_sc_hd__and2_1
XFILLER_0_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08488_ _15221_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _08488_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_92_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_397_wb_clk_i clkbuf_6_36_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17889_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10450_ hold3610/X _10646_/B _10449_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _10450_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_326_wb_clk_i clkbuf_6_46_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17843_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09109_ hold1748/X _09106_/B _09108_/X _15284_/A vssd1 vssd1 vccd1 vccd1 _09109_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10381_ hold3593/X _10571_/B _10380_/X _14769_/C1 vssd1 vssd1 vccd1 vccd1 _10381_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12120_ _12216_/A _12120_/B vssd1 vssd1 vccd1 vccd1 _12120_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12051_ _12243_/A _12051_/B vssd1 vssd1 vccd1 vccd1 _12051_/X sky130_fd_sc_hd__or2_1
Xhold380 hold380/A vssd1 vssd1 vccd1 vccd1 hold380/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold391 hold391/A vssd1 vssd1 vccd1 vccd1 hold391/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11002_ hold5020/X _11195_/B _11001_/X _14526_/C1 vssd1 vssd1 vccd1 vccd1 _11002_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout860 hold5976/X vssd1 vssd1 vccd1 vccd1 _13056_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15810_ _17690_/CLK _15810_/D vssd1 vssd1 vccd1 vccd1 _15810_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout871 _07781_/Y vssd1 vssd1 vccd1 vccd1 _15219_/A sky130_fd_sc_hd__buf_12
XFILLER_0_176_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16790_ _17929_/CLK _16790_/D vssd1 vssd1 vccd1 vccd1 _16790_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout882 hold932/X vssd1 vssd1 vccd1 vccd1 hold933/A sky130_fd_sc_hd__buf_8
Xfanout893 hold945/X vssd1 vssd1 vccd1 vccd1 _14457_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_204_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15741_ _17744_/CLK _15741_/D vssd1 vssd1 vccd1 vccd1 _15741_/Q sky130_fd_sc_hd__dfxtp_1
X_12953_ hold3759/X _12952_/X _12986_/S vssd1 vssd1 vccd1 vccd1 _12953_/X sky130_fd_sc_hd__mux2_1
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1080 _08150_/X vssd1 vssd1 vccd1 vccd1 _08151_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1091 _15618_/Q vssd1 vssd1 vccd1 vccd1 hold1091/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ _13797_/A _11904_/B vssd1 vssd1 vccd1 vccd1 _11904_/X sky130_fd_sc_hd__or2_1
X_18460_ _18460_/CLK _18460_/D vssd1 vssd1 vccd1 vccd1 _18460_/Q sky130_fd_sc_hd__dfxtp_2
X_15672_ _17260_/CLK _15672_/D vssd1 vssd1 vccd1 vccd1 _15672_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_42_wb_clk_i clkbuf_6_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18427_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ hold3335/X _12883_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12884_/X sky130_fd_sc_hd__mux2_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ hold1724/X _14610_/B _14622_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14623_/X
+ sky130_fd_sc_hd__o211a_1
X_17411_ _17753_/CLK _17411_/D vssd1 vssd1 vccd1 vccd1 _17411_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18391_ _18391_/CLK _18391_/D vssd1 vssd1 vccd1 vccd1 _18391_/Q sky130_fd_sc_hd__dfxtp_1
X_11835_ _13482_/A _11835_/B vssd1 vssd1 vccd1 vccd1 _11835_/X sky130_fd_sc_hd__or2_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17347_/CLK hold36/X vssd1 vssd1 vccd1 vccd1 _17342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ hold6074/X _14537_/B hold550/X _13897_/A vssd1 vssd1 vccd1 vccd1 hold551/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ hold4337/X _11670_/A _11765_/X vssd1 vssd1 vccd1 vccd1 _11766_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13505_ hold963/X _17622_/Q _13766_/S vssd1 vssd1 vccd1 vccd1 _13506_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17273_ _17608_/CLK _17273_/D vssd1 vssd1 vccd1 vccd1 _17273_/Q sky130_fd_sc_hd__dfxtp_1
X_10717_ hold4135/X _11210_/B _10716_/X _14528_/C1 vssd1 vssd1 vccd1 vccd1 _10717_/X
+ sky130_fd_sc_hd__o211a_1
X_14485_ _15165_/A _14487_/B vssd1 vssd1 vccd1 vccd1 _14485_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_181_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11697_ _11697_/A _11697_/B vssd1 vssd1 vccd1 vccd1 _11697_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16224_ _17456_/CLK _16224_/D vssd1 vssd1 vccd1 vccd1 _16224_/Q sky130_fd_sc_hd__dfxtp_1
X_13436_ hold3076/X hold3763/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13437_/B sky130_fd_sc_hd__mux2_1
X_10648_ _11218_/A _10648_/B vssd1 vssd1 vccd1 vccd1 _10648_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_153_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16155_ _17493_/CLK _16155_/D vssd1 vssd1 vccd1 vccd1 _16155_/Q sky130_fd_sc_hd__dfxtp_1
X_13367_ hold1378/X hold3527/X _13868_/C vssd1 vssd1 vccd1 vccd1 _13368_/B sky130_fd_sc_hd__mux2_1
X_10579_ _10603_/A _10579_/B vssd1 vssd1 vccd1 vccd1 _16683_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_183_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15106_ hold6068/X hold340/X hold642/X _15404_/A vssd1 vssd1 vccd1 vccd1 hold643/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_239_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12318_ hold4315/X _12285_/A _12317_/X vssd1 vssd1 vccd1 vccd1 _12318_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16086_ _16086_/CLK _16086_/D vssd1 vssd1 vccd1 vccd1 hold716/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13298_ _17588_/Q _17122_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13298_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15037_ _15199_/A hold3099/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15038_/B sky130_fd_sc_hd__mux2_1
X_12249_ _13749_/A _12249_/B vssd1 vssd1 vccd1 vccd1 _12249_/X sky130_fd_sc_hd__or2_1
XFILLER_0_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2709 _18344_/Q vssd1 vssd1 vccd1 vccd1 hold2709/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07790_ hold353/X vssd1 vssd1 vccd1 vccd1 _14555_/B sky130_fd_sc_hd__inv_2
X_16988_ _17887_/CLK _16988_/D vssd1 vssd1 vccd1 vccd1 _16988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15939_ _18409_/CLK _15939_/D vssd1 vssd1 vccd1 vccd1 hold472/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09460_ _09463_/C _09463_/D _09463_/B vssd1 vssd1 vccd1 vccd1 _09462_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_204_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08411_ _15525_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08411_/X sky130_fd_sc_hd__or2_1
X_17609_ _17737_/CLK _17609_/D vssd1 vssd1 vccd1 vccd1 _17609_/Q sky130_fd_sc_hd__dfxtp_1
X_09391_ _16283_/Q _09342_/B _09342_/Y _09390_/X _12412_/A vssd1 vssd1 vccd1 vccd1
+ _09391_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_47_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08342_ hold915/X hold1669/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08343_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08273_ hold1327/X _08268_/B _08272_/X _12738_/A vssd1 vssd1 vccd1 vccd1 _08273_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6003 _16905_/Q vssd1 vssd1 vccd1 vccd1 hold6003/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6014 _17538_/Q vssd1 vssd1 vccd1 vccd1 hold6014/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6025 _17544_/Q vssd1 vssd1 vccd1 vccd1 hold6025/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6036 _17526_/Q vssd1 vssd1 vccd1 vccd1 hold6036/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6047 data_in[29] vssd1 vssd1 vccd1 vccd1 hold492/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5302 _12262_/X vssd1 vssd1 vccd1 vccd1 _17244_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6058 _17515_/Q vssd1 vssd1 vccd1 vccd1 hold6058/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5313 _16991_/Q vssd1 vssd1 vccd1 vccd1 hold5313/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6069 _16203_/Q vssd1 vssd1 vccd1 vccd1 hold6069/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5324 _12190_/X vssd1 vssd1 vccd1 vccd1 _17220_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5335 _16793_/Q vssd1 vssd1 vccd1 vccd1 hold5335/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4601 _10165_/X vssd1 vssd1 vccd1 vccd1 _16545_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5346 _11941_/X vssd1 vssd1 vccd1 vccd1 _17137_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5357 _17605_/Q vssd1 vssd1 vccd1 vccd1 hold5357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4612 _17727_/Q vssd1 vssd1 vccd1 vccd1 hold4612/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4623 _09823_/X vssd1 vssd1 vccd1 vccd1 _16431_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5368 _17001_/Q vssd1 vssd1 vccd1 vccd1 hold5368/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4634 _16709_/Q vssd1 vssd1 vccd1 vccd1 hold4634/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5379 _13681_/X vssd1 vssd1 vccd1 vccd1 _17680_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3900 _10219_/X vssd1 vssd1 vccd1 vccd1 _16563_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4645 _11745_/Y vssd1 vssd1 vccd1 vccd1 _11746_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3911 _16391_/Q vssd1 vssd1 vccd1 vccd1 hold3911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4656 _16401_/Q vssd1 vssd1 vccd1 vccd1 hold4656/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3922 _10345_/X vssd1 vssd1 vccd1 vccd1 _16605_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4667 _10675_/X vssd1 vssd1 vccd1 vccd1 _16715_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4678 _09514_/X vssd1 vssd1 vccd1 vccd1 _16328_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3933 _16821_/Q vssd1 vssd1 vccd1 vccd1 hold3933/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3944 _16510_/Q vssd1 vssd1 vccd1 vccd1 hold3944/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4689 _17662_/Q vssd1 vssd1 vccd1 vccd1 hold4689/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3955 _10240_/X vssd1 vssd1 vccd1 vccd1 _16570_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3966 _12833_/X vssd1 vssd1 vccd1 vccd1 _12834_/B sky130_fd_sc_hd__dlygate4sd3_1
Xfanout156 _12986_/S vssd1 vssd1 vccd1 vccd1 _13001_/S sky130_fd_sc_hd__buf_6
Xhold3977 _11866_/X vssd1 vssd1 vccd1 vccd1 _17112_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3988 _10162_/X vssd1 vssd1 vccd1 vccd1 _16544_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout167 _13795_/A2 vssd1 vssd1 vccd1 vccd1 _13862_/B sky130_fd_sc_hd__buf_4
XFILLER_0_226_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3999 _16570_/Q vssd1 vssd1 vccd1 vccd1 hold3999/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout178 _11741_/B vssd1 vssd1 vccd1 vccd1 _12317_/B sky130_fd_sc_hd__buf_4
Xfanout189 _12332_/B vssd1 vssd1 vccd1 vccd1 _12350_/B sky130_fd_sc_hd__buf_4
X_07988_ _15557_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07988_/X sky130_fd_sc_hd__or2_1
XFILLER_0_199_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09727_ hold4557/X _10004_/B _09726_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _09727_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09658_ hold4919/X _10070_/B _09657_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _09658_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ hold147/X hold560/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08610_/B sky130_fd_sc_hd__mux2_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09589_ hold3270/X _10568_/B _09588_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _09589_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11620_ hold5567/X _12305_/B _11619_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _11620_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11551_ hold4087/X _11741_/B _11550_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _11551_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10502_ hold1244/X _16658_/Q _11183_/C vssd1 vssd1 vccd1 vccd1 _10503_/B sky130_fd_sc_hd__mux2_1
X_14270_ _15219_/A _14272_/B vssd1 vssd1 vccd1 vccd1 _14270_/Y sky130_fd_sc_hd__nand2_1
X_11482_ hold4875/X _11798_/B _11481_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _11482_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_160_wb_clk_i clkbuf_6_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17295_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_135_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13221_ _13220_/X hold3515/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13221_/X sky130_fd_sc_hd__mux2_1
X_10433_ _18193_/Q _16635_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10434_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_208_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13152_ _13145_/X _13151_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17537_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_27_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10364_ hold1919/X _16612_/Q _10985_/S vssd1 vssd1 vccd1 vccd1 _10365_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12103_ hold4825/X _12293_/B _12102_/X _12103_/C1 vssd1 vssd1 vccd1 vccd1 _12103_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5880 output80/X vssd1 vssd1 vccd1 vccd1 data_out[17] sky130_fd_sc_hd__buf_12
XFILLER_0_209_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17960_ _17960_/CLK _17960_/D vssd1 vssd1 vccd1 vccd1 _17960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _13082_/X _16903_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13083_/X sky130_fd_sc_hd__mux2_1
Xhold5891 hold6030/X vssd1 vssd1 vccd1 vccd1 _13297_/A sky130_fd_sc_hd__buf_1
X_10295_ hold2049/X hold3995/X _10595_/C vssd1 vssd1 vccd1 vccd1 _10296_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12034_ hold4791/X _12353_/B _12033_/X _12289_/C1 vssd1 vssd1 vccd1 vccd1 _12034_/X
+ sky130_fd_sc_hd__o211a_1
X_16911_ _17825_/CLK _16911_/D vssd1 vssd1 vccd1 vccd1 _16911_/Q sky130_fd_sc_hd__dfxtp_1
X_17891_ _17891_/CLK _17891_/D vssd1 vssd1 vccd1 vccd1 _17891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16842_ _17981_/CLK _16842_/D vssd1 vssd1 vccd1 vccd1 _16842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout690 _12987_/A vssd1 vssd1 vccd1 vccd1 _12948_/A sky130_fd_sc_hd__buf_4
XFILLER_0_189_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16773_ _17976_/CLK _16773_/D vssd1 vssd1 vccd1 vccd1 _16773_/Q sky130_fd_sc_hd__dfxtp_1
X_13985_ hold2455/X _13986_/B _13984_/Y _13935_/A vssd1 vssd1 vccd1 vccd1 _13985_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12936_ _12948_/A _12936_/B vssd1 vssd1 vccd1 vccd1 _17488_/D sky130_fd_sc_hd__and2_1
X_15724_ _17730_/CLK _15724_/D vssd1 vssd1 vccd1 vccd1 _15724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18443_ _18443_/CLK _18443_/D vssd1 vssd1 vccd1 vccd1 _18443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15655_ _17229_/CLK _15655_/D vssd1 vssd1 vccd1 vccd1 _15655_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ _12888_/A _12867_/B vssd1 vssd1 vccd1 vccd1 _17465_/D sky130_fd_sc_hd__and2_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14606_ _15215_/A _14610_/B vssd1 vssd1 vccd1 vccd1 _14606_/Y sky130_fd_sc_hd__nand2_1
X_11818_ hold4805/X _13811_/B _11817_/X _08363_/A vssd1 vssd1 vccd1 vccd1 _11818_/X
+ sky130_fd_sc_hd__o211a_1
X_18374_ _18374_/CLK _18374_/D vssd1 vssd1 vccd1 vccd1 _18374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15586_ _17590_/CLK _15586_/D vssd1 vssd1 vccd1 vccd1 _15586_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_248_wb_clk_i clkbuf_6_59_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18154_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12798_ _12798_/A _12798_/B vssd1 vssd1 vccd1 vccd1 _17442_/D sky130_fd_sc_hd__and2_1
XFILLER_0_12_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _17325_/CLK hold75/X vssd1 vssd1 vccd1 vccd1 _17325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14537_ _15163_/A _14537_/B vssd1 vssd1 vccd1 vccd1 _14537_/Y sky130_fd_sc_hd__nand2_1
X_11749_ _12301_/A _11749_/B vssd1 vssd1 vccd1 vccd1 _11749_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_84_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14468_ hold2962/X _14481_/B _14467_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _14468_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17256_ _18443_/CLK _17256_/D vssd1 vssd1 vccd1 vccd1 _17256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13419_ _13722_/A _13419_/B vssd1 vssd1 vccd1 vccd1 _13419_/X sky130_fd_sc_hd__or2_1
X_16207_ _17446_/CLK hold983/X vssd1 vssd1 vccd1 vccd1 hold982/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17187_ _17187_/CLK _17187_/D vssd1 vssd1 vccd1 vccd1 _17187_/Q sky130_fd_sc_hd__dfxtp_1
X_14399_ hold911/X _14445_/B vssd1 vssd1 vccd1 vccd1 _14399_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16138_ _17339_/CLK _16138_/D vssd1 vssd1 vccd1 vccd1 hold571/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3207 _10614_/Y vssd1 vssd1 vccd1 vccd1 _10615_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08960_ _15491_/A hold250/X vssd1 vssd1 vccd1 vccd1 _16097_/D sky130_fd_sc_hd__and2_1
X_16069_ _18408_/CLK _16069_/D vssd1 vssd1 vccd1 vccd1 hold724/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3218 _16367_/Q vssd1 vssd1 vccd1 vccd1 hold3218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3229 _09676_/X vssd1 vssd1 vccd1 vccd1 _16382_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07911_ hold2703/X _07918_/B _07910_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _07911_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2506 _14173_/X vssd1 vssd1 vccd1 vccd1 _17889_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2517 _14637_/X vssd1 vssd1 vccd1 vccd1 _18111_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08891_ _15344_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _16063_/D sky130_fd_sc_hd__and2_1
Xhold2528 _18203_/Q vssd1 vssd1 vccd1 vccd1 hold2528/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2539 _15571_/Q vssd1 vssd1 vccd1 vccd1 hold2539/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1805 _18395_/Q vssd1 vssd1 vccd1 vccd1 hold1805/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1816 _14685_/X vssd1 vssd1 vccd1 vccd1 _18134_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07842_ hold1025/X _07865_/B _07841_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _07842_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1827 _18284_/Q vssd1 vssd1 vccd1 vccd1 hold1827/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1838 _07998_/X vssd1 vssd1 vccd1 vccd1 _15640_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1849 _17861_/Q vssd1 vssd1 vccd1 vccd1 hold1849/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09512_ hold1017/X _13094_/A _09992_/C vssd1 vssd1 vccd1 vccd1 _09513_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09443_ _09447_/C _09447_/D _09442_/Y vssd1 vssd1 vccd1 vccd1 _09443_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_231_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09374_ hold593/X _09365_/B _09362_/D hold344/X _09373_/X vssd1 vssd1 vccd1 vccd1
+ _09375_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_192_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08325_ _15549_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08325_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08256_ _14529_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08256_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08187_ _14461_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08187_/X sky130_fd_sc_hd__or2_1
Xhold5110 _10963_/X vssd1 vssd1 vccd1 vccd1 _16811_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5121 _17151_/Q vssd1 vssd1 vccd1 vccd1 hold5121/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5132 _10798_/X vssd1 vssd1 vccd1 vccd1 _16756_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5143 _10138_/X vssd1 vssd1 vccd1 vccd1 _16536_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5154 _16829_/Q vssd1 vssd1 vccd1 vccd1 hold5154/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4420 _11733_/Y vssd1 vssd1 vccd1 vccd1 _11734_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5165 _16818_/Q vssd1 vssd1 vccd1 vccd1 hold5165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5176 _12184_/X vssd1 vssd1 vccd1 vccd1 _17218_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4431 _11748_/Y vssd1 vssd1 vccd1 vccd1 _11749_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5187 _16805_/Q vssd1 vssd1 vccd1 vccd1 hold5187/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4442 _17582_/Q vssd1 vssd1 vccd1 vccd1 hold4442/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4453 _10420_/X vssd1 vssd1 vccd1 vccd1 _16630_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5198 _11635_/X vssd1 vssd1 vccd1 vccd1 _17035_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4464 _09622_/X vssd1 vssd1 vccd1 vccd1 _16364_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4475 _16558_/Q vssd1 vssd1 vccd1 vccd1 hold4475/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3730 _16688_/Q vssd1 vssd1 vccd1 vccd1 hold3730/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3741 _10084_/X vssd1 vssd1 vccd1 vccd1 _16518_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10080_ _10560_/A _10080_/B vssd1 vssd1 vccd1 vccd1 _10080_/X sky130_fd_sc_hd__or2_1
Xhold4486 _17363_/Q vssd1 vssd1 vccd1 vccd1 hold4486/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3752 _17444_/Q vssd1 vssd1 vccd1 vccd1 hold3752/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4497 _13852_/Y vssd1 vssd1 vccd1 vccd1 _17737_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3763 _17599_/Q vssd1 vssd1 vccd1 vccd1 hold3763/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3774 _09781_/X vssd1 vssd1 vccd1 vccd1 _16417_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3785 _16639_/Q vssd1 vssd1 vccd1 vccd1 hold3785/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3796 _10363_/X vssd1 vssd1 vccd1 vccd1 _16611_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_230_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_230_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13770_ _13776_/A _13770_/B vssd1 vssd1 vccd1 vccd1 _13770_/X sky130_fd_sc_hd__or2_1
X_10982_ hold1067/X _16818_/Q _11753_/C vssd1 vssd1 vccd1 vccd1 _10983_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12721_ hold2552/X hold3400/X _12766_/S vssd1 vssd1 vccd1 vccd1 _12721_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15440_ hold523/X _09365_/B _09362_/D hold755/X _15438_/X vssd1 vssd1 vccd1 vccd1
+ _15442_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_84_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12652_ hold2155/X hold3143/X _12850_/S vssd1 vssd1 vccd1 vccd1 _12652_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_341_wb_clk_i clkbuf_6_43_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17735_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11603_ hold1570/X hold4941/X _12173_/S vssd1 vssd1 vccd1 vccd1 _11604_/B sky130_fd_sc_hd__mux2_1
X_15371_ _16301_/Q _15477_/A2 _15487_/B1 hold754/X _15370_/X vssd1 vssd1 vccd1 vccd1
+ _15372_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_38_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12583_ hold3029/X hold3131/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12583_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14322_ _15163_/A _14326_/B vssd1 vssd1 vccd1 vccd1 _14322_/Y sky130_fd_sc_hd__nand2_1
X_17110_ _17272_/CLK _17110_/D vssd1 vssd1 vccd1 vccd1 _17110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18090_ _18220_/CLK _18090_/D vssd1 vssd1 vccd1 vccd1 _18090_/Q sky130_fd_sc_hd__dfxtp_1
X_11534_ hold2871/X _17002_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _11535_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_52_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17041_ _17889_/CLK _17041_/D vssd1 vssd1 vccd1 vccd1 _17041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14253_ hold2952/X _14272_/B _14252_/X _14528_/C1 vssd1 vssd1 vccd1 vccd1 _14253_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11465_ hold1409/X hold5261/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11466_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13204_ hold4318/X _13203_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13204_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10416_ _10554_/A _10416_/B vssd1 vssd1 vccd1 vccd1 _10416_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14184_ _15203_/A _14204_/B vssd1 vssd1 vccd1 vccd1 _14184_/X sky130_fd_sc_hd__or2_1
X_11396_ hold1457/X _16956_/Q _11741_/C vssd1 vssd1 vccd1 vccd1 _11397_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13135_ _13199_/A1 _13133_/X _13134_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13135_/X
+ sky130_fd_sc_hd__o211a_1
X_10347_ _10515_/A _10347_/B vssd1 vssd1 vccd1 vccd1 _10347_/X sky130_fd_sc_hd__or2_1
XFILLER_0_221_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17943_ _18073_/CLK hold584/X vssd1 vssd1 vccd1 vccd1 hold583/A sky130_fd_sc_hd__dfxtp_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _17559_/Q _17093_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13066_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_221_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10278_ _10470_/A _10278_/B vssd1 vssd1 vccd1 vccd1 _10278_/X sky130_fd_sc_hd__or2_1
X_12017_ hold2396/X _17163_/Q _12305_/C vssd1 vssd1 vccd1 vccd1 _12018_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17874_ _17874_/CLK _17874_/D vssd1 vssd1 vccd1 vccd1 _17874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16825_ _18060_/CLK _16825_/D vssd1 vssd1 vccd1 vccd1 _16825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16756_ _18023_/CLK _16756_/D vssd1 vssd1 vccd1 vccd1 _16756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13968_ _15529_/A _13994_/B vssd1 vssd1 vccd1 vccd1 _13968_/X sky130_fd_sc_hd__or2_1
XFILLER_0_159_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_429_wb_clk_i clkbuf_6_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17709_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_216_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15707_ _17741_/CLK _15707_/D vssd1 vssd1 vccd1 vccd1 hold535/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12919_ hold1334/X hold3314/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12919_/X sky130_fd_sc_hd__mux2_1
X_16687_ _18213_/CLK _16687_/D vssd1 vssd1 vccd1 vccd1 _16687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13899_ _13901_/A _13899_/B vssd1 vssd1 vccd1 vccd1 _17757_/D sky130_fd_sc_hd__and2_1
XFILLER_0_186_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_236_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18426_ _18428_/CLK _18426_/D vssd1 vssd1 vccd1 vccd1 _18426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15638_ _17266_/CLK _15638_/D vssd1 vssd1 vccd1 vccd1 _15638_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18357_ _18357_/CLK _18357_/D vssd1 vssd1 vccd1 vccd1 _18357_/Q sky130_fd_sc_hd__dfxtp_1
X_15569_ _17269_/CLK _15569_/D vssd1 vssd1 vccd1 vccd1 _15569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08110_ _14850_/A hold2525/X hold108/X vssd1 vssd1 vccd1 vccd1 _08111_/B sky130_fd_sc_hd__mux2_1
X_17308_ _17328_/CLK _17308_/D vssd1 vssd1 vccd1 vccd1 hold653/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09090_ _14596_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _09090_/X sky130_fd_sc_hd__or2_1
X_18288_ _18352_/CLK _18288_/D vssd1 vssd1 vccd1 vccd1 _18288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08041_ _14960_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08041_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17239_ _17271_/CLK _17239_/D vssd1 vssd1 vccd1 vccd1 _17239_/Q sky130_fd_sc_hd__dfxtp_1
Xhold902 hold902/A vssd1 vssd1 vccd1 vccd1 hold902/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold913 hold913/A vssd1 vssd1 vccd1 vccd1 hold913/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold924 hold924/A vssd1 vssd1 vccd1 vccd1 hold924/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold935 hold935/A vssd1 vssd1 vccd1 vccd1 hold935/X sky130_fd_sc_hd__clkbuf_4
Xhold946 hold946/A vssd1 vssd1 vccd1 vccd1 hold946/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 hold957/A vssd1 vssd1 vccd1 vccd1 hold957/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 hold968/A vssd1 vssd1 vccd1 vccd1 hold968/X sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ _16488_/Q _09992_/B _09992_/C vssd1 vssd1 vccd1 vccd1 _09992_/X sky130_fd_sc_hd__and3_1
XFILLER_0_126_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3004 _16210_/Q vssd1 vssd1 vccd1 vccd1 hold3004/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold979 hold979/A vssd1 vssd1 vccd1 vccd1 hold979/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3015 _14197_/X vssd1 vssd1 vccd1 vccd1 _17901_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3026 _13955_/X vssd1 vssd1 vccd1 vccd1 _17784_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08943_ hold71/X hold754/X _08991_/S vssd1 vssd1 vccd1 vccd1 _08944_/B sky130_fd_sc_hd__mux2_1
Xhold3037 _16188_/Q vssd1 vssd1 vccd1 vccd1 hold3037/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2303 _14717_/X vssd1 vssd1 vccd1 vccd1 _18150_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3048 _08083_/X vssd1 vssd1 vccd1 vccd1 _15681_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3059 _17789_/Q vssd1 vssd1 vccd1 vccd1 hold3059/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2314 _18065_/Q vssd1 vssd1 vccd1 vccd1 hold2314/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2325 _14041_/X vssd1 vssd1 vccd1 vccd1 _17826_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2336 _08514_/X vssd1 vssd1 vccd1 vccd1 _15884_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08874_ hold131/X hold187/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold188/A sky130_fd_sc_hd__mux2_1
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2347 _17935_/Q vssd1 vssd1 vccd1 vccd1 hold2347/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1602 _15608_/Q vssd1 vssd1 vccd1 vccd1 hold1602/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2358 _08322_/X vssd1 vssd1 vccd1 vccd1 _15794_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1613 _17779_/Q vssd1 vssd1 vccd1 vccd1 hold1613/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1624 _18342_/Q vssd1 vssd1 vccd1 vccd1 hold1624/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2369 _18248_/Q vssd1 vssd1 vccd1 vccd1 hold2369/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1635 _17513_/Q vssd1 vssd1 vccd1 vccd1 hold1635/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07825_ _07809_/X _07810_/Y hold2254/X _09362_/A vssd1 vssd1 vccd1 vccd1 _07825_/X
+ sky130_fd_sc_hd__a2bb2o_1
Xhold1646 _09073_/X vssd1 vssd1 vccd1 vccd1 _16151_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1657 _13959_/X vssd1 vssd1 vccd1 vccd1 _17786_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1668 _16243_/Q vssd1 vssd1 vccd1 vccd1 hold1668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1679 _07917_/X vssd1 vssd1 vccd1 vccd1 _15602_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09426_ hold704/X _16299_/Q vssd1 vssd1 vccd1 vccd1 _09426_/X sky130_fd_sc_hd__or2_1
XFILLER_0_17_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09357_ _09357_/A _09392_/A vssd1 vssd1 vccd1 vccd1 _09386_/B sky130_fd_sc_hd__or2_1
XFILLER_0_19_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08308_ hold1203/X _08323_/B _08307_/X _13795_/C1 vssd1 vssd1 vccd1 vccd1 _08308_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09288_ hold1706/X _09325_/B _09287_/X _12948_/A vssd1 vssd1 vccd1 vccd1 _09288_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08239_ hold2400/X _08262_/B _08238_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _08239_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11250_ _11637_/A _11250_/B vssd1 vssd1 vccd1 vccd1 _11250_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10201_ hold3995/X _10619_/B _10200_/X _14853_/C1 vssd1 vssd1 vccd1 vccd1 _10201_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11181_ hold4350/X _11091_/A _11180_/X vssd1 vssd1 vccd1 vccd1 _11181_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4250 _12334_/Y vssd1 vssd1 vccd1 vccd1 _17268_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10132_ hold4436/X _10628_/B _10131_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10132_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4261 _11155_/Y vssd1 vssd1 vccd1 vccd1 _16875_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4272 _13813_/Y vssd1 vssd1 vccd1 vccd1 _17724_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4283 _11161_/Y vssd1 vssd1 vccd1 vccd1 _16877_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4294 _13864_/Y vssd1 vssd1 vccd1 vccd1 _17741_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3560 _16371_/Q vssd1 vssd1 vccd1 vccd1 hold3560/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10063_ _10603_/A _10063_/B vssd1 vssd1 vccd1 vccd1 _16511_/D sky130_fd_sc_hd__nor2_1
XTAP_6478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14940_ _15209_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14940_/X sky130_fd_sc_hd__or2_1
Xhold3571 _12770_/X vssd1 vssd1 vccd1 vccd1 _12771_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3582 _16475_/Q vssd1 vssd1 vccd1 vccd1 hold3582/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3593 _16649_/Q vssd1 vssd1 vccd1 vccd1 hold3593/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_238_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2870 _14891_/X vssd1 vssd1 vccd1 vccd1 _18234_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14871_ hold2153/X hold332/X _14870_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14871_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2881 _18436_/Q vssd1 vssd1 vccd1 vccd1 hold2881/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2892 _14701_/X vssd1 vssd1 vccd1 vccd1 _18142_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16610_ _18220_/CLK _16610_/D vssd1 vssd1 vccd1 vccd1 _16610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13822_ _13864_/A _13822_/B vssd1 vssd1 vccd1 vccd1 _13822_/Y sky130_fd_sc_hd__nor2_1
X_17590_ _17590_/CLK _17590_/D vssd1 vssd1 vccd1 vccd1 _17590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16541_ _18099_/CLK _16541_/D vssd1 vssd1 vccd1 vccd1 _16541_/Q sky130_fd_sc_hd__dfxtp_1
X_13753_ hold5486/X _13847_/B _13752_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13753_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10965_ _11061_/A _10965_/B vssd1 vssd1 vccd1 vccd1 _10965_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12704_ hold3969/X _12703_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12705_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_214_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16472_ _18385_/CLK _16472_/D vssd1 vssd1 vccd1 vccd1 _16472_/Q sky130_fd_sc_hd__dfxtp_1
X_13684_ hold5527/X _13874_/B _13683_/X _13684_/C1 vssd1 vssd1 vccd1 vccd1 _13684_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10896_ _11088_/A _10896_/B vssd1 vssd1 vccd1 vccd1 _10896_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18211_ _18211_/CLK _18211_/D vssd1 vssd1 vccd1 vccd1 _18211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15423_ _15481_/A1 _15415_/X _15422_/X _15481_/B1 hold5952/A vssd1 vssd1 vccd1 vccd1
+ _15423_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_182_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12635_ hold3357/X _12634_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12635_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18142_ _18174_/CLK _18142_/D vssd1 vssd1 vccd1 vccd1 _18142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15354_ _15394_/A _15354_/B vssd1 vssd1 vccd1 vccd1 _18411_/D sky130_fd_sc_hd__and2_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12566_ hold3636/X _12565_/X _12986_/S vssd1 vssd1 vccd1 vccd1 _12566_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_53_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14305_ hold3112/X _14333_/A2 _14304_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _14305_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11517_ _12285_/A _11517_/B vssd1 vssd1 vccd1 vccd1 _11517_/X sky130_fd_sc_hd__or2_1
X_15285_ hold766/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15285_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18073_ _18073_/CLK hold551/X vssd1 vssd1 vccd1 vccd1 _18073_/Q sky130_fd_sc_hd__dfxtp_1
X_12497_ hold41/X _12509_/A2 _12501_/A3 _12496_/X _09003_/A vssd1 vssd1 vccd1 vccd1
+ hold42/A sky130_fd_sc_hd__o311a_1
XFILLER_0_151_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold209 hold22/X vssd1 vssd1 vccd1 vccd1 input6/A sky130_fd_sc_hd__dlygate4sd3_1
X_14236_ _14970_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14236_/X sky130_fd_sc_hd__or2_1
X_17024_ _17904_/CLK _17024_/D vssd1 vssd1 vccd1 vccd1 _17024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11448_ _11649_/A _11448_/B vssd1 vssd1 vccd1 vccd1 _11448_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_238_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14167_ hold1698/X _14198_/B _14166_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _14167_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11379_ _11661_/A _11379_/B vssd1 vssd1 vccd1 vccd1 _11379_/X sky130_fd_sc_hd__or2_1
XFILLER_0_221_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _13118_/A _13294_/B vssd1 vssd1 vccd1 vccd1 _13118_/X sky130_fd_sc_hd__or2_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ hold992/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14098_/X sky130_fd_sc_hd__or2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ hold5938/X hold907/X _13055_/C vssd1 vssd1 vccd1 vccd1 _13049_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_186_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17926_ _17967_/CLK _17926_/D vssd1 vssd1 vccd1 vccd1 _17926_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17857_ _17890_/CLK _17857_/D vssd1 vssd1 vccd1 vccd1 _17857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16808_ _18043_/CLK _16808_/D vssd1 vssd1 vccd1 vccd1 _16808_/Q sky130_fd_sc_hd__dfxtp_1
X_08590_ hold495/X hold599/X _08592_/S vssd1 vssd1 vccd1 vccd1 hold600/A sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_263_wb_clk_i clkbuf_6_56_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17997_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17788_ _17820_/CLK _17788_/D vssd1 vssd1 vccd1 vccd1 _17788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16739_ _18036_/CLK _16739_/D vssd1 vssd1 vccd1 vccd1 _16739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09211_ hold1823/X _09214_/B _09210_/X _12822_/A vssd1 vssd1 vccd1 vccd1 _09211_/X
+ sky130_fd_sc_hd__o211a_1
X_18409_ _18409_/CLK _18409_/D vssd1 vssd1 vccd1 vccd1 _18409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09142_ _15525_/A _09156_/B vssd1 vssd1 vccd1 vccd1 _09142_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09073_ hold1645/X _09106_/B _09072_/X _12987_/A vssd1 vssd1 vccd1 vccd1 _09073_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08024_ hold1546/X _08029_/B _08023_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _08024_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold710 hold710/A vssd1 vssd1 vccd1 vccd1 hold710/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_241_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold721 hold721/A vssd1 vssd1 vccd1 vccd1 hold721/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold732 hold732/A vssd1 vssd1 vccd1 vccd1 hold732/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold743 hold743/A vssd1 vssd1 vccd1 vccd1 hold743/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 hold754/A vssd1 vssd1 vccd1 vccd1 hold754/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold765 hold765/A vssd1 vssd1 vccd1 vccd1 hold765/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold776 hold776/A vssd1 vssd1 vccd1 vccd1 hold776/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold787 hold787/A vssd1 vssd1 vccd1 vccd1 hold787/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold798 hold798/A vssd1 vssd1 vccd1 vccd1 hold798/X sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ _10986_/A _09975_/B vssd1 vssd1 vccd1 vccd1 _09975_/X sky130_fd_sc_hd__or2_1
Xhold2100 _18174_/Q vssd1 vssd1 vccd1 vccd1 hold2100/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2111 _18172_/Q vssd1 vssd1 vccd1 vccd1 hold2111/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08926_ hold87/X hold516/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold517/A sky130_fd_sc_hd__mux2_1
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2122 _14031_/X vssd1 vssd1 vccd1 vccd1 _17821_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2133 _18048_/Q vssd1 vssd1 vccd1 vccd1 hold2133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2144 _14945_/X vssd1 vssd1 vccd1 vccd1 _18259_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1410 _14043_/X vssd1 vssd1 vccd1 vccd1 _17827_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2155 _18446_/Q vssd1 vssd1 vccd1 vccd1 hold2155/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2166 _14235_/X vssd1 vssd1 vccd1 vccd1 _17918_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1421 _14283_/X vssd1 vssd1 vccd1 vccd1 _17942_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1432 _18288_/Q vssd1 vssd1 vccd1 vccd1 hold1432/X sky130_fd_sc_hd__dlygate4sd3_1
X_08857_ _15473_/A _08857_/B vssd1 vssd1 vccd1 vccd1 _16047_/D sky130_fd_sc_hd__and2_1
XFILLER_0_207_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2177 _18237_/Q vssd1 vssd1 vccd1 vccd1 hold2177/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2188 _14995_/X vssd1 vssd1 vccd1 vccd1 _18283_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1443 _08493_/X vssd1 vssd1 vccd1 vccd1 _15875_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2199 _17919_/Q vssd1 vssd1 vccd1 vccd1 hold2199/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1454 _15532_/X vssd1 vssd1 vccd1 vccd1 _18444_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1465 hold1465/A vssd1 vssd1 vccd1 vccd1 _15195_/A sky130_fd_sc_hd__buf_12
X_07808_ _15314_/A _13048_/A _07803_/Y hold2275/X vssd1 vssd1 vccd1 vccd1 _07808_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1476 _15180_/X vssd1 vssd1 vccd1 vccd1 _18373_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08788_ _15482_/A hold464/X vssd1 vssd1 vccd1 vccd1 _16014_/D sky130_fd_sc_hd__and2_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1487 _18032_/Q vssd1 vssd1 vccd1 vccd1 hold1487/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1498 _08497_/X vssd1 vssd1 vccd1 vccd1 _15877_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ hold4085/X _11071_/A2 _10749_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _10750_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09409_ _07804_/A _09447_/B _09440_/B _09408_/X vssd1 vssd1 vccd1 vccd1 _09409_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10681_ hold4668/X _11162_/B _10680_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _10681_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12420_ _12420_/A _12420_/B vssd1 vssd1 vccd1 vccd1 _17303_/D sky130_fd_sc_hd__and2_1
XFILLER_0_164_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12351_ hold5714/X _12255_/A _12350_/X vssd1 vssd1 vccd1 vccd1 _12351_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_wb_clk_i clkbuf_6_19_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17291_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11302_ hold4109/X _12323_/B _11301_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11302_/X
+ sky130_fd_sc_hd__o211a_1
X_15070_ _15070_/A hold290/X vssd1 vssd1 vccd1 vccd1 hold291/A sky130_fd_sc_hd__and2_1
XFILLER_0_205_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12282_ _13407_/A _12282_/B vssd1 vssd1 vccd1 vccd1 _12282_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_1365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14021_ hold1859/X _14038_/B _14020_/X _12588_/A vssd1 vssd1 vccd1 vccd1 _14021_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11233_ hold4091/X _11717_/B _11232_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11233_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11164_ _11203_/A _11164_/B vssd1 vssd1 vccd1 vccd1 _11164_/Y sky130_fd_sc_hd__nor2_1
XTAP_6231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4080 _11140_/X vssd1 vssd1 vccd1 vccd1 _16870_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10115_ hold3033/X hold3499/X _10595_/C vssd1 vssd1 vccd1 vccd1 _10116_/B sky130_fd_sc_hd__mux2_1
Xhold4091 _16933_/Q vssd1 vssd1 vccd1 vccd1 hold4091/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15972_ _18462_/CLK _15972_/D vssd1 vssd1 vccd1 vccd1 hold846/A sky130_fd_sc_hd__dfxtp_1
X_11095_ hold5152/X _11225_/B _11094_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _11095_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17711_ _17744_/CLK _17711_/D vssd1 vssd1 vccd1 vccd1 _17711_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3390 _17453_/Q vssd1 vssd1 vccd1 vccd1 hold3390/X sky130_fd_sc_hd__dlygate4sd3_1
X_14923_ hold2369/X _14946_/B _14922_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _14923_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10046_ _16506_/Q _10046_/B _10067_/C vssd1 vssd1 vccd1 vccd1 _10046_/X sky130_fd_sc_hd__and3_1
XFILLER_0_234_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__buf_1
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_153_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17642_ _17738_/CLK _17642_/D vssd1 vssd1 vccd1 vccd1 _17642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14854_ _15085_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14854_/X sky130_fd_sc_hd__or2_1
XFILLER_0_203_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13805_ _17722_/Q _13808_/B _13814_/C vssd1 vssd1 vccd1 vccd1 _13805_/X sky130_fd_sc_hd__and3_1
XFILLER_0_188_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17573_ _17739_/CLK _17573_/D vssd1 vssd1 vccd1 vccd1 _17573_/Q sky130_fd_sc_hd__dfxtp_1
X_14785_ hold1598/X _14772_/B _14784_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14785_/X
+ sky130_fd_sc_hd__o211a_1
X_11997_ _12093_/A _11997_/B vssd1 vssd1 vccd1 vccd1 _11997_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16524_ _18146_/CLK _16524_/D vssd1 vssd1 vccd1 vccd1 _16524_/Q sky130_fd_sc_hd__dfxtp_1
X_10948_ hold5241/X _11732_/B _10947_/X _13895_/A vssd1 vssd1 vccd1 vccd1 _10948_/X
+ sky130_fd_sc_hd__o211a_1
X_13736_ hold2322/X hold4764/X _13862_/C vssd1 vssd1 vccd1 vccd1 _13737_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_58_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16455_ _18368_/CLK _16455_/D vssd1 vssd1 vccd1 vccd1 _16455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13667_ hold1115/X _17676_/Q _13883_/C vssd1 vssd1 vccd1 vccd1 _13668_/B sky130_fd_sc_hd__mux2_1
X_10879_ hold5066/X _11165_/B _10878_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _10879_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15406_ _17344_/Q _15486_/B1 _15485_/B1 hold280/X vssd1 vssd1 vccd1 vccd1 _15406_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12618_ _12864_/A _12618_/B vssd1 vssd1 vccd1 vccd1 _17382_/D sky130_fd_sc_hd__and2_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16386_ _18363_/CLK _16386_/D vssd1 vssd1 vccd1 vccd1 _16386_/Q sky130_fd_sc_hd__dfxtp_1
X_13598_ hold1566/X _17653_/Q _13877_/C vssd1 vssd1 vccd1 vccd1 _13599_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_170_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18125_ _18125_/CLK _18125_/D vssd1 vssd1 vccd1 vccd1 _18125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15337_ hold575/X _09357_/A _09386_/D hold741/X _15336_/X vssd1 vssd1 vccd1 vccd1
+ _15342_/B sky130_fd_sc_hd__a221o_1
X_12549_ _12924_/A _12549_/B vssd1 vssd1 vccd1 vccd1 _17359_/D sky130_fd_sc_hd__and2_1
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5709 _12360_/Y vssd1 vssd1 vccd1 vccd1 _12361_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_1 _13052_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_26_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_26_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_18056_ _18056_/CLK _18056_/D vssd1 vssd1 vccd1 vccd1 _18056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15268_ hold539/X _09386_/A _09392_/D hold847/X vssd1 vssd1 vccd1 vccd1 _15268_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17007_ _17887_/CLK _17007_/D vssd1 vssd1 vccd1 vccd1 _17007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14219_ hold2119/X _14216_/Y _14218_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _14219_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15199_ _15199_/A _15227_/B vssd1 vssd1 vccd1 vccd1 _15199_/X sky130_fd_sc_hd__or2_1
XFILLER_0_238_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout508 _10538_/S vssd1 vssd1 vccd1 vccd1 _10604_/C sky130_fd_sc_hd__buf_4
Xfanout519 _10619_/C vssd1 vssd1 vccd1 vccd1 _10595_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09760_ hold3614/X _10046_/B _09759_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09760_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_225_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_444_wb_clk_i clkbuf_6_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _15886_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08711_ hold92/X hold533/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold534/A sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17909_ _18428_/CLK _17909_/D vssd1 vssd1 vccd1 vccd1 _17909_/Q sky130_fd_sc_hd__dfxtp_1
X_09691_ hold3584/X _10601_/B _09690_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09691_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08642_ _15324_/A _08642_/B vssd1 vssd1 vccd1 vccd1 _15943_/D sky130_fd_sc_hd__and2_1
XFILLER_0_221_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08573_ _09047_/A _08573_/B vssd1 vssd1 vccd1 vccd1 _15910_/D sky130_fd_sc_hd__and2_1
XFILLER_0_156_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_234_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09125_ _15128_/A hold363/X vssd1 vssd1 vccd1 vccd1 _09156_/B sky130_fd_sc_hd__or2_2
XFILLER_0_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09056_ hold87/X hold124/X _09056_/S vssd1 vssd1 vccd1 vccd1 hold125/A sky130_fd_sc_hd__mux2_1
XFILLER_0_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08007_ _15521_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08007_/X sky130_fd_sc_hd__or2_1
Xhold540 hold540/A vssd1 vssd1 vccd1 vccd1 hold540/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_241_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold551 hold551/A vssd1 vssd1 vccd1 vccd1 hold551/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 hold562/A vssd1 vssd1 vccd1 vccd1 hold562/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold573 hold573/A vssd1 vssd1 vccd1 vccd1 hold573/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold584 hold584/A vssd1 vssd1 vccd1 vccd1 hold584/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold595 hold595/A vssd1 vssd1 vccd1 vccd1 input45/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_229_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_217_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09958_ hold3554/X _10052_/B _09957_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _09958_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_217_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_185_wb_clk_i clkbuf_6_54_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18361_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08909_ _12420_/A _08909_/B vssd1 vssd1 vccd1 vccd1 _16072_/D sky130_fd_sc_hd__and2_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_114_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17335_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09889_ hold4528/X _10025_/B _09888_/X _08954_/A vssd1 vssd1 vccd1 vccd1 _09889_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1240 _13971_/X vssd1 vssd1 vccd1 vccd1 _17792_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1251 hold640/X vssd1 vssd1 vccd1 vccd1 input43/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1262 _18309_/Q vssd1 vssd1 vccd1 vccd1 hold1262/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ hold4787/X _12293_/B _11919_/X _12103_/C1 vssd1 vssd1 vccd1 vccd1 _11920_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1273 _17895_/Q vssd1 vssd1 vccd1 vccd1 hold1273/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1284 _14895_/X vssd1 vssd1 vccd1 vccd1 _18236_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1295 _18055_/Q vssd1 vssd1 vccd1 vccd1 hold1295/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ hold5699/X _12329_/B _11850_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _11851_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ hold2408/X hold4909/X _11186_/C vssd1 vssd1 vccd1 vccd1 _10803_/B sky130_fd_sc_hd__mux2_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _15492_/A _14573_/B hold2238/X vssd1 vssd1 vccd1 vccd1 _14570_/X sky130_fd_sc_hd__a21o_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11782_ _13864_/A _11782_/B vssd1 vssd1 vccd1 vccd1 _11782_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_32_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10733_ hold1915/X hold4347/X _11213_/C vssd1 vssd1 vccd1 vccd1 _10734_/B sky130_fd_sc_hd__mux2_1
X_13521_ _13722_/A _13521_/B vssd1 vssd1 vccd1 vccd1 _13521_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13452_ _13773_/A _13452_/B vssd1 vssd1 vccd1 vccd1 _13452_/X sky130_fd_sc_hd__or2_1
X_16240_ _17661_/CLK _16240_/D vssd1 vssd1 vccd1 vccd1 _16240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10664_ hold1117/X hold3508/X _11144_/C vssd1 vssd1 vccd1 vccd1 _10665_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12403_ hold163/X hold749/X _12441_/S vssd1 vssd1 vccd1 vccd1 hold750/A sky130_fd_sc_hd__mux2_1
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16171_ _17492_/CLK _16171_/D vssd1 vssd1 vccd1 vccd1 _16171_/Q sky130_fd_sc_hd__dfxtp_1
X_13383_ _13737_/A _13383_/B vssd1 vssd1 vccd1 vccd1 _13383_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10595_ _16689_/Q _10619_/B _10595_/C vssd1 vssd1 vccd1 vccd1 _10595_/X sky130_fd_sc_hd__and3_1
XFILLER_0_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15122_ hold2950/X hold340/X _15121_/X _15176_/C1 vssd1 vssd1 vccd1 vccd1 _15122_/X
+ sky130_fd_sc_hd__o211a_1
X_12334_ _13873_/A _12334_/B vssd1 vssd1 vccd1 vccd1 _12334_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_105_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15053_ hold384/X hold833/X _15071_/S vssd1 vssd1 vccd1 vccd1 hold834/A sky130_fd_sc_hd__mux2_1
XFILLER_0_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12265_ hold5737/X _12362_/B _12264_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _12265_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14004_ hold915/X _14042_/B vssd1 vssd1 vccd1 vccd1 _14004_/X sky130_fd_sc_hd__or2_1
XFILLER_0_142_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11216_ _16896_/Q _11225_/B _11216_/C vssd1 vssd1 vccd1 vccd1 _11216_/X sky130_fd_sc_hd__and3_1
XFILLER_0_103_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12196_ hold4795/X _12308_/B _12195_/X _08167_/A vssd1 vssd1 vccd1 vccd1 _12196_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput82 _13209_/A vssd1 vssd1 vccd1 vccd1 output82/X sky130_fd_sc_hd__buf_6
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput93 _13289_/A vssd1 vssd1 vccd1 vccd1 output93/X sky130_fd_sc_hd__buf_6
XTAP_6050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11147_ _16873_/Q _11153_/B _11153_/C vssd1 vssd1 vccd1 vccd1 _11147_/X sky130_fd_sc_hd__and3_1
XTAP_6061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15955_ _16098_/CLK _15955_/D vssd1 vssd1 vccd1 vccd1 hold791/A sky130_fd_sc_hd__dfxtp_1
XTAP_5360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11078_ hold2800/X _16850_/Q _11753_/C vssd1 vssd1 vccd1 vccd1 _11079_/B sky130_fd_sc_hd__mux2_1
XTAP_5371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10029_ _13190_/A _09933_/A _10028_/X vssd1 vssd1 vccd1 vccd1 _10029_/Y sky130_fd_sc_hd__a21oi_1
X_14906_ hold945/X _14910_/B vssd1 vssd1 vccd1 vccd1 _14906_/X sky130_fd_sc_hd__or2_1
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15886_ _15886_/CLK _15886_/D vssd1 vssd1 vccd1 vccd1 _15886_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17625_ _17722_/CLK _17625_/D vssd1 vssd1 vccd1 vccd1 _17625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14837_ hold2936/X _14828_/B _14836_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _14837_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17556_ _18191_/CLK _17556_/D vssd1 vssd1 vccd1 vccd1 _17556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14768_ _15161_/A _14772_/B vssd1 vssd1 vccd1 vccd1 _14768_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16507_ _18396_/CLK _16507_/D vssd1 vssd1 vccd1 vccd1 _16507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13719_ _13719_/A _13719_/B vssd1 vssd1 vccd1 vccd1 _13719_/X sky130_fd_sc_hd__or2_1
XFILLER_0_89_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17487_ _17491_/CLK _17487_/D vssd1 vssd1 vccd1 vccd1 _17487_/Q sky130_fd_sc_hd__dfxtp_1
X_14699_ hold3082/X _14718_/B _14698_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _14699_/X
+ sky130_fd_sc_hd__o211a_1
X_16438_ _18383_/CLK _16438_/D vssd1 vssd1 vccd1 vccd1 _16438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16369_ _18323_/CLK _16369_/D vssd1 vssd1 vccd1 vccd1 _16369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18108_ _18214_/CLK _18108_/D vssd1 vssd1 vccd1 vccd1 _18108_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5506 _11350_/X vssd1 vssd1 vccd1 vccd1 _16940_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5517 _16970_/Q vssd1 vssd1 vccd1 vccd1 hold5517/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5528 _13684_/X vssd1 vssd1 vccd1 vccd1 _17681_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5539 _16974_/Q vssd1 vssd1 vccd1 vccd1 hold5539/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4805 _17128_/Q vssd1 vssd1 vccd1 vccd1 hold4805/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18039_ _18039_/CLK _18039_/D vssd1 vssd1 vccd1 vccd1 _18039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4816 _12067_/X vssd1 vssd1 vccd1 vccd1 _17179_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4827 _17194_/Q vssd1 vssd1 vccd1 vccd1 hold4827/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4838 _10777_/X vssd1 vssd1 vccd1 vccd1 _16749_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4849 _16466_/Q vssd1 vssd1 vccd1 vccd1 hold4849/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout305 _11106_/A vssd1 vssd1 vccd1 vccd1 _09987_/A sky130_fd_sc_hd__buf_4
Xfanout316 _10539_/A vssd1 vssd1 vccd1 vccd1 _10563_/A sky130_fd_sc_hd__buf_4
Xfanout327 _10386_/A vssd1 vssd1 vccd1 vccd1 _09954_/A sky130_fd_sc_hd__buf_4
X_09812_ hold2605/X hold4509/X _10028_/C vssd1 vssd1 vccd1 vccd1 _09813_/B sky130_fd_sc_hd__mux2_1
Xfanout338 _12506_/B vssd1 vssd1 vccd1 vccd1 _12498_/B sky130_fd_sc_hd__clkbuf_8
Xfanout349 _08934_/X vssd1 vssd1 vccd1 vccd1 _08997_/S sky130_fd_sc_hd__buf_8
XFILLER_0_201_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09743_ hold2536/X hold4034/X _10031_/C vssd1 vssd1 vccd1 vccd1 _09744_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_236_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09674_ hold1235/X _16382_/Q _10538_/S vssd1 vssd1 vccd1 vccd1 _09675_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08625_ hold169/X hold585/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold586/A sky130_fd_sc_hd__mux2_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08556_ hold77/X hold587/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08557_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08487_ hold2386/X _08486_/B _08486_/Y _08133_/A vssd1 vssd1 vccd1 vccd1 _08487_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09108_ _15169_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09108_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10380_ _10476_/A _10380_/B vssd1 vssd1 vccd1 vccd1 _10380_/X sky130_fd_sc_hd__or2_1
XFILLER_0_143_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09039_ _15374_/A _09039_/B vssd1 vssd1 vccd1 vccd1 _16136_/D sky130_fd_sc_hd__and2_1
XFILLER_0_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_366_wb_clk_i clkbuf_6_34_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17606_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12050_ hold1352/X hold4863/X _12242_/S vssd1 vssd1 vccd1 vccd1 _12051_/B sky130_fd_sc_hd__mux2_1
Xhold370 hold370/A vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 la_data_in[16] vssd1 vssd1 vccd1 vccd1 hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 hold392/A vssd1 vssd1 vccd1 vccd1 hold392/X sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ _11661_/A _11001_/B vssd1 vssd1 vccd1 vccd1 _11001_/X sky130_fd_sc_hd__or2_1
Xfanout850 _17754_/Q vssd1 vssd1 vccd1 vccd1 _12337_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_232_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout872 _14952_/A vssd1 vssd1 vccd1 vccd1 _15547_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_102_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout883 hold932/X vssd1 vssd1 vccd1 vccd1 _14517_/A sky130_fd_sc_hd__buf_12
Xfanout894 hold945/X vssd1 vssd1 vccd1 vccd1 _15191_/A sky130_fd_sc_hd__buf_8
X_15740_ _17744_/CLK _15740_/D vssd1 vssd1 vccd1 vccd1 _15740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12952_ hold1386/X _17495_/Q _12985_/S vssd1 vssd1 vccd1 vccd1 _12952_/X sky130_fd_sc_hd__mux2_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1070 _17866_/Q vssd1 vssd1 vccd1 vccd1 hold1070/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1081 _15816_/Q vssd1 vssd1 vccd1 vccd1 hold1081/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ hold2077/X hold4670/X _13796_/S vssd1 vssd1 vccd1 vccd1 _11904_/B sky130_fd_sc_hd__mux2_1
Xhold1092 _07951_/X vssd1 vssd1 vccd1 vccd1 _15618_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _17878_/CLK _15671_/D vssd1 vssd1 vccd1 vccd1 _15671_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ hold3037/X _17472_/Q _12916_/S vssd1 vssd1 vccd1 vccd1 _12883_/X sky130_fd_sc_hd__mux2_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _17434_/CLK _17410_/D vssd1 vssd1 vccd1 vccd1 _17410_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14622_ _15231_/A _14622_/B vssd1 vssd1 vccd1 vccd1 _14622_/X sky130_fd_sc_hd__or2_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _18390_/CLK _18390_/D vssd1 vssd1 vccd1 vccd1 _18390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11834_ hold2525/X hold4267/X _13481_/S vssd1 vssd1 vccd1 vccd1 _11835_/B sky130_fd_sc_hd__mux2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _17341_/CLK hold42/X vssd1 vssd1 vccd1 vccd1 _17341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _17079_/Q _11765_/B _11765_/C vssd1 vssd1 vccd1 vccd1 _11765_/X sky130_fd_sc_hd__and3_1
X_14553_ hold579/A _14553_/B vssd1 vssd1 vccd1 vccd1 hold550/A sky130_fd_sc_hd__or2_1
XFILLER_0_166_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_82_wb_clk_i clkbuf_6_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17491_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13504_ hold4154/X _13880_/B _13503_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13504_/X
+ sky130_fd_sc_hd__o211a_1
X_10716_ _11100_/A _10716_/B vssd1 vssd1 vccd1 vccd1 _10716_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17272_ _17272_/CLK _17272_/D vssd1 vssd1 vccd1 vccd1 _17272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_1300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_wb_clk_i clkbuf_6_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18447_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11696_ hold2603/X hold5400/X _12335_/C vssd1 vssd1 vccd1 vccd1 _11697_/B sky130_fd_sc_hd__mux2_1
X_14484_ hold1348/X _14487_/B _14483_/Y _14376_/A vssd1 vssd1 vccd1 vccd1 _14484_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16223_ _17452_/CLK _16223_/D vssd1 vssd1 vccd1 vccd1 _16223_/Q sky130_fd_sc_hd__dfxtp_1
X_10647_ hold4245/X _10551_/A _10646_/X vssd1 vssd1 vccd1 vccd1 _10647_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13435_ hold3646/X _13829_/B _13434_/X _13795_/C1 vssd1 vssd1 vccd1 vccd1 _13435_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16154_ _17491_/CLK _16154_/D vssd1 vssd1 vccd1 vccd1 _16154_/Q sky130_fd_sc_hd__dfxtp_1
X_13366_ hold4985/X _13886_/B _13365_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _13366_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10578_ hold3423/X _10386_/A _10577_/X vssd1 vssd1 vccd1 vccd1 _10578_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_183_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15105_ hold641/X _15125_/B vssd1 vssd1 vccd1 vccd1 hold642/A sky130_fd_sc_hd__or2_1
XFILLER_0_121_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12317_ _17263_/Q _12317_/B _12317_/C vssd1 vssd1 vccd1 vccd1 _12317_/X sky130_fd_sc_hd__and3_1
X_13297_ _13297_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13297_/X sky130_fd_sc_hd__and2_1
X_16085_ _17293_/CLK _16085_/D vssd1 vssd1 vccd1 vccd1 hold720/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15036_ _15394_/A hold368/X vssd1 vssd1 vccd1 vccd1 hold369/A sky130_fd_sc_hd__and2_1
XFILLER_0_20_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12248_ hold1205/X hold4913/X _13748_/S vssd1 vssd1 vccd1 vccd1 _12249_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_208_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12179_ hold1556/X hold5078/X _13748_/S vssd1 vssd1 vccd1 vccd1 _12180_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_208_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16987_ _17823_/CLK _16987_/D vssd1 vssd1 vccd1 vccd1 _16987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15938_ _17297_/CLK _15938_/D vssd1 vssd1 vccd1 vccd1 _15938_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15869_ _17740_/CLK _15869_/D vssd1 vssd1 vccd1 vccd1 _15869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08410_ hold1052/X _08442_/A2 _08409_/X _13795_/C1 vssd1 vssd1 vccd1 vccd1 _08410_/X
+ sky130_fd_sc_hd__o211a_1
X_17608_ _17608_/CLK _17608_/D vssd1 vssd1 vccd1 vccd1 _17608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09390_ _09369_/C _09389_/X _07809_/B vssd1 vssd1 vccd1 vccd1 _09390_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08341_ _08347_/A _08341_/B vssd1 vssd1 vccd1 vccd1 _15802_/D sky130_fd_sc_hd__and2_1
XFILLER_0_59_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17539_ _18380_/CLK _17539_/D vssd1 vssd1 vccd1 vccd1 _17539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08272_ hold992/X _08280_/B vssd1 vssd1 vccd1 vccd1 _08272_/X sky130_fd_sc_hd__or2_1
XFILLER_0_6_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_229_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6004 _17552_/Q vssd1 vssd1 vccd1 vccd1 hold6004/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6015 _17535_/Q vssd1 vssd1 vccd1 vccd1 hold6015/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6026 _17545_/Q vssd1 vssd1 vccd1 vccd1 hold6026/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6037 data_in[15] vssd1 vssd1 vccd1 vccd1 hold177/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5303 _16791_/Q vssd1 vssd1 vccd1 vccd1 hold5303/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6048 data_in[30] vssd1 vssd1 vccd1 vccd1 hold317/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold6059 _18290_/Q vssd1 vssd1 vccd1 vccd1 hold6059/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5314 _11407_/X vssd1 vssd1 vccd1 vccd1 _16959_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5325 _17617_/Q vssd1 vssd1 vccd1 vccd1 hold5325/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5336 _10813_/X vssd1 vssd1 vccd1 vccd1 _16761_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4602 _16674_/Q vssd1 vssd1 vccd1 vccd1 hold4602/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5347 _16990_/Q vssd1 vssd1 vccd1 vccd1 hold5347/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5358 _13360_/X vssd1 vssd1 vccd1 vccd1 _17573_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4613 _13726_/X vssd1 vssd1 vccd1 vccd1 _17695_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4624 _17730_/Q vssd1 vssd1 vccd1 vccd1 hold4624/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5369 _11437_/X vssd1 vssd1 vccd1 vccd1 _16969_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4635 _11137_/X vssd1 vssd1 vccd1 vccd1 _16869_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3901 _16562_/Q vssd1 vssd1 vccd1 vccd1 hold3901/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4646 _17134_/Q vssd1 vssd1 vccd1 vccd1 hold4646/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3912 _09607_/X vssd1 vssd1 vccd1 vccd1 _16359_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4657 _09637_/X vssd1 vssd1 vccd1 vccd1 _16369_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4668 _16749_/Q vssd1 vssd1 vccd1 vccd1 hold4668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3923 _17728_/Q vssd1 vssd1 vccd1 vccd1 _13823_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3934 _10897_/X vssd1 vssd1 vccd1 vccd1 _16789_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4679 _16392_/Q vssd1 vssd1 vccd1 vccd1 hold4679/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3945 _09964_/X vssd1 vssd1 vccd1 vccd1 _16478_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3956 _16863_/Q vssd1 vssd1 vccd1 vccd1 hold3956/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3967 _17658_/Q vssd1 vssd1 vccd1 vccd1 hold3967/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3978 _16740_/Q vssd1 vssd1 vccd1 vccd1 hold3978/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout157 _12971_/S vssd1 vssd1 vccd1 vccd1 _12986_/S sky130_fd_sc_hd__buf_4
Xhold3989 _17679_/Q vssd1 vssd1 vccd1 vccd1 hold3989/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout168 _12217_/A2 vssd1 vssd1 vccd1 vccd1 _13795_/A2 sky130_fd_sc_hd__clkbuf_8
X_07987_ hold1604/X _07978_/B _07986_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _07987_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout179 _11741_/B vssd1 vssd1 vccd1 vccd1 _12323_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_226_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09726_ _09984_/A _09726_/B vssd1 vssd1 vccd1 vccd1 _09726_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_215_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09657_ _11109_/A _09657_/B vssd1 vssd1 vccd1 vccd1 _09657_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08608_ _15244_/A _08608_/B vssd1 vssd1 vccd1 vccd1 _15926_/D sky130_fd_sc_hd__and2_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09588_ _10476_/A _09588_/B vssd1 vssd1 vccd1 vccd1 _09588_/X sky130_fd_sc_hd__or2_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08539_ _12440_/A hold816/X vssd1 vssd1 vccd1 vccd1 _15893_/D sky130_fd_sc_hd__and2_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11550_ _11553_/A _11550_/B vssd1 vssd1 vccd1 vccd1 _11550_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10501_ hold3832/X _10619_/B _10500_/X _14853_/C1 vssd1 vssd1 vccd1 vccd1 _10501_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11481_ _12174_/A _11481_/B vssd1 vssd1 vccd1 vccd1 _11481_/X sky130_fd_sc_hd__or2_1
XFILLER_0_208_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13220_ hold4531/X _13219_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13220_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10432_ hold3761/X _10649_/B _10431_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10432_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13151_ _13311_/A1 hold5997/X _13150_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13151_/X
+ sky130_fd_sc_hd__o211a_1
X_10363_ hold3795/X _10649_/B _10362_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10363_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12102_ _12198_/A _12102_/B vssd1 vssd1 vccd1 vccd1 _12102_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5870 output74/X vssd1 vssd1 vccd1 vccd1 data_out[11] sky130_fd_sc_hd__buf_12
X_13082_ _17561_/Q _17095_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13082_/X sky130_fd_sc_hd__mux2_1
Xhold5881 hold6025/X vssd1 vssd1 vccd1 vccd1 _13201_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10294_ hold3668/X _10625_/B _10293_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _10294_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5892 output95/X vssd1 vssd1 vccd1 vccd1 data_out[30] sky130_fd_sc_hd__buf_12
XFILLER_0_40_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12033_ _13314_/A _12033_/B vssd1 vssd1 vccd1 vccd1 _12033_/X sky130_fd_sc_hd__or2_1
X_16910_ _17886_/CLK _16910_/D vssd1 vssd1 vccd1 vccd1 _16910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17890_ _17890_/CLK _17890_/D vssd1 vssd1 vccd1 vccd1 _17890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16841_ _18461_/CLK _16841_/D vssd1 vssd1 vccd1 vccd1 _16841_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout680 _14356_/A vssd1 vssd1 vccd1 vccd1 _13895_/A sky130_fd_sc_hd__buf_4
XFILLER_0_137_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout691 _12987_/A vssd1 vssd1 vccd1 vccd1 _12984_/A sky130_fd_sc_hd__buf_4
X_16772_ _18039_/CLK _16772_/D vssd1 vssd1 vccd1 vccd1 _16772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13984_ _15545_/A _13986_/B vssd1 vssd1 vccd1 vccd1 _13984_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_189_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15723_ _17259_/CLK _15723_/D vssd1 vssd1 vccd1 vccd1 _15723_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ hold4447/X _12934_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12935_/X sky130_fd_sc_hd__mux2_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ _18453_/CLK _18442_/D vssd1 vssd1 vccd1 vccd1 _18442_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15654_ _17167_/CLK _15654_/D vssd1 vssd1 vccd1 vccd1 _15654_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ hold3288/X _12865_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12866_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_185_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ hold1984/X _14612_/B _14604_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14605_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_1331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18373_ _18373_/CLK _18373_/D vssd1 vssd1 vccd1 vccd1 _18373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11817_ _13716_/A _11817_/B vssd1 vssd1 vccd1 vccd1 _11817_/X sky130_fd_sc_hd__or2_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _17264_/CLK _15585_/D vssd1 vssd1 vccd1 vccd1 _15585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12797_ hold3392/X _12796_/X _12812_/S vssd1 vssd1 vccd1 vccd1 _12797_/X sky130_fd_sc_hd__mux2_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17324_ _17324_/CLK hold204/X vssd1 vssd1 vccd1 vccd1 _17324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ hold3017/X _14541_/B _14535_/Y _14348_/A vssd1 vssd1 vccd1 vccd1 _14536_/X
+ sky130_fd_sc_hd__o211a_1
X_11748_ hold4430/X _12219_/A _11747_/X vssd1 vssd1 vccd1 vccd1 _11748_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17255_ _18445_/CLK _17255_/D vssd1 vssd1 vccd1 vccd1 _17255_/Q sky130_fd_sc_hd__dfxtp_1
X_14467_ _15201_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14467_/X sky130_fd_sc_hd__or2_1
X_11679_ _12243_/A _11679_/B vssd1 vssd1 vccd1 vccd1 _11679_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_288_wb_clk_i clkbuf_6_37_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18052_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16206_ _17435_/CLK _16206_/D vssd1 vssd1 vccd1 vccd1 _16206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13418_ hold2987/X _17593_/Q _13817_/C vssd1 vssd1 vccd1 vccd1 _13419_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17186_ _17250_/CLK _17186_/D vssd1 vssd1 vccd1 vccd1 _17186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14398_ hold2083/X _14446_/A2 _14397_/X _14342_/A vssd1 vssd1 vccd1 vccd1 _14398_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_217_wb_clk_i clkbuf_6_61_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18087_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16137_ _17297_/CLK _16137_/D vssd1 vssd1 vccd1 vccd1 hold156/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13349_ hold998/X hold4239/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13350_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_11_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3208 _16547_/Q vssd1 vssd1 vccd1 vccd1 hold3208/X sky130_fd_sc_hd__dlygate4sd3_1
X_16068_ _17300_/CLK _16068_/D vssd1 vssd1 vccd1 vccd1 hold728/A sky130_fd_sc_hd__dfxtp_1
Xhold3219 _09535_/X vssd1 vssd1 vccd1 vccd1 _16335_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15019_ hold1235/X hold447/X _15018_/X _15019_/C1 vssd1 vssd1 vccd1 vccd1 _15019_/X
+ sky130_fd_sc_hd__o211a_1
X_07910_ _15533_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07910_/X sky130_fd_sc_hd__or2_1
X_08890_ hold23/X hold322/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08891_/B sky130_fd_sc_hd__mux2_1
Xhold2507 _17963_/Q vssd1 vssd1 vccd1 vccd1 hold2507/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2518 _18137_/Q vssd1 vssd1 vccd1 vccd1 hold2518/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2529 _14827_/X vssd1 vssd1 vccd1 vccd1 _18203_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07841_ _15085_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07841_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1806 _15226_/X vssd1 vssd1 vccd1 vccd1 _18395_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1817 _15633_/Q vssd1 vssd1 vccd1 vccd1 hold1817/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1828 _14997_/X vssd1 vssd1 vccd1 vccd1 _18284_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1839 _18165_/Q vssd1 vssd1 vccd1 vccd1 hold1839/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09511_ hold3648/X _10004_/B _09510_/X _15482_/A vssd1 vssd1 vccd1 vccd1 _09511_/X
+ sky130_fd_sc_hd__o211a_1
X_09442_ _09447_/C _09447_/D _09478_/B vssd1 vssd1 vccd1 vccd1 _09442_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ _17325_/Q _15487_/A2 _09392_/B _16102_/Q vssd1 vssd1 vccd1 vccd1 _09373_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_231_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08324_ hold2326/X _08323_/B _08323_/Y _13801_/C1 vssd1 vssd1 vccd1 vccd1 _08324_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08255_ hold2861/X _08262_/B _08254_/X _08347_/A vssd1 vssd1 vccd1 vccd1 _08255_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08186_ hold1123/X _08209_/B _08185_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _08186_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5100 _11815_/X vssd1 vssd1 vccd1 vccd1 _17095_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5111 _17010_/Q vssd1 vssd1 vccd1 vccd1 hold5111/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5122 _11887_/X vssd1 vssd1 vccd1 vccd1 _17119_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5133 _17048_/Q vssd1 vssd1 vccd1 vccd1 hold5133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5144 _16682_/Q vssd1 vssd1 vccd1 vccd1 hold5144/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4410 _13858_/Y vssd1 vssd1 vccd1 vccd1 _17739_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5155 _10921_/X vssd1 vssd1 vccd1 vccd1 _16797_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4421 _17578_/Q vssd1 vssd1 vccd1 vccd1 hold4421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5166 _10888_/X vssd1 vssd1 vccd1 vccd1 _16786_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5177 _16454_/Q vssd1 vssd1 vccd1 vccd1 hold5177/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4432 _11749_/Y vssd1 vssd1 vccd1 vccd1 _17073_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4443 _13866_/Y vssd1 vssd1 vccd1 vccd1 _13867_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5188 _10849_/X vssd1 vssd1 vccd1 vccd1 _16773_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5199 _17060_/Q vssd1 vssd1 vccd1 vccd1 hold5199/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4454 _16906_/Q vssd1 vssd1 vccd1 vccd1 hold4454/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3720 _16646_/Q vssd1 vssd1 vccd1 vccd1 hold3720/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4465 _16630_/Q vssd1 vssd1 vccd1 vccd1 hold4465/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4476 _10108_/X vssd1 vssd1 vccd1 vccd1 _16526_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3731 _10498_/X vssd1 vssd1 vccd1 vccd1 _16656_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3742 _16613_/Q vssd1 vssd1 vccd1 vccd1 hold3742/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4487 _12560_/X vssd1 vssd1 vccd1 vccd1 _12561_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3753 _16624_/Q vssd1 vssd1 vccd1 vccd1 hold3753/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4498 _17574_/Q vssd1 vssd1 vccd1 vccd1 hold4498/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3764 _13342_/X vssd1 vssd1 vccd1 vccd1 _17567_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3775 _16647_/Q vssd1 vssd1 vccd1 vccd1 hold3775/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3786 _10351_/X vssd1 vssd1 vccd1 vccd1 _16607_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3797 _16325_/Q vssd1 vssd1 vccd1 vccd1 _13070_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09709_ hold3746/X _10013_/B _09708_/X _15042_/A vssd1 vssd1 vccd1 vccd1 _09709_/X
+ sky130_fd_sc_hd__o211a_1
X_10981_ hold4997/X _11165_/B _10980_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _10981_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12720_ _12810_/A _12720_/B vssd1 vssd1 vccd1 vccd1 _17416_/D sky130_fd_sc_hd__and2_1
XFILLER_0_214_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12651_ _12849_/A _12651_/B vssd1 vssd1 vccd1 vccd1 _17393_/D sky130_fd_sc_hd__and2_1
XFILLER_0_214_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ hold5400/X _12335_/B _11601_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _11602_/X
+ sky130_fd_sc_hd__o211a_1
X_15370_ hold722/X _15448_/A2 _15446_/B1 hold561/X vssd1 vssd1 vccd1 vccd1 _15370_/X
+ sky130_fd_sc_hd__a22o_1
X_12582_ _12894_/A _12582_/B vssd1 vssd1 vccd1 vccd1 _17370_/D sky130_fd_sc_hd__and2_1
XFILLER_0_66_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14321_ hold2850/X _14326_/B _14320_/Y _14344_/A vssd1 vssd1 vccd1 vccd1 _14321_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11533_ hold5374/X _11726_/B _11532_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _11533_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_381_wb_clk_i clkbuf_6_33_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17262_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17040_ _17885_/CLK _17040_/D vssd1 vssd1 vccd1 vccd1 _17040_/Q sky130_fd_sc_hd__dfxtp_1
X_14252_ _14413_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14252_/X sky130_fd_sc_hd__or2_1
X_11464_ hold5111/X _11753_/B _11463_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _11464_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_310_wb_clk_i clkbuf_6_45_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17973_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10415_ hold2064/X hold3345/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10416_/B sky130_fd_sc_hd__mux2_1
X_13203_ _13202_/X _16918_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13203_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11395_ hold5349/X _12323_/B _11394_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _11395_/X
+ sky130_fd_sc_hd__o211a_1
X_14183_ hold3006/X _14202_/B _14182_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _14183_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13134_ _13134_/A _13294_/B vssd1 vssd1 vccd1 vccd1 _13134_/X sky130_fd_sc_hd__or2_1
X_10346_ hold2493/X hold4493/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10347_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_238_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _13065_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13065_/X sky130_fd_sc_hd__and2_1
XFILLER_0_209_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17942_ _18061_/CLK _17942_/D vssd1 vssd1 vccd1 vccd1 _17942_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10277_ hold3082/X _16583_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10278_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12016_ hold4827/X _12293_/B _12015_/X _12103_/C1 vssd1 vssd1 vccd1 vccd1 _12016_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_218_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17873_ _17873_/CLK _17873_/D vssd1 vssd1 vccd1 vccd1 _17873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16824_ _18059_/CLK _16824_/D vssd1 vssd1 vccd1 vccd1 _16824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16755_ _17967_/CLK _16755_/D vssd1 vssd1 vccd1 vccd1 _16755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13967_ hold1787/X _13995_/A2 _13966_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _13967_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_232_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15706_ _17576_/CLK _15706_/D vssd1 vssd1 vccd1 vccd1 _15706_/Q sky130_fd_sc_hd__dfxtp_1
X_12918_ _12924_/A _12918_/B vssd1 vssd1 vccd1 vccd1 _17482_/D sky130_fd_sc_hd__and2_1
X_16686_ _18212_/CLK _16686_/D vssd1 vssd1 vccd1 vccd1 _16686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13898_ _15513_/A hold2903/X hold297/X vssd1 vssd1 vccd1 vccd1 _13899_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18425_ _18425_/CLK _18425_/D vssd1 vssd1 vccd1 vccd1 _18425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15637_ _17266_/CLK _15637_/D vssd1 vssd1 vccd1 vccd1 _15637_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _12849_/A _12849_/B vssd1 vssd1 vccd1 vccd1 _17459_/D sky130_fd_sc_hd__and2_1
XFILLER_0_158_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18356_ _18356_/CLK _18356_/D vssd1 vssd1 vccd1 vccd1 _18356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ _17236_/CLK _15568_/D vssd1 vssd1 vccd1 vccd1 _15568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17307_ _17331_/CLK _17307_/D vssd1 vssd1 vccd1 vccd1 hold126/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14519_ _15199_/A _14543_/B vssd1 vssd1 vccd1 vccd1 _14519_/X sky130_fd_sc_hd__or2_1
XFILLER_0_56_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18287_ _18325_/CLK _18287_/D vssd1 vssd1 vccd1 vccd1 _18287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15499_ _15515_/A hold2223/X _15505_/S vssd1 vssd1 vccd1 vccd1 _15500_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_182_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08040_ hold2775/X _08033_/B _08039_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _08040_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17238_ _17898_/CLK _17238_/D vssd1 vssd1 vccd1 vccd1 _17238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold903 hold903/A vssd1 vssd1 vccd1 vccd1 hold903/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold914 hold914/A vssd1 vssd1 vccd1 vccd1 hold914/X sky130_fd_sc_hd__clkbuf_2
X_17169_ _17902_/CLK _17169_/D vssd1 vssd1 vccd1 vccd1 _17169_/Q sky130_fd_sc_hd__dfxtp_1
Xhold925 hold925/A vssd1 vssd1 vccd1 vccd1 hold925/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 hold936/A vssd1 vssd1 vccd1 vccd1 hold936/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold947 hold947/A vssd1 vssd1 vccd1 vccd1 hold947/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 hold958/A vssd1 vssd1 vccd1 vccd1 hold958/X sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ _11203_/A _09991_/B vssd1 vssd1 vccd1 vccd1 _09991_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_161_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold969 hold969/A vssd1 vssd1 vccd1 vccd1 hold969/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3005 _09197_/X vssd1 vssd1 vccd1 vccd1 _16210_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3016 _15810_/Q vssd1 vssd1 vccd1 vccd1 hold3016/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3027 _15609_/Q vssd1 vssd1 vccd1 vccd1 hold3027/X sky130_fd_sc_hd__dlygate4sd3_1
X_08942_ _15344_/A hold685/X vssd1 vssd1 vccd1 vccd1 _16088_/D sky130_fd_sc_hd__and2_1
XFILLER_0_23_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3038 _09151_/X vssd1 vssd1 vccd1 vccd1 _16188_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2304 _15741_/Q vssd1 vssd1 vccd1 vccd1 hold2304/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3049 _17862_/Q vssd1 vssd1 vccd1 vccd1 hold3049/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2315 _14538_/X vssd1 vssd1 vccd1 vccd1 _18065_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2326 _15795_/Q vssd1 vssd1 vccd1 vccd1 hold2326/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2337 _16234_/Q vssd1 vssd1 vccd1 vccd1 hold2337/X sky130_fd_sc_hd__dlygate4sd3_1
X_08873_ _15414_/A hold798/X vssd1 vssd1 vccd1 vccd1 _16054_/D sky130_fd_sc_hd__and2_1
Xhold2348 _14269_/X vssd1 vssd1 vccd1 vccd1 _17935_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1603 _07929_/X vssd1 vssd1 vccd1 vccd1 _15608_/D sky130_fd_sc_hd__dlygate4sd3_1
Xload_slew861 _09498_/A vssd1 vssd1 vccd1 vccd1 _14681_/A sky130_fd_sc_hd__buf_6
XFILLER_0_208_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1614 _16227_/Q vssd1 vssd1 vccd1 vccd1 hold1614/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2359 _15684_/Q vssd1 vssd1 vccd1 vccd1 hold2359/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1625 _15116_/X vssd1 vssd1 vccd1 vccd1 _18342_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07824_ _09366_/A _09122_/A _07824_/C _09121_/B vssd1 vssd1 vccd1 vccd1 _07824_/Y
+ sky130_fd_sc_hd__nor4_2
Xhold1636 _13010_/X vssd1 vssd1 vccd1 vccd1 _17513_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1647 hold6120/X vssd1 vssd1 vccd1 vccd1 hold1647/X sky130_fd_sc_hd__buf_1
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1658 _17788_/Q vssd1 vssd1 vccd1 vccd1 hold1658/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1669 _15803_/Q vssd1 vssd1 vccd1 vccd1 hold1669/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09425_ _07804_/A _09472_/C _15274_/A _09424_/X vssd1 vssd1 vccd1 vccd1 _09425_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09356_ _09366_/A _09366_/B _09356_/C vssd1 vssd1 vccd1 vccd1 _09356_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_139_wb_clk_i clkbuf_6_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18419_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08307_ _15531_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08307_/X sky130_fd_sc_hd__or2_1
X_09287_ hold927/X _09337_/B vssd1 vssd1 vccd1 vccd1 _09287_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08238_ _14457_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08238_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08169_ _15502_/A _08169_/B vssd1 vssd1 vccd1 vccd1 _15722_/D sky130_fd_sc_hd__and2_1
XFILLER_0_127_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10200_ _10524_/A _10200_/B vssd1 vssd1 vccd1 vccd1 _10200_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11180_ _16884_/Q _11186_/B _11186_/C vssd1 vssd1 vccd1 vccd1 _11180_/X sky130_fd_sc_hd__and3_1
XFILLER_0_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4240 _13830_/Y vssd1 vssd1 vccd1 vccd1 _13831_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10131_ _10515_/A _10131_/B vssd1 vssd1 vccd1 vccd1 _10131_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4251 _16721_/Q vssd1 vssd1 vccd1 vccd1 hold4251/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4262 _17568_/Q vssd1 vssd1 vccd1 vccd1 hold4262/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4273 _17115_/Q vssd1 vssd1 vccd1 vccd1 hold4273/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4284 _16718_/Q vssd1 vssd1 vccd1 vccd1 hold4284/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3550 _16581_/Q vssd1 vssd1 vccd1 vccd1 hold3550/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4295 _16930_/Q vssd1 vssd1 vccd1 vccd1 hold4295/X sky130_fd_sc_hd__dlygate4sd3_1
X_10062_ _13278_/A _10482_/A _10061_/X vssd1 vssd1 vccd1 vccd1 _10062_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3561 _09547_/X vssd1 vssd1 vccd1 vccd1 _16339_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3572 _16389_/Q vssd1 vssd1 vccd1 vccd1 hold3572/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3583 _09859_/X vssd1 vssd1 vccd1 vccd1 _16443_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3594 _10381_/X vssd1 vssd1 vccd1 vccd1 _16617_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2860 _07961_/X vssd1 vssd1 vccd1 vccd1 _15623_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14870_ _15209_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14870_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2871 _17850_/Q vssd1 vssd1 vccd1 vccd1 hold2871/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2882 _15516_/X vssd1 vssd1 vccd1 vccd1 _18436_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2893 _15766_/Q vssd1 vssd1 vccd1 vccd1 hold2893/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13821_ hold4242/X _13734_/A _13820_/X vssd1 vssd1 vccd1 vccd1 _13821_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_230_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_214_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16540_ _18162_/CLK _16540_/D vssd1 vssd1 vccd1 vccd1 _16540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13752_ _13752_/A _13752_/B vssd1 vssd1 vccd1 vccd1 _13752_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10964_ hold2613/X _16812_/Q _10964_/S vssd1 vssd1 vccd1 vccd1 _10965_/B sky130_fd_sc_hd__mux2_1
X_12703_ hold2284/X hold3722/X _12766_/S vssd1 vssd1 vccd1 vccd1 _12703_/X sky130_fd_sc_hd__mux2_1
X_16471_ _18384_/CLK _16471_/D vssd1 vssd1 vccd1 vccd1 _16471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13683_ _13758_/A _13683_/B vssd1 vssd1 vccd1 vccd1 _13683_/X sky130_fd_sc_hd__or2_1
X_10895_ hold2511/X _16789_/Q _11183_/C vssd1 vssd1 vccd1 vccd1 _10896_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18210_ _18210_/CLK _18210_/D vssd1 vssd1 vccd1 vccd1 _18210_/Q sky130_fd_sc_hd__dfxtp_1
X_15422_ _15480_/A _15422_/B _15422_/C _15422_/D vssd1 vssd1 vccd1 vccd1 _15422_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_39_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12634_ hold1414/X _17389_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12634_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18141_ _18205_/CLK _18141_/D vssd1 vssd1 vccd1 vccd1 _18141_/Q sky130_fd_sc_hd__dfxtp_1
X_15353_ _15481_/A1 _15345_/X _15352_/X _15481_/B1 hold4185/X vssd1 vssd1 vccd1 vccd1
+ _15353_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_38_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12565_ hold2767/X _17366_/Q _12985_/S vssd1 vssd1 vccd1 vccd1 _12565_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14304_ _15199_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14304_/X sky130_fd_sc_hd__or2_1
X_18072_ _18072_/CLK _18072_/D vssd1 vssd1 vccd1 vccd1 _18072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11516_ hold1258/X hold4050/X _12317_/C vssd1 vssd1 vccd1 vccd1 _11517_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15284_ _15284_/A _15284_/B vssd1 vssd1 vccd1 vccd1 _18404_/D sky130_fd_sc_hd__and2_1
Xclkbuf_6_16_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_16_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12496_ _17341_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12496_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17023_ _17871_/CLK _17023_/D vssd1 vssd1 vccd1 vccd1 _17023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14235_ hold2165/X _14268_/B _14234_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _14235_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11447_ hold2121/X _16973_/Q _11738_/C vssd1 vssd1 vccd1 vccd1 _11448_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14166_ _14166_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14166_/X sky130_fd_sc_hd__or2_1
X_11378_ hold2312/X _16950_/Q _11660_/S vssd1 vssd1 vccd1 vccd1 _11379_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13117_ _13116_/X hold3423/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13117_/X sky130_fd_sc_hd__mux2_1
X_10329_ _11088_/A _10329_/B vssd1 vssd1 vccd1 vccd1 _10329_/X sky130_fd_sc_hd__or2_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ hold2071/X _14107_/A2 _14096_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _14097_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13048_ _13048_/A _13048_/B vssd1 vssd1 vccd1 vccd1 _13048_/X sky130_fd_sc_hd__and2_1
X_17925_ _18020_/CLK _17925_/D vssd1 vssd1 vccd1 vccd1 _17925_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_234_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17856_ _17856_/CLK hold710/X vssd1 vssd1 vccd1 vccd1 _17856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16807_ _18042_/CLK _16807_/D vssd1 vssd1 vccd1 vccd1 _16807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17787_ _17883_/CLK _17787_/D vssd1 vssd1 vccd1 vccd1 _17787_/Q sky130_fd_sc_hd__dfxtp_1
X_14999_ hold1891/X hold447/X _14998_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _14999_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_178_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16738_ _18005_/CLK _16738_/D vssd1 vssd1 vccd1 vccd1 _16738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16669_ _18227_/CLK _16669_/D vssd1 vssd1 vccd1 vccd1 _16669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_6_55_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_55_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_202_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09210_ _15539_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09210_/X sky130_fd_sc_hd__or2_1
X_18408_ _18408_/CLK _18408_/D vssd1 vssd1 vccd1 vccd1 _18408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_232_wb_clk_i clkbuf_6_62_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18233_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_118_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ hold1186/X _09177_/A2 _09140_/X _12873_/A vssd1 vssd1 vccd1 vccd1 _09141_/X
+ sky130_fd_sc_hd__o211a_1
X_18339_ _18371_/CLK _18339_/D vssd1 vssd1 vccd1 vccd1 _18339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09072_ _14972_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09072_/X sky130_fd_sc_hd__or2_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08023_ _15537_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08023_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold700 hold700/A vssd1 vssd1 vccd1 vccd1 hold700/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 slv_done vssd1 vssd1 vccd1 vccd1 hold711/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold722 hold722/A vssd1 vssd1 vccd1 vccd1 hold722/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 hold733/A vssd1 vssd1 vccd1 vccd1 hold733/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold744 hold744/A vssd1 vssd1 vccd1 vccd1 hold744/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold755 hold755/A vssd1 vssd1 vccd1 vccd1 hold755/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold766 hold766/A vssd1 vssd1 vccd1 vccd1 hold766/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 hold777/A vssd1 vssd1 vccd1 vccd1 hold777/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold788 hold788/A vssd1 vssd1 vccd1 vccd1 hold788/X sky130_fd_sc_hd__buf_1
Xhold799 hold799/A vssd1 vssd1 vccd1 vccd1 hold799/X sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ hold1805/X _16482_/Q _10040_/C vssd1 vssd1 vccd1 vccd1 _09975_/B sky130_fd_sc_hd__mux2_1
Xhold2101 _14767_/X vssd1 vssd1 vccd1 vccd1 _18174_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2112 _14763_/X vssd1 vssd1 vccd1 vccd1 _18172_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08925_ _15284_/A hold469/X vssd1 vssd1 vccd1 vccd1 _16080_/D sky130_fd_sc_hd__and2_1
Xhold2123 _17880_/Q vssd1 vssd1 vccd1 vccd1 hold2123/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2134 _14504_/X vssd1 vssd1 vccd1 vccd1 _18048_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1400 _16265_/Q vssd1 vssd1 vccd1 vccd1 hold1400/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2145 _16268_/Q vssd1 vssd1 vccd1 vccd1 hold2145/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1411 _15704_/Q vssd1 vssd1 vccd1 vccd1 hold1411/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2156 _15536_/X vssd1 vssd1 vccd1 vccd1 _18446_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1422 _18427_/Q vssd1 vssd1 vccd1 vccd1 hold1422/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2167 _17872_/Q vssd1 vssd1 vccd1 vccd1 hold2167/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1433 _15005_/X vssd1 vssd1 vccd1 vccd1 _18288_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08856_ hold315/X hold346/X _08866_/S vssd1 vssd1 vccd1 vccd1 _08857_/B sky130_fd_sc_hd__mux2_1
Xhold2178 _14899_/X vssd1 vssd1 vccd1 vccd1 _18237_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1444 _16315_/Q vssd1 vssd1 vccd1 vccd1 _09463_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2189 _17847_/Q vssd1 vssd1 vccd1 vccd1 hold2189/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1455 _18118_/Q vssd1 vssd1 vccd1 vccd1 hold1455/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1466 _15087_/X vssd1 vssd1 vccd1 vccd1 hold1466/X sky130_fd_sc_hd__dlygate4sd3_1
X_07807_ _07785_/Y _07789_/A _07805_/A _07806_/Y vssd1 vssd1 vccd1 vccd1 _07807_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1477 _18433_/Q vssd1 vssd1 vccd1 vccd1 hold1477/X sky130_fd_sc_hd__dlygate4sd3_1
X_08787_ hold87/X hold463/X _08793_/S vssd1 vssd1 vccd1 vccd1 hold464/A sky130_fd_sc_hd__mux2_1
Xhold1488 _14470_/X vssd1 vssd1 vccd1 vccd1 _18032_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 _16277_/Q vssd1 vssd1 vccd1 vccd1 hold1499/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09408_ _09438_/B _16290_/Q vssd1 vssd1 vccd1 vccd1 _09408_/X sky130_fd_sc_hd__or2_1
X_10680_ _11067_/A _10680_/B vssd1 vssd1 vccd1 vccd1 _10680_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09339_ _09339_/A _09339_/B vssd1 vssd1 vccd1 vccd1 _09339_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12350_ _17274_/Q _12350_/B _13463_/S vssd1 vssd1 vccd1 vccd1 _12350_/X sky130_fd_sc_hd__and3_1
XFILLER_0_50_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11301_ _11553_/A _11301_/B vssd1 vssd1 vccd1 vccd1 _11301_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12281_ hold2714/X hold5255/X _13886_/C vssd1 vssd1 vccd1 vccd1 _12282_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_160_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14020_ hold951/X _14042_/B vssd1 vssd1 vccd1 vccd1 _14020_/X sky130_fd_sc_hd__or2_1
X_11232_ _12093_/A _11232_/B vssd1 vssd1 vccd1 vccd1 _11232_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_1377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11163_ hold4284/X _11010_/A _11162_/X vssd1 vssd1 vccd1 vccd1 _11163_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_36_wb_clk_i clkbuf_6_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17847_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4070 _16766_/Q vssd1 vssd1 vccd1 vccd1 hold4070/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10114_ hold3684/X _10598_/B _10113_/X _15218_/C1 vssd1 vssd1 vccd1 vccd1 _10114_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4081 _16798_/Q vssd1 vssd1 vccd1 vccd1 hold4081/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15971_ _17309_/CLK _15971_/D vssd1 vssd1 vccd1 vccd1 hold263/A sky130_fd_sc_hd__dfxtp_1
X_11094_ _11121_/A _11094_/B vssd1 vssd1 vccd1 vccd1 _11094_/X sky130_fd_sc_hd__or2_1
Xhold4092 _11233_/X vssd1 vssd1 vccd1 vccd1 _16901_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17710_ _17742_/CLK _17710_/D vssd1 vssd1 vccd1 vccd1 _17710_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3380 _17449_/Q vssd1 vssd1 vccd1 vccd1 hold3380/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10045_ _10603_/A _10045_/B vssd1 vssd1 vccd1 vccd1 _16505_/D sky130_fd_sc_hd__nor2_1
XTAP_6298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14922_ _15191_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14922_/X sky130_fd_sc_hd__or2_1
XTAP_5553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3391 _12830_/X vssd1 vssd1 vccd1 vccd1 _12831_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__buf_4
XTAP_5586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__buf_4
Xhold2690 _14665_/X vssd1 vssd1 vccd1 vccd1 _18125_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17641_ _17737_/CLK _17641_/D vssd1 vssd1 vccd1 vccd1 _17641_/Q sky130_fd_sc_hd__dfxtp_1
X_14853_ hold2483/X _14880_/B _14852_/X _14853_/C1 vssd1 vssd1 vccd1 vccd1 _14853_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_230_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _13819_/A _13804_/B vssd1 vssd1 vccd1 vccd1 _13804_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_76_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17572_ _17648_/CLK _17572_/D vssd1 vssd1 vccd1 vccd1 _17572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14784_ _15231_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14784_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11996_ hold1346/X hold4596/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11997_/B sky130_fd_sc_hd__mux2_1
X_16523_ _18081_/CLK _16523_/D vssd1 vssd1 vccd1 vccd1 _16523_/Q sky130_fd_sc_hd__dfxtp_1
X_13735_ hold4624/X _13829_/B _13734_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13735_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10947_ _11637_/A _10947_/B vssd1 vssd1 vccd1 vccd1 _10947_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16454_ _18271_/CLK _16454_/D vssd1 vssd1 vccd1 vccd1 _16454_/Q sky130_fd_sc_hd__dfxtp_1
X_13666_ hold5386/X _13856_/B _13665_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13666_/X
+ sky130_fd_sc_hd__o211a_1
X_10878_ _11655_/A _10878_/B vssd1 vssd1 vccd1 vccd1 _10878_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15405_ hold574/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15405_/X sky130_fd_sc_hd__or2_1
XFILLER_0_13_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12617_ _17382_/Q _12616_/X _12626_/S vssd1 vssd1 vccd1 vccd1 _12617_/X sky130_fd_sc_hd__mux2_1
X_16385_ _18298_/CLK _16385_/D vssd1 vssd1 vccd1 vccd1 _16385_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13597_ hold5494/X _13883_/B _13596_/X _08347_/A vssd1 vssd1 vccd1 vccd1 _13597_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18124_ _18124_/CLK _18124_/D vssd1 vssd1 vccd1 vccd1 _18124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15336_ _17337_/Q _15486_/B1 _09362_/D hold502/X vssd1 vssd1 vccd1 vccd1 _15336_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12548_ hold3381/X _12547_/X _12923_/S vssd1 vssd1 vccd1 vccd1 _12548_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18055_ _18063_/CLK _18055_/D vssd1 vssd1 vccd1 vccd1 _18055_/Q sky130_fd_sc_hd__dfxtp_1
X_15267_ hold760/X _09357_/A _09386_/D hold514/X _15266_/X vssd1 vssd1 vccd1 vccd1
+ _15272_/B sky130_fd_sc_hd__a221o_1
X_12479_ hold185/X _12445_/A _12445_/B _12478_/X _09057_/A vssd1 vssd1 vccd1 vccd1
+ hold15/A sky130_fd_sc_hd__o311a_1
XANTENNA_2 _13068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17006_ _17886_/CLK _17006_/D vssd1 vssd1 vccd1 vccd1 _17006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14218_ hold927/X _14230_/B vssd1 vssd1 vccd1 vccd1 _14218_/X sky130_fd_sc_hd__or2_1
X_15198_ hold1002/X _15221_/B _15197_/X _15048_/A vssd1 vssd1 vccd1 vccd1 _15198_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14149_ hold2460/X _14148_/B _14148_/Y _15494_/A vssd1 vssd1 vccd1 vccd1 _14149_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout509 _09499_/Y vssd1 vssd1 vccd1 vccd1 _10538_/S sky130_fd_sc_hd__buf_4
XFILLER_0_238_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08710_ _12412_/A _08710_/B vssd1 vssd1 vccd1 vccd1 _15976_/D sky130_fd_sc_hd__and2_1
X_17908_ _17908_/CLK _17908_/D vssd1 vssd1 vccd1 vccd1 _17908_/Q sky130_fd_sc_hd__dfxtp_1
X_09690_ _10482_/A _09690_/B vssd1 vssd1 vccd1 vccd1 _09690_/X sky130_fd_sc_hd__or2_1
XFILLER_0_241_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08641_ hold373/X hold497/X _08657_/S vssd1 vssd1 vccd1 vccd1 _08642_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_174_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17839_ _17871_/CLK _17839_/D vssd1 vssd1 vccd1 vccd1 _17839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08572_ hold5/X hold639/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08573_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_178_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_413_wb_clk_i clkbuf_6_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17856_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09124_ _15128_/A hold363/A vssd1 vssd1 vccd1 vccd1 _09124_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_165_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09055_ _12440_/A hold397/X vssd1 vssd1 vccd1 vccd1 _16144_/D sky130_fd_sc_hd__and2_1
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08006_ hold1346/X _08029_/B _08005_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _08006_/X
+ sky130_fd_sc_hd__o211a_1
Xhold530 hold530/A vssd1 vssd1 vccd1 vccd1 hold530/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold541 hold541/A vssd1 vssd1 vccd1 vccd1 hold541/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold552 hold594/X vssd1 vssd1 vccd1 vccd1 hold595/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 hold563/A vssd1 vssd1 vccd1 vccd1 hold563/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold574 hold574/A vssd1 vssd1 vccd1 vccd1 hold574/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold585 hold585/A vssd1 vssd1 vccd1 vccd1 hold585/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold596 input45/X vssd1 vssd1 vccd1 vccd1 hold596/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09957_ _09957_/A _09957_/B vssd1 vssd1 vccd1 vccd1 _09957_/X sky130_fd_sc_hd__or2_1
XFILLER_0_99_1256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08908_ hold215/X hold532/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08909_/B sky130_fd_sc_hd__mux2_1
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09888_ _09912_/A _09888_/B vssd1 vssd1 vccd1 vccd1 _09888_/X sky130_fd_sc_hd__or2_1
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1230 _08014_/X vssd1 vssd1 vccd1 vccd1 _15648_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1241 _15716_/Q vssd1 vssd1 vccd1 vccd1 hold1241/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1252 input43/X vssd1 vssd1 vccd1 vccd1 hold641/A sky130_fd_sc_hd__buf_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08839_ _12394_/A _08839_/B vssd1 vssd1 vccd1 vccd1 _16038_/D sky130_fd_sc_hd__and2_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1263 _15817_/Q vssd1 vssd1 vccd1 vccd1 hold1263/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1274 _14185_/X vssd1 vssd1 vccd1 vccd1 _17895_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_234_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1285 _17906_/Q vssd1 vssd1 vccd1 vccd1 hold1285/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1296 _14518_/X vssd1 vssd1 vccd1 vccd1 _18055_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _12234_/A _11850_/B vssd1 vssd1 vccd1 vccd1 _11850_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_154_wb_clk_i clkbuf_6_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18418_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10801_ hold5267/X _10616_/B _10800_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _10801_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ hold4405/X _12219_/A _11780_/X vssd1 vssd1 vccd1 vccd1 _11781_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13520_ hold2541/X _17627_/Q _13817_/C vssd1 vssd1 vccd1 vccd1 _13521_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10732_ hold4070/X _11210_/B _10731_/X _14528_/C1 vssd1 vssd1 vccd1 vccd1 _10732_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13451_ hold1548/X hold5034/X _13871_/C vssd1 vssd1 vccd1 vccd1 _13452_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10663_ hold3872/X _11144_/B _10662_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _10663_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12402_ _15344_/A _12402_/B vssd1 vssd1 vccd1 vccd1 _17294_/D sky130_fd_sc_hd__and2_1
XFILLER_0_180_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16170_ _17506_/CLK _16170_/D vssd1 vssd1 vccd1 vccd1 _16170_/Q sky130_fd_sc_hd__dfxtp_1
X_10594_ _11206_/A _10594_/B vssd1 vssd1 vccd1 vccd1 _16688_/D sky130_fd_sc_hd__nor2_1
X_13382_ hold2895/X hold4293/X _13481_/S vssd1 vssd1 vccd1 vccd1 _13383_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15121_ _15229_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15121_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12333_ hold4248/X _12159_/A _12332_/X vssd1 vssd1 vccd1 vccd1 _12333_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_181_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15052_ _15054_/A _15052_/B vssd1 vssd1 vccd1 vccd1 _18311_/D sky130_fd_sc_hd__and2_1
XFILLER_0_142_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12264_ _12267_/A _12264_/B vssd1 vssd1 vccd1 vccd1 _12264_/X sky130_fd_sc_hd__or2_1
X_14003_ hold1970/X _14040_/B _14002_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _14003_/X
+ sky130_fd_sc_hd__o211a_1
X_11215_ _11218_/A _11215_/B vssd1 vssd1 vccd1 vccd1 _11215_/Y sky130_fd_sc_hd__nor2_1
X_12195_ _13797_/A _12195_/B vssd1 vssd1 vccd1 vccd1 _12195_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput72 _13051_/A vssd1 vssd1 vccd1 vccd1 output72/X sky130_fd_sc_hd__buf_6
Xoutput83 _13065_/A vssd1 vssd1 vccd1 vccd1 output83/X sky130_fd_sc_hd__buf_6
XTAP_6040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ _11158_/A _11146_/B vssd1 vssd1 vccd1 vccd1 _16872_/D sky130_fd_sc_hd__nor2_1
Xoutput94 _13073_/A vssd1 vssd1 vccd1 vccd1 output94/X sky130_fd_sc_hd__buf_6
XTAP_6051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15954_ _17301_/CLK _15954_/D vssd1 vssd1 vccd1 vccd1 hold743/A sky130_fd_sc_hd__dfxtp_1
X_11077_ hold5038/X _11165_/B _11076_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _11077_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14905_ hold1779/X _14896_/Y _14904_/X _15482_/A vssd1 vssd1 vccd1 vccd1 _14905_/X
+ sky130_fd_sc_hd__o211a_1
X_10028_ _16500_/Q _10028_/B _10028_/C vssd1 vssd1 vccd1 vccd1 _10028_/X sky130_fd_sc_hd__and3_1
XTAP_5394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15885_ _17561_/CLK _15885_/D vssd1 vssd1 vccd1 vccd1 _15885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14836_ _15229_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14836_/X sky130_fd_sc_hd__or2_1
X_17624_ _17624_/CLK _17624_/D vssd1 vssd1 vccd1 vccd1 _17624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17555_ _18229_/CLK _17555_/D vssd1 vssd1 vccd1 vccd1 _17555_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14767_ hold2100/X _14772_/B _14766_/X _14769_/C1 vssd1 vssd1 vccd1 vccd1 _14767_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11979_ _12267_/A _11979_/B vssd1 vssd1 vccd1 vccd1 _11979_/X sky130_fd_sc_hd__or2_1
XFILLER_0_188_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16506_ _18387_/CLK _16506_/D vssd1 vssd1 vccd1 vccd1 _16506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13718_ hold1267/X hold5777/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13719_/B sky130_fd_sc_hd__mux2_1
X_17486_ _17486_/CLK _17486_/D vssd1 vssd1 vccd1 vccd1 _17486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14698_ _15199_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14698_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16437_ _18382_/CLK _16437_/D vssd1 vssd1 vccd1 vccd1 _16437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13649_ hold1744/X _17670_/Q _13841_/C vssd1 vssd1 vccd1 vccd1 _13650_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_229_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16368_ _18315_/CLK _16368_/D vssd1 vssd1 vccd1 vccd1 _16368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18107_ _18262_/CLK _18107_/D vssd1 vssd1 vccd1 vccd1 _18107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15319_ hold638/X _15485_/A2 _15488_/A2 hold590/X _15318_/X vssd1 vssd1 vccd1 vccd1
+ _15322_/C sky130_fd_sc_hd__a221o_1
Xhold5507 _17620_/Q vssd1 vssd1 vccd1 vccd1 hold5507/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16299_ _18460_/CLK hold740/X vssd1 vssd1 vccd1 vccd1 _16299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5518 _11344_/X vssd1 vssd1 vccd1 vccd1 _16938_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5529 _17020_/Q vssd1 vssd1 vccd1 vccd1 hold5529/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18038_ _18070_/CLK _18038_/D vssd1 vssd1 vccd1 vccd1 _18038_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4806 _11818_/X vssd1 vssd1 vccd1 vccd1 _17096_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4817 _16834_/Q vssd1 vssd1 vccd1 vccd1 hold4817/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4828 _12016_/X vssd1 vssd1 vccd1 vccd1 _17162_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4839 _16434_/Q vssd1 vssd1 vccd1 vccd1 hold4839/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout306 _11061_/A vssd1 vssd1 vccd1 vccd1 _11106_/A sky130_fd_sc_hd__buf_4
XFILLER_0_22_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09811_ hold3576/X _10025_/B _09810_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09811_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_201_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout317 _11088_/A vssd1 vssd1 vccd1 vccd1 _11103_/A sky130_fd_sc_hd__buf_4
Xfanout328 _10386_/A vssd1 vssd1 vccd1 vccd1 _10482_/A sky130_fd_sc_hd__buf_4
Xfanout339 _12508_/B vssd1 vssd1 vccd1 vccd1 _12506_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09742_ hold4581/X _10028_/B _09741_/X _15048_/A vssd1 vssd1 vccd1 vccd1 _09742_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_236_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09673_ hold3617/X _10049_/B _09672_/X _15212_/C1 vssd1 vssd1 vccd1 vccd1 _09673_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _15364_/A hold752/X vssd1 vssd1 vccd1 vccd1 _15934_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _15434_/A hold282/X vssd1 vssd1 vccd1 vccd1 _15901_/D sky130_fd_sc_hd__and2_1
XFILLER_0_204_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08486_ _15545_/A _08486_/B vssd1 vssd1 vccd1 vccd1 _08486_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_37_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09107_ hold2468/X _09102_/B _09106_/Y _12987_/A vssd1 vssd1 vccd1 vccd1 _09107_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09038_ hold215/X hold301/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09039_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_14_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold360 input61/X vssd1 vssd1 vccd1 vccd1 hold360/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_104_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold371 hold46/X vssd1 vssd1 vccd1 vccd1 input18/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 hold382/A vssd1 vssd1 vccd1 vccd1 input44/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 hold393/A vssd1 vssd1 vccd1 vccd1 input32/A sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ hold2601/X hold4959/X _11660_/S vssd1 vssd1 vccd1 vccd1 _11001_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_229_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout840 _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14881_/C1 sky130_fd_sc_hd__buf_4
Xfanout851 _11203_/A vssd1 vssd1 vccd1 vccd1 _11158_/A sky130_fd_sc_hd__buf_6
Xfanout862 _07785_/Y vssd1 vssd1 vccd1 vccd1 _07804_/A sky130_fd_sc_hd__clkbuf_8
Xfanout873 _14952_/A vssd1 vssd1 vccd1 vccd1 _15221_/A sky130_fd_sc_hd__buf_12
Xfanout884 hold932/X vssd1 vssd1 vccd1 vccd1 _15197_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_335_wb_clk_i clkbuf_6_43_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17187_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_102_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout895 hold944/X vssd1 vssd1 vccd1 vccd1 hold945/A sky130_fd_sc_hd__buf_6
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _12984_/A _12951_/B vssd1 vssd1 vccd1 vccd1 _17493_/D sky130_fd_sc_hd__and2_1
XFILLER_0_198_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1060 _18230_/Q vssd1 vssd1 vccd1 vccd1 hold1060/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1071 _14125_/X vssd1 vssd1 vccd1 vccd1 _17866_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11902_ hold4596/X _12308_/B _11901_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _11902_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1082 _15594_/Q vssd1 vssd1 vccd1 vccd1 hold1082/X sky130_fd_sc_hd__dlygate4sd3_1
X_15670_ _17127_/CLK _15670_/D vssd1 vssd1 vccd1 vccd1 _15670_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1093 _17778_/Q vssd1 vssd1 vccd1 vccd1 hold1093/X sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ _12888_/A _12882_/B vssd1 vssd1 vccd1 vccd1 _17470_/D sky130_fd_sc_hd__and2_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ hold2652/X _14612_/B _14620_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14621_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11833_ hold5022/X _12217_/A2 _11832_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _11833_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17340_ _17344_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 _17340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ hold1893/X _14537_/B _14551_/X _14552_/C1 vssd1 vssd1 vccd1 vccd1 _14552_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _12331_/A _11764_/B vssd1 vssd1 vccd1 vccd1 _11764_/Y sky130_fd_sc_hd__nor2_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13503_ _13599_/A _13503_/B vssd1 vssd1 vccd1 vccd1 _13503_/X sky130_fd_sc_hd__or2_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _17271_/CLK _17271_/D vssd1 vssd1 vccd1 vccd1 _17271_/Q sky130_fd_sc_hd__dfxtp_1
X_10715_ hold2004/X hold3590/X _11210_/C vssd1 vssd1 vccd1 vccd1 _10716_/B sky130_fd_sc_hd__mux2_1
X_14483_ _15217_/A _14487_/B vssd1 vssd1 vccd1 vccd1 _14483_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_193_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11695_ hold5311/X _11789_/B _11694_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _11695_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16222_ _17452_/CLK _16222_/D vssd1 vssd1 vccd1 vccd1 _16222_/Q sky130_fd_sc_hd__dfxtp_1
X_13434_ _13794_/A _13434_/B vssd1 vssd1 vccd1 vccd1 _13434_/X sky130_fd_sc_hd__or2_1
X_10646_ _16706_/Q _10646_/B _10646_/C vssd1 vssd1 vccd1 vccd1 _10646_/X sky130_fd_sc_hd__and3_1
XFILLER_0_3_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16153_ _17492_/CLK _16153_/D vssd1 vssd1 vccd1 vccd1 _16153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13365_ _13407_/A _13365_/B vssd1 vssd1 vccd1 vccd1 _13365_/X sky130_fd_sc_hd__or2_1
X_10577_ _16683_/Q _10577_/B _10601_/C vssd1 vssd1 vccd1 vccd1 _10577_/X sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_51_wb_clk_i clkbuf_6_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18039_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_210_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15104_ hold1789/X hold341/X _15103_/X _08954_/A vssd1 vssd1 vccd1 vccd1 _15104_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ _13819_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _12316_/Y sky130_fd_sc_hd__nor2_1
X_16084_ _18404_/CLK _16084_/D vssd1 vssd1 vccd1 vccd1 hold649/A sky130_fd_sc_hd__dfxtp_1
X_13296_ _13289_/X _13295_/X _13296_/B1 vssd1 vssd1 vccd1 vccd1 _17555_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_224_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15035_ hold932/A _18303_/Q _15071_/S vssd1 vssd1 vccd1 vccd1 hold368/A sky130_fd_sc_hd__mux2_1
XFILLER_0_139_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12247_ _12341_/A _12365_/B _12246_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _12247_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12178_ hold5167/X _12365_/B _12177_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _12178_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11129_ hold2546/X hold4701/X _11765_/C vssd1 vssd1 vccd1 vccd1 _11130_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16986_ _17834_/CLK _16986_/D vssd1 vssd1 vccd1 vccd1 _16986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_1316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15937_ _17284_/CLK _15937_/D vssd1 vssd1 vccd1 vccd1 hold525/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15868_ _17606_/CLK _15868_/D vssd1 vssd1 vccd1 vccd1 _15868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14819_ hold1845/X _14828_/B _14818_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14819_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17607_ _17703_/CLK _17607_/D vssd1 vssd1 vccd1 vccd1 _17607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15799_ _17425_/CLK _15799_/D vssd1 vssd1 vccd1 vccd1 _15799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08340_ _14395_/A hold1450/X hold115/X vssd1 vssd1 vccd1 vccd1 _08341_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_58_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17538_ _18380_/CLK _17538_/D vssd1 vssd1 vccd1 vccd1 _17538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08271_ hold1370/X _08268_/B _08270_/X _08361_/A vssd1 vssd1 vccd1 vccd1 _08271_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17469_ _17471_/CLK _17469_/D vssd1 vssd1 vccd1 vccd1 _17469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6005 _17541_/Q vssd1 vssd1 vccd1 vccd1 hold6005/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6016 _17536_/Q vssd1 vssd1 vccd1 vccd1 hold6016/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6027 _17533_/Q vssd1 vssd1 vccd1 vccd1 hold6027/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6038 data_in[17] vssd1 vssd1 vccd1 vccd1 hold251/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6049 becStatus[1] vssd1 vssd1 vccd1 vccd1 hold6049/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5304 _10807_/X vssd1 vssd1 vccd1 vccd1 _16759_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5315 _17038_/Q vssd1 vssd1 vccd1 vccd1 hold5315/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5326 _13396_/X vssd1 vssd1 vccd1 vccd1 _17585_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5337 _17683_/Q vssd1 vssd1 vccd1 vccd1 hold5337/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4603 _10456_/X vssd1 vssd1 vccd1 vccd1 _16642_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5348 _11404_/X vssd1 vssd1 vccd1 vccd1 _16958_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4614 _16837_/Q vssd1 vssd1 vccd1 vccd1 hold4614/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5359 _16969_/Q vssd1 vssd1 vccd1 vccd1 hold5359/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4625 _13735_/X vssd1 vssd1 vccd1 vccd1 _17698_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4636 _16909_/Q vssd1 vssd1 vccd1 vccd1 hold4636/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3902 _10120_/X vssd1 vssd1 vccd1 vccd1 _16530_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4647 _11836_/X vssd1 vssd1 vccd1 vccd1 _17102_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3913 _16592_/Q vssd1 vssd1 vccd1 vccd1 hold3913/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4658 _17718_/Q vssd1 vssd1 vccd1 vccd1 hold4658/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4669 _10681_/X vssd1 vssd1 vccd1 vccd1 _16717_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3924 _13729_/X vssd1 vssd1 vccd1 vccd1 _17696_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3935 _17164_/Q vssd1 vssd1 vccd1 vccd1 hold3935/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3946 _16373_/Q vssd1 vssd1 vccd1 vccd1 hold3946/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3957 _11023_/X vssd1 vssd1 vccd1 vccd1 _16831_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_238_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout147 _12812_/S vssd1 vssd1 vccd1 vccd1 _12800_/S sky130_fd_sc_hd__buf_6
Xhold3968 _13519_/X vssd1 vssd1 vccd1 vccd1 _17626_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout158 _12905_/S vssd1 vssd1 vccd1 vccd1 _12971_/S sky130_fd_sc_hd__buf_4
Xhold3979 _10654_/X vssd1 vssd1 vccd1 vccd1 _16708_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07986_ _15555_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07986_/X sky130_fd_sc_hd__or2_1
Xfanout169 _12217_/A2 vssd1 vssd1 vccd1 vccd1 _12353_/B sky130_fd_sc_hd__buf_4
XFILLER_0_226_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09725_ hold833/X hold3734/X _10028_/C vssd1 vssd1 vccd1 vccd1 _09726_/B sky130_fd_sc_hd__mux2_1
X_09656_ hold2424/X hold3622/X _11204_/C vssd1 vssd1 vccd1 vccd1 _09657_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08607_ hold71/X hold829/X _08657_/S vssd1 vssd1 vccd1 vccd1 _08608_/B sky130_fd_sc_hd__mux2_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09587_ hold2838/X _16353_/Q _10475_/S vssd1 vssd1 vccd1 vccd1 _09588_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_139_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ hold684/X hold815/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold816/A sky130_fd_sc_hd__mux2_1
XFILLER_0_194_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08469_ hold2716/X _08486_/B _08468_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08469_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10500_ _10524_/A _10500_/B vssd1 vssd1 vccd1 vccd1 _10500_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11480_ hold1035/X hold4783/X _12173_/S vssd1 vssd1 vccd1 vccd1 _11481_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_163_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10431_ _10554_/A _10431_/B vssd1 vssd1 vccd1 vccd1 _10431_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13150_ _13150_/A _13294_/B vssd1 vssd1 vccd1 vccd1 _13150_/X sky130_fd_sc_hd__or2_1
X_10362_ _10554_/A _10362_/B vssd1 vssd1 vccd1 vccd1 _10362_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12101_ hold1650/X hold4793/X _13811_/C vssd1 vssd1 vccd1 vccd1 _12102_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_60_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5860 output79/X vssd1 vssd1 vccd1 vccd1 data_out[16] sky130_fd_sc_hd__buf_12
XFILLER_0_103_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5871 hold6016/X vssd1 vssd1 vccd1 vccd1 _13137_/A sky130_fd_sc_hd__dlygate4sd3_1
X_13081_ _13081_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _13081_/X sky130_fd_sc_hd__and2_1
X_10293_ _10530_/A _10293_/B vssd1 vssd1 vccd1 vccd1 _10293_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5882 output81/X vssd1 vssd1 vccd1 vccd1 data_out[18] sky130_fd_sc_hd__buf_12
Xhold5893 hold6035/X vssd1 vssd1 vccd1 vccd1 _13065_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12032_ hold2298/X hold3818/X _13409_/S vssd1 vssd1 vccd1 vccd1 _12033_/B sky130_fd_sc_hd__mux2_1
Xhold190 hold190/A vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ _18043_/CLK _16840_/D vssd1 vssd1 vccd1 vccd1 _16840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout670 _08351_/A vssd1 vssd1 vccd1 vccd1 _08367_/A sky130_fd_sc_hd__buf_4
XFILLER_0_219_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout681 _14356_/A vssd1 vssd1 vccd1 vccd1 _13897_/A sky130_fd_sc_hd__buf_4
XFILLER_0_189_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout692 _08851_/A vssd1 vssd1 vccd1 vccd1 _12987_/A sky130_fd_sc_hd__buf_4
X_16771_ _18036_/CLK _16771_/D vssd1 vssd1 vccd1 vccd1 _16771_/Q sky130_fd_sc_hd__dfxtp_1
X_13983_ hold2312/X _13986_/B _13982_/Y _14392_/A vssd1 vssd1 vccd1 vccd1 _13983_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_232_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15722_ _17161_/CLK _15722_/D vssd1 vssd1 vccd1 vccd1 _15722_/Q sky130_fd_sc_hd__dfxtp_1
X_12934_ hold2916/X _17489_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12934_/X sky130_fd_sc_hd__mux2_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15653_ _17262_/CLK _15653_/D vssd1 vssd1 vccd1 vccd1 _15653_/Q sky130_fd_sc_hd__dfxtp_1
X_18441_ _18453_/CLK _18441_/D vssd1 vssd1 vccd1 vccd1 _18441_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ hold2657/X _17466_/Q _12916_/S vssd1 vssd1 vccd1 vccd1 _12865_/X sky130_fd_sc_hd__mux2_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _14604_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14604_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _18372_/CLK _18372_/D vssd1 vssd1 vccd1 vccd1 _18372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11816_ hold2375/X hold4323/X _13811_/C vssd1 vssd1 vccd1 vccd1 _11817_/B sky130_fd_sc_hd__mux2_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _17899_/CLK _15584_/D vssd1 vssd1 vccd1 vccd1 _15584_/Q sky130_fd_sc_hd__dfxtp_1
X_12796_ _16211_/Q hold3350/X _12838_/S vssd1 vssd1 vccd1 vccd1 _12796_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17323_ _17338_/CLK hold193/X vssd1 vssd1 vccd1 vccd1 _17323_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14535_ _15215_/A _14541_/B vssd1 vssd1 vccd1 vccd1 _14535_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_230_1281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _17073_/Q _12323_/B _12323_/C vssd1 vssd1 vccd1 vccd1 _11747_/X sky130_fd_sc_hd__and3_1
XFILLER_0_12_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17254_ _17719_/CLK _17254_/D vssd1 vssd1 vccd1 vccd1 _17254_/Q sky130_fd_sc_hd__dfxtp_1
X_14466_ hold3110/X _14487_/B _14465_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _14466_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11678_ hold1611/X hold5161/X _12242_/S vssd1 vssd1 vccd1 vccd1 _11679_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_181_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16205_ _17437_/CLK _16205_/D vssd1 vssd1 vccd1 vccd1 _16205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13417_ hold5263/X _13814_/B _13416_/X _13417_/C1 vssd1 vssd1 vccd1 vccd1 _13417_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10629_ hold4225/X _10515_/A _10628_/X vssd1 vssd1 vccd1 vccd1 _10629_/Y sky130_fd_sc_hd__a21oi_1
X_17185_ _17279_/CLK _17185_/D vssd1 vssd1 vccd1 vccd1 _17185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14397_ hold915/X _14445_/B vssd1 vssd1 vccd1 vccd1 _14397_/X sky130_fd_sc_hd__or2_1
X_16136_ _18413_/CLK _16136_/D vssd1 vssd1 vccd1 vccd1 hold301/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13348_ hold4672/X _13862_/B _13347_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13348_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16067_ _16090_/CLK _16067_/D vssd1 vssd1 vccd1 vccd1 hold802/A sky130_fd_sc_hd__dfxtp_1
X_13279_ _13311_/A1 _13277_/X _13278_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13279_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3209 _10650_/Y vssd1 vssd1 vccd1 vccd1 _10651_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_257_wb_clk_i clkbuf_6_58_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18058_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15018_ _15233_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _15018_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2508 _14327_/X vssd1 vssd1 vccd1 vccd1 _17963_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2519 _14691_/X vssd1 vssd1 vccd1 vccd1 _18137_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07840_ hold2365/X _07865_/B _07839_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _07840_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1807 _16308_/Q vssd1 vssd1 vccd1 vccd1 _09447_/B sky130_fd_sc_hd__buf_1
Xhold1818 _07981_/X vssd1 vssd1 vccd1 vccd1 _15633_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1829 _18235_/Q vssd1 vssd1 vccd1 vccd1 hold1829/X sky130_fd_sc_hd__dlygate4sd3_1
X_16969_ _17850_/CLK _16969_/D vssd1 vssd1 vccd1 vccd1 _16969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09510_ _09984_/A _09510_/B vssd1 vssd1 vccd1 vccd1 _09510_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ _09447_/D _09478_/B vssd1 vssd1 vccd1 vccd1 _16306_/D sky130_fd_sc_hd__and2b_1
XFILLER_0_188_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09372_ _07805_/A _09362_/A _09386_/A hold856/X vssd1 vssd1 vccd1 vccd1 _09375_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08323_ _15547_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08323_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08254_ _15533_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08254_/X sky130_fd_sc_hd__or2_1
XFILLER_0_172_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08185_ _15085_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08185_/X sky130_fd_sc_hd__or2_1
XFILLER_0_166_1286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5101 _17613_/Q vssd1 vssd1 vccd1 vccd1 hold5101/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5112 _11464_/X vssd1 vssd1 vccd1 vccd1 _16978_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5123 _17229_/Q vssd1 vssd1 vccd1 vccd1 hold5123/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5134 _11578_/X vssd1 vssd1 vccd1 vccd1 _17016_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5145 _10480_/X vssd1 vssd1 vccd1 vccd1 _16650_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4400 _11208_/Y vssd1 vssd1 vccd1 vccd1 _11209_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4411 _16929_/Q vssd1 vssd1 vccd1 vccd1 hold4411/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5156 _17219_/Q vssd1 vssd1 vccd1 vccd1 hold5156/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4422 _13854_/Y vssd1 vssd1 vccd1 vccd1 _13855_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5167 _17248_/Q vssd1 vssd1 vccd1 vccd1 hold5167/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5178 _09796_/X vssd1 vssd1 vccd1 vccd1 _16422_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4433 _17109_/Q vssd1 vssd1 vccd1 vccd1 hold4433/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4444 _13867_/Y vssd1 vssd1 vccd1 vccd1 _17742_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5189 _17047_/Q vssd1 vssd1 vccd1 vccd1 hold5189/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3710 _16698_/Q vssd1 vssd1 vccd1 vccd1 hold3710/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4455 _11727_/Y vssd1 vssd1 vccd1 vccd1 _11728_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3721 _10372_/X vssd1 vssd1 vccd1 vccd1 _16614_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4466 _10324_/X vssd1 vssd1 vccd1 vccd1 _16598_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3732 _16483_/Q vssd1 vssd1 vccd1 vccd1 hold3732/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4477 _17349_/Q vssd1 vssd1 vccd1 vccd1 hold4477/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3743 _10273_/X vssd1 vssd1 vccd1 vccd1 _16581_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4488 _17588_/Q vssd1 vssd1 vccd1 vccd1 hold4488/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3754 _10306_/X vssd1 vssd1 vccd1 vccd1 _16592_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4499 _13842_/Y vssd1 vssd1 vccd1 vccd1 _13843_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3765 _16693_/Q vssd1 vssd1 vccd1 vccd1 hold3765/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3776 _10375_/X vssd1 vssd1 vccd1 vccd1 _16615_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3787 _17502_/Q vssd1 vssd1 vccd1 vccd1 hold3787/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3798 _09985_/X vssd1 vssd1 vccd1 vccd1 _16485_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07969_ hold1650/X _07978_/B _07968_/X _12103_/C1 vssd1 vssd1 vccd1 vccd1 _07969_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09708_ _09984_/A _09708_/B vssd1 vssd1 vccd1 vccd1 _09708_/X sky130_fd_sc_hd__or2_1
XFILLER_0_202_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10980_ _11655_/A _10980_/B vssd1 vssd1 vccd1 vccd1 _10980_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09639_ _11010_/A _09639_/B vssd1 vssd1 vccd1 vccd1 _09639_/X sky130_fd_sc_hd__or2_1
XFILLER_0_210_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12650_ hold3356/X _12649_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12651_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_183_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11601_ _12240_/A _11601_/B vssd1 vssd1 vccd1 vccd1 _11601_/X sky130_fd_sc_hd__or2_1
XFILLER_0_155_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12581_ hold3389/X _12580_/X _12923_/S vssd1 vssd1 vccd1 vccd1 _12582_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ _15215_/A _14326_/B vssd1 vssd1 vccd1 vccd1 _14320_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11532_ _11631_/A _11532_/B vssd1 vssd1 vccd1 vccd1 _11532_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14251_ hold3104/X _14268_/B _14250_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _14251_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11463_ _11658_/A _11463_/B vssd1 vssd1 vccd1 vccd1 _11463_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13202_ _17576_/Q _17110_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13202_/X sky130_fd_sc_hd__mux2_1
X_10414_ hold3642/X _10604_/B _10413_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _10414_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14182_ _14413_/A _14204_/B vssd1 vssd1 vccd1 vccd1 _14182_/X sky130_fd_sc_hd__or2_1
X_11394_ _12219_/A _11394_/B vssd1 vssd1 vccd1 vccd1 _11394_/X sky130_fd_sc_hd__or2_1
XFILLER_0_238_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13133_ _13132_/X hold3501/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13133_/X sky130_fd_sc_hd__mux2_1
X_10345_ hold3921/X _10631_/B _10344_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10345_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_350_wb_clk_i clkbuf_6_40_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17620_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_237_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5690 _12205_/X vssd1 vssd1 vccd1 vccd1 _17225_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13064_ _13051_/X _13063_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17526_/D sky130_fd_sc_hd__o21a_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941_ _18005_/CLK _17941_/D vssd1 vssd1 vccd1 vccd1 _17941_/Q sky130_fd_sc_hd__dfxtp_1
X_10276_ hold3846/X _10625_/B _10275_/X _14769_/C1 vssd1 vssd1 vccd1 vccd1 _10276_/X
+ sky130_fd_sc_hd__o211a_1
X_12015_ _12198_/A _12015_/B vssd1 vssd1 vccd1 vccd1 _12015_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17872_ _17904_/CLK _17872_/D vssd1 vssd1 vccd1 vccd1 _17872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16823_ _18056_/CLK _16823_/D vssd1 vssd1 vccd1 vccd1 _16823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_232_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_219_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13966_ hold951/X _13998_/B vssd1 vssd1 vccd1 vccd1 _13966_/X sky130_fd_sc_hd__or2_1
X_16754_ _18021_/CLK _16754_/D vssd1 vssd1 vccd1 vccd1 _16754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15705_ _17608_/CLK _15705_/D vssd1 vssd1 vccd1 vccd1 _15705_/Q sky130_fd_sc_hd__dfxtp_1
X_12917_ hold3312/X _12916_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12917_/X sky130_fd_sc_hd__mux2_1
X_16685_ _18211_/CLK _16685_/D vssd1 vssd1 vccd1 vccd1 _16685_/Q sky130_fd_sc_hd__dfxtp_1
X_13897_ _13897_/A _13897_/B vssd1 vssd1 vccd1 vccd1 _17756_/D sky130_fd_sc_hd__and2_1
XFILLER_0_152_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_45_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_45_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_18424_ _18424_/CLK _18424_/D vssd1 vssd1 vccd1 vccd1 _18424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12848_ hold3398/X _12847_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12849_/B sky130_fd_sc_hd__mux2_1
X_15636_ _17264_/CLK _15636_/D vssd1 vssd1 vccd1 vccd1 _15636_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18355_ _18387_/CLK hold985/X vssd1 vssd1 vccd1 vccd1 hold984/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15567_ _17204_/CLK _15567_/D vssd1 vssd1 vccd1 vccd1 _15567_/Q sky130_fd_sc_hd__dfxtp_1
X_12779_ hold4065/X _12778_/X _12839_/S vssd1 vssd1 vccd1 vccd1 _12780_/B sky130_fd_sc_hd__mux2_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17306_ _17321_/CLK _17306_/D vssd1 vssd1 vccd1 vccd1 hold457/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14518_ hold1295/X _14541_/B _14517_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _14518_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18286_ _18324_/CLK _18286_/D vssd1 vssd1 vccd1 vccd1 _18286_/Q sky130_fd_sc_hd__dfxtp_1
X_15498_ _15498_/A _15498_/B vssd1 vssd1 vccd1 vccd1 _18428_/D sky130_fd_sc_hd__and2_1
XFILLER_0_25_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14449_ hold927/X _14499_/B vssd1 vssd1 vccd1 vccd1 _14449_/X sky130_fd_sc_hd__or2_1
X_17237_ _17269_/CLK _17237_/D vssd1 vssd1 vccd1 vccd1 _17237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_438_wb_clk_i clkbuf_6_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17626_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_226_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold904 hold904/A vssd1 vssd1 vccd1 vccd1 hold904/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17168_ _17229_/CLK _17168_/D vssd1 vssd1 vccd1 vccd1 _17168_/Q sky130_fd_sc_hd__dfxtp_1
Xhold915 hold915/A vssd1 vssd1 vccd1 vccd1 hold915/X sky130_fd_sc_hd__buf_12
Xhold926 hold926/A vssd1 vssd1 vccd1 vccd1 hold926/X sky130_fd_sc_hd__clkbuf_2
Xhold937 hold948/X vssd1 vssd1 vccd1 vccd1 hold937/X sky130_fd_sc_hd__clkbuf_4
X_16119_ _17347_/CLK _16119_/D vssd1 vssd1 vccd1 vccd1 hold175/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold948 hold948/A vssd1 vssd1 vccd1 vccd1 hold948/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09990_ _13086_/A _09984_/A _09989_/X vssd1 vssd1 vccd1 vccd1 _09990_/Y sky130_fd_sc_hd__a21oi_1
Xhold959 hold959/A vssd1 vssd1 vccd1 vccd1 hold959/X sky130_fd_sc_hd__dlygate4sd3_1
X_17099_ _17878_/CLK _17099_/D vssd1 vssd1 vccd1 vccd1 _17099_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3006 _17894_/Q vssd1 vssd1 vccd1 vccd1 hold3006/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08941_ hold684/X _16088_/Q _08991_/S vssd1 vssd1 vccd1 vccd1 hold685/A sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3017 _18064_/Q vssd1 vssd1 vccd1 vccd1 hold3017/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3028 _07931_/X vssd1 vssd1 vccd1 vccd1 _15609_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3039 _17875_/Q vssd1 vssd1 vccd1 vccd1 hold3039/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2305 _08210_/X vssd1 vssd1 vccd1 vccd1 _15741_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2316 _18052_/Q vssd1 vssd1 vccd1 vccd1 hold2316/X sky130_fd_sc_hd__dlygate4sd3_1
X_08872_ hold618/X hold797/X _08930_/S vssd1 vssd1 vccd1 vccd1 hold798/A sky130_fd_sc_hd__mux2_1
Xhold2327 _08324_/X vssd1 vssd1 vccd1 vccd1 _15795_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2338 _15655_/Q vssd1 vssd1 vccd1 vccd1 hold2338/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2349 _18378_/Q vssd1 vssd1 vccd1 vccd1 hold2349/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1604 _15636_/Q vssd1 vssd1 vccd1 vccd1 hold1604/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1615 _09231_/X vssd1 vssd1 vccd1 vccd1 _16227_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07823_ hold597/X hold384/X _09496_/A _15169_/A vssd1 vssd1 vccd1 vccd1 _09121_/B
+ sky130_fd_sc_hd__or4b_1
Xhold1626 _16199_/Q vssd1 vssd1 vccd1 vccd1 hold1626/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1637 _15881_/Q vssd1 vssd1 vccd1 vccd1 hold1637/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1648 _18347_/Q vssd1 vssd1 vccd1 vccd1 hold1648/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1659 _13963_/X vssd1 vssd1 vccd1 vccd1 _17788_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_237_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09424_ _09438_/B _16298_/Q vssd1 vssd1 vccd1 vccd1 _09424_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09355_ _15547_/A _15165_/A _09359_/C vssd1 vssd1 vccd1 vccd1 _09356_/C sky130_fd_sc_hd__or3_1
XFILLER_0_212_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08306_ hold1566/X _08336_/A2 _08305_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _08306_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09286_ hold406/X hold363/X vssd1 vssd1 vccd1 vccd1 _09315_/B sky130_fd_sc_hd__or2_2
XFILLER_0_191_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08237_ hold2687/X _08262_/B _08236_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _08237_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_179_wb_clk_i clkbuf_6_49_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18325_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08168_ _15519_/A hold1506/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08169_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_108_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17331_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_120_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08099_ hold1256/X _08088_/B _08098_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _08099_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4230 _17569_/Q vssd1 vssd1 vccd1 vccd1 hold4230/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10130_ hold1271/X hold4238/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10131_/B sky130_fd_sc_hd__mux2_1
Xhold4241 _13831_/Y vssd1 vssd1 vccd1 vccd1 _17730_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4252 _11172_/Y vssd1 vssd1 vccd1 vccd1 _11173_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4263 _13825_/Y vssd1 vssd1 vccd1 vccd1 _17728_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4274 _12354_/Y vssd1 vssd1 vccd1 vccd1 _12355_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4285 _11163_/Y vssd1 vssd1 vccd1 vccd1 _11164_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3540 _17441_/Q vssd1 vssd1 vccd1 vccd1 hold3540/X sky130_fd_sc_hd__dlygate4sd3_1
X_10061_ _16511_/Q _10601_/B _10385_/S vssd1 vssd1 vccd1 vccd1 _10061_/X sky130_fd_sc_hd__and3_1
XTAP_6458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3551 _10177_/X vssd1 vssd1 vccd1 vccd1 _16549_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4296 _11799_/Y vssd1 vssd1 vccd1 vccd1 _11800_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_234_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3562 _16412_/Q vssd1 vssd1 vccd1 vccd1 hold3562/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3573 _09601_/X vssd1 vssd1 vccd1 vccd1 _16357_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3584 _16419_/Q vssd1 vssd1 vccd1 vccd1 hold3584/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3595 _16548_/Q vssd1 vssd1 vccd1 vccd1 hold3595/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2850 _17960_/Q vssd1 vssd1 vccd1 vccd1 hold2850/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2861 _15762_/Q vssd1 vssd1 vccd1 vccd1 hold2861/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2872 _14091_/X vssd1 vssd1 vccd1 vccd1 _17850_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2883 _15720_/Q vssd1 vssd1 vccd1 vccd1 hold2883/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2894 _08263_/X vssd1 vssd1 vccd1 vccd1 _15766_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13820_ _17727_/Q _13829_/B _13829_/C vssd1 vssd1 vccd1 vccd1 _13820_/X sky130_fd_sc_hd__and3_1
XFILLER_0_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13751_ hold2758/X hold5233/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13752_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_202_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10963_ hold5109/X _11153_/B _10962_/X _14354_/A vssd1 vssd1 vccd1 vccd1 _10963_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12702_ _12786_/A _12702_/B vssd1 vssd1 vccd1 vccd1 _17410_/D sky130_fd_sc_hd__and2_1
X_16470_ _18325_/CLK _16470_/D vssd1 vssd1 vccd1 vccd1 _16470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13682_ hold2861/X hold5460/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13683_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10894_ hold4979/X _11186_/B _10893_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10894_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15421_ hold489/X _15441_/A2 _09386_/D hold849/X _15416_/X vssd1 vssd1 vccd1 vccd1
+ _15422_/D sky130_fd_sc_hd__a221o_1
X_12633_ _12864_/A _12633_/B vssd1 vssd1 vccd1 vccd1 _17387_/D sky130_fd_sc_hd__and2_1
XFILLER_0_39_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18140_ _18210_/CLK _18140_/D vssd1 vssd1 vccd1 vccd1 _18140_/Q sky130_fd_sc_hd__dfxtp_1
X_15352_ _15480_/A _15352_/B _15352_/C _15352_/D vssd1 vssd1 vccd1 vccd1 _15352_/X
+ sky130_fd_sc_hd__or4_1
X_12564_ _12906_/A _12564_/B vssd1 vssd1 vccd1 vccd1 _17364_/D sky130_fd_sc_hd__and2_1
XFILLER_0_81_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14303_ hold1588/X _14333_/A2 _14302_/X _14552_/C1 vssd1 vssd1 vccd1 vccd1 _14303_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11515_ hold4115/X _11792_/B _11514_/X _14143_/C1 vssd1 vssd1 vccd1 vccd1 _11515_/X
+ sky130_fd_sc_hd__o211a_1
X_18071_ _18073_/CLK hold822/X vssd1 vssd1 vccd1 vccd1 _18071_/Q sky130_fd_sc_hd__dfxtp_1
X_15283_ _15490_/A1 _15275_/X _15282_/X _15490_/B1 hold5912/A vssd1 vssd1 vccd1 vccd1
+ _15283_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_0_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12495_ hold17/X _12445_/A _12445_/B _12494_/X _09057_/A vssd1 vssd1 vccd1 vccd1
+ hold18/A sky130_fd_sc_hd__o311a_1
XFILLER_0_108_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17022_ _17902_/CLK _17022_/D vssd1 vssd1 vccd1 vccd1 _17022_/Q sky130_fd_sc_hd__dfxtp_1
X_14234_ hold927/X _14284_/B vssd1 vssd1 vccd1 vccd1 _14234_/X sky130_fd_sc_hd__or2_1
XFILLER_0_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11446_ hold5376/X _11732_/B _11445_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _11446_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14165_ hold2215/X _14198_/B _14164_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _14165_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11377_ hold5082/X _11765_/B _11376_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _11377_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13116_ hold4259/X _13115_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13116_/X sky130_fd_sc_hd__mux2_2
X_10328_ hold1220/X _16600_/Q _11183_/C vssd1 vssd1 vccd1 vccd1 _10329_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _15549_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14096_/X sky130_fd_sc_hd__or2_1
XFILLER_0_147_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _13056_/C _13044_/X _13046_/X _09339_/A vssd1 vssd1 vccd1 vccd1 _13047_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_17924_ _18052_/CLK _17924_/D vssd1 vssd1 vccd1 vccd1 _17924_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ hold1700/X _16577_/Q _10646_/C vssd1 vssd1 vccd1 vccd1 _10260_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_147_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_218_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17855_ _17867_/CLK _17855_/D vssd1 vssd1 vccd1 vccd1 _17855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16806_ _18041_/CLK _16806_/D vssd1 vssd1 vccd1 vccd1 _16806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17786_ _18432_/CLK _17786_/D vssd1 vssd1 vccd1 vccd1 _17786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14998_ _15213_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14998_/X sky130_fd_sc_hd__or2_1
XFILLER_0_88_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16737_ _18036_/CLK _16737_/D vssd1 vssd1 vccd1 vccd1 _16737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13949_ hold2039/X _13995_/A2 _13948_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _13949_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16668_ _18226_/CLK _16668_/D vssd1 vssd1 vccd1 vccd1 _16668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18407_ _18462_/CLK _18407_/D vssd1 vssd1 vccd1 vccd1 _18407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15619_ _17905_/CLK _15619_/D vssd1 vssd1 vccd1 vccd1 _15619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16599_ _18221_/CLK _16599_/D vssd1 vssd1 vccd1 vccd1 _16599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09140_ hold933/X _09176_/B vssd1 vssd1 vccd1 vccd1 _09140_/X sky130_fd_sc_hd__or2_1
X_18338_ _18376_/CLK _18338_/D vssd1 vssd1 vccd1 vccd1 _18338_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_6_wb_clk_i clkbuf_6_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17452_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_115_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09071_ hold1301/X _09106_/B _09070_/X _12987_/A vssd1 vssd1 vccd1 vccd1 _09071_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18269_ _18375_/CLK _18269_/D vssd1 vssd1 vccd1 vccd1 _18269_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_272_wb_clk_i clkbuf_6_57_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18164_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08022_ hold1953/X _08029_/B _08021_/X _08167_/A vssd1 vssd1 vccd1 vccd1 _08022_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold701 hold701/A vssd1 vssd1 vccd1 vccd1 hold701/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold712 hold712/A vssd1 vssd1 vccd1 vccd1 input70/A sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_201_wb_clk_i clkbuf_6_53_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18356_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold723 hold723/A vssd1 vssd1 vccd1 vccd1 hold723/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold734 hold734/A vssd1 vssd1 vccd1 vccd1 hold734/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold745 hold745/A vssd1 vssd1 vccd1 vccd1 hold745/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold756 hold756/A vssd1 vssd1 vccd1 vccd1 hold756/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold767 hold767/A vssd1 vssd1 vccd1 vccd1 hold767/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 hold778/A vssd1 vssd1 vccd1 vccd1 hold778/X sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _10067_/A _10067_/B _09972_/X _15228_/C1 vssd1 vssd1 vccd1 vccd1 _09973_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_228_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold789 hold789/A vssd1 vssd1 vccd1 vccd1 hold789/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08924_ hold82/X hold468/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold469/A sky130_fd_sc_hd__mux2_1
Xhold2102 hold2225/X vssd1 vssd1 vccd1 vccd1 hold2226/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2113 _18133_/Q vssd1 vssd1 vccd1 vccd1 hold2113/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2124 _14153_/X vssd1 vssd1 vccd1 vccd1 _17880_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2135 _18161_/Q vssd1 vssd1 vccd1 vccd1 hold2135/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1401 _09310_/X vssd1 vssd1 vccd1 vccd1 _16265_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2146 _09316_/X vssd1 vssd1 vccd1 vccd1 _16268_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08855_ _12426_/A _08855_/B vssd1 vssd1 vccd1 vccd1 _16046_/D sky130_fd_sc_hd__and2_1
Xhold2157 _18361_/Q vssd1 vssd1 vccd1 vccd1 hold2157/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1412 _08130_/X vssd1 vssd1 vccd1 vccd1 _08131_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1423 _18307_/Q vssd1 vssd1 vccd1 vccd1 hold1423/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2168 _14137_/X vssd1 vssd1 vccd1 vccd1 _17872_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 _18386_/Q vssd1 vssd1 vccd1 vccd1 hold1434/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2179 _18447_/Q vssd1 vssd1 vccd1 vccd1 hold2179/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1445 _09423_/X vssd1 vssd1 vccd1 vccd1 _16297_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1456 _14651_/X vssd1 vssd1 vccd1 vccd1 _18118_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07806_ _07786_/A _07801_/B _09339_/B vssd1 vssd1 vccd1 vccd1 _07806_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1467 _15088_/X vssd1 vssd1 vccd1 vccd1 _18328_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08786_ _15473_/A hold155/X vssd1 vssd1 vccd1 vccd1 _16013_/D sky130_fd_sc_hd__and2_1
XFILLER_0_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1478 _15510_/X vssd1 vssd1 vccd1 vccd1 _18433_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1489 _15745_/Q vssd1 vssd1 vccd1 vccd1 hold1489/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09407_ _07804_/A _09447_/C _15284_/A _09406_/X vssd1 vssd1 vccd1 vccd1 _09407_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09338_ hold1297/X _09325_/B _09337_/X _12924_/A vssd1 vssd1 vccd1 vccd1 _09338_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09269_ hold220/X _16246_/Q hold271/X vssd1 vssd1 vccd1 vccd1 hold365/A sky130_fd_sc_hd__mux2_1
XFILLER_0_145_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11300_ _17772_/Q _16924_/Q _11741_/C vssd1 vssd1 vccd1 vccd1 _11301_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_16_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12280_ hold5107/X _12374_/B _12279_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _12280_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11231_ hold1422/X _16901_/Q _11717_/C vssd1 vssd1 vccd1 vccd1 _11232_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11162_ _16878_/Q _11162_/B _11162_/C vssd1 vssd1 vccd1 vccd1 _11162_/X sky130_fd_sc_hd__and3_1
XTAP_6211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4060 _10792_/X vssd1 vssd1 vccd1 vccd1 _16754_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10113_ _10563_/A _10113_/B vssd1 vssd1 vccd1 vccd1 _10113_/X sky130_fd_sc_hd__or2_1
Xhold4071 _10732_/X vssd1 vssd1 vccd1 vccd1 _16734_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4082 _10828_/X vssd1 vssd1 vccd1 vccd1 _16766_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15970_ _16129_/CLK _15970_/D vssd1 vssd1 vccd1 vccd1 hold205/A sky130_fd_sc_hd__dfxtp_1
XTAP_5510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11093_ hold2781/X hold5070/X _11216_/C vssd1 vssd1 vccd1 vccd1 _11094_/B sky130_fd_sc_hd__mux2_1
Xhold4093 _17059_/Q vssd1 vssd1 vccd1 vccd1 hold4093/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_234_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3370 _17389_/Q vssd1 vssd1 vccd1 vccd1 hold3370/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10044_ _13230_/A _10386_/A _10043_/X vssd1 vssd1 vccd1 vccd1 _10044_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14921_ hold3182/X _14952_/B _14920_/X _15202_/C1 vssd1 vssd1 vccd1 vccd1 _14921_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3381 _17359_/Q vssd1 vssd1 vccd1 vccd1 hold3381/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3392 _17442_/Q vssd1 vssd1 vccd1 vccd1 hold3392/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__clkbuf_2
XTAP_5565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_76_wb_clk_i clkbuf_6_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17514_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2680 _14707_/X vssd1 vssd1 vccd1 vccd1 _18145_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17640_ _17672_/CLK _17640_/D vssd1 vssd1 vccd1 vccd1 _17640_/Q sky130_fd_sc_hd__dfxtp_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ _15191_/A _14892_/B vssd1 vssd1 vccd1 vccd1 _14852_/X sky130_fd_sc_hd__or2_1
XTAP_5598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2691 _15616_/Q vssd1 vssd1 vccd1 vccd1 hold2691/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1990 _16263_/Q vssd1 vssd1 vccd1 vccd1 hold1990/X sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ hold4300/X _13719_/A _13802_/X vssd1 vssd1 vccd1 vccd1 _13803_/Y sky130_fd_sc_hd__a21oi_1
X_14783_ hold2583/X _14774_/B _14782_/X _15218_/C1 vssd1 vssd1 vccd1 vccd1 _14783_/X
+ sky130_fd_sc_hd__o211a_1
X_17571_ _17648_/CLK _17571_/D vssd1 vssd1 vccd1 vccd1 _17571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11995_ hold4857/X _13886_/B _11994_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _11995_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16522_ _18176_/CLK _16522_/D vssd1 vssd1 vccd1 vccd1 _16522_/Q sky130_fd_sc_hd__dfxtp_1
X_13734_ _13734_/A _13734_/B vssd1 vssd1 vccd1 vccd1 _13734_/X sky130_fd_sc_hd__or2_1
X_10946_ hold2109/X _16806_/Q _11732_/C vssd1 vssd1 vccd1 vccd1 _10947_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16453_ _18334_/CLK _16453_/D vssd1 vssd1 vccd1 vccd1 _16453_/Q sky130_fd_sc_hd__dfxtp_1
X_13665_ _13773_/A _13665_/B vssd1 vssd1 vccd1 vccd1 _13665_/X sky130_fd_sc_hd__or2_1
X_10877_ hold783/X _16783_/Q _11654_/S vssd1 vssd1 vccd1 vccd1 _10878_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_156_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _15404_/A _15404_/B vssd1 vssd1 vccd1 vccd1 _18416_/D sky130_fd_sc_hd__and2_1
X_12616_ hold1155/X _17383_/Q _12850_/S vssd1 vssd1 vccd1 vccd1 _12616_/X sky130_fd_sc_hd__mux2_1
X_16384_ _16480_/CLK _16384_/D vssd1 vssd1 vccd1 vccd1 _16384_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _13788_/A _13596_/B vssd1 vssd1 vccd1 vccd1 _13596_/X sky130_fd_sc_hd__or2_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18123_ _18149_/CLK _18123_/D vssd1 vssd1 vccd1 vccd1 _18123_/Q sky130_fd_sc_hd__dfxtp_1
X_15335_ hold343/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15335_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12547_ hold2361/X _17360_/Q _12925_/S vssd1 vssd1 vccd1 vccd1 _12547_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_227_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15266_ _17330_/Q _09362_/C _09362_/D hold753/X vssd1 vssd1 vccd1 vccd1 _15266_/X
+ sky130_fd_sc_hd__a22o_1
X_18054_ _18054_/CLK _18054_/D vssd1 vssd1 vccd1 vccd1 _18054_/Q sky130_fd_sc_hd__dfxtp_1
X_12478_ _17332_/Q _12506_/B vssd1 vssd1 vccd1 vccd1 _12478_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_3 _13068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17005_ _17853_/CLK _17005_/D vssd1 vssd1 vccd1 vccd1 _17005_/Q sky130_fd_sc_hd__dfxtp_1
X_14217_ _14897_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14230_/B sky130_fd_sc_hd__or2_2
X_11429_ hold3114/X hold5659/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11430_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_111_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15197_ _15197_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15197_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14148_ _15547_/A _14148_/B vssd1 vssd1 vccd1 vccd1 _14148_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14079_ hold1258/X _14094_/B _14078_/X _14211_/C1 vssd1 vssd1 vccd1 vccd1 _14079_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_225_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17907_ _17907_/CLK _17907_/D vssd1 vssd1 vccd1 vccd1 _17907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08640_ _15374_/A _08640_/B vssd1 vssd1 vccd1 vccd1 _15942_/D sky130_fd_sc_hd__and2_1
XFILLER_0_83_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17838_ _17838_/CLK _17838_/D vssd1 vssd1 vccd1 vccd1 _17838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08571_ _12390_/A _08571_/B vssd1 vssd1 vccd1 vccd1 _15909_/D sky130_fd_sc_hd__and2_1
XFILLER_0_117_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17769_ _17865_/CLK _17769_/D vssd1 vssd1 vccd1 vccd1 _17769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_453_wb_clk_i clkbuf_6_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17690_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_228_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09123_ _07788_/A _09120_/Y _09122_/Y hold6085/X vssd1 vssd1 vccd1 vccd1 _09123_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09054_ hold82/X hold396/X _09060_/S vssd1 vssd1 vccd1 vccd1 hold397/A sky130_fd_sc_hd__mux2_1
XFILLER_0_32_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08005_ _15519_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08005_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold520 hold520/A vssd1 vssd1 vccd1 vccd1 hold520/X sky130_fd_sc_hd__buf_4
Xhold531 hold531/A vssd1 vssd1 vccd1 vccd1 hold531/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold542 hold542/A vssd1 vssd1 vccd1 vccd1 hold542/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold553 hold596/X vssd1 vssd1 vccd1 vccd1 hold597/A sky130_fd_sc_hd__buf_6
Xhold564 hold564/A vssd1 vssd1 vccd1 vccd1 hold564/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold575 hold575/A vssd1 vssd1 vccd1 vccd1 hold575/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 hold586/A vssd1 vssd1 vccd1 vccd1 hold586/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold597 hold597/A vssd1 vssd1 vccd1 vccd1 hold597/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_198_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09956_ hold1949/X _16476_/Q _10040_/C vssd1 vssd1 vccd1 vccd1 _09957_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08907_ _12418_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _16071_/D sky130_fd_sc_hd__and2_1
XFILLER_0_148_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ hold2550/X _16453_/Q _10031_/C vssd1 vssd1 vccd1 vccd1 _09888_/B sky130_fd_sc_hd__mux2_1
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1220 _18158_/Q vssd1 vssd1 vccd1 vccd1 hold1220/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1231 _17905_/Q vssd1 vssd1 vccd1 vccd1 hold1231/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08838_ hold254/X hold386/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08839_/B sky130_fd_sc_hd__mux2_1
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1242 _16255_/Q vssd1 vssd1 vccd1 vccd1 hold1242/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1253 hold641/X vssd1 vssd1 vccd1 vccd1 hold1253/X sky130_fd_sc_hd__buf_4
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1264 _16248_/Q vssd1 vssd1 vccd1 vccd1 hold1264/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1275 _15678_/Q vssd1 vssd1 vccd1 vccd1 hold1275/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1286 _14207_/X vssd1 vssd1 vccd1 vccd1 _17906_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ hold215/X hold660/X _08779_/S vssd1 vssd1 vccd1 vccd1 _08770_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1297 _16279_/Q vssd1 vssd1 vccd1 vccd1 hold1297/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _11088_/A _10800_/B vssd1 vssd1 vccd1 vccd1 _10800_/X sky130_fd_sc_hd__or2_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11780_ _17084_/Q _12323_/B _12323_/C vssd1 vssd1 vccd1 vccd1 _11780_/X sky130_fd_sc_hd__and3_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10731_ _11100_/A _10731_/B vssd1 vssd1 vccd1 vccd1 _10731_/X sky130_fd_sc_hd__or2_1
XFILLER_0_177_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_194_wb_clk_i clkbuf_6_52_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18378_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13450_ hold4867/X _13862_/B _13449_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13450_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10662_ _11049_/A _10662_/B vssd1 vssd1 vccd1 vccd1 _10662_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_123_wb_clk_i clkbuf_6_22_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17320_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12401_ hold23/X hold357/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12402_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_137_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13381_ hold5470/X _13847_/B _13380_/X _13765_/C1 vssd1 vssd1 vccd1 vccd1 _13381_/X
+ sky130_fd_sc_hd__o211a_1
X_10593_ hold3468/X _10563_/A _10592_/X vssd1 vssd1 vccd1 vccd1 _10593_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15120_ hold2709/X hold341/X _15119_/X _15048_/A vssd1 vssd1 vccd1 vccd1 _15120_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12332_ _17268_/Q _12332_/B _12332_/C vssd1 vssd1 vccd1 vccd1 _12332_/X sky130_fd_sc_hd__and3_1
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15051_ _15213_/A hold2224/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15052_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12263_ hold3043/X _17245_/Q _12362_/C vssd1 vssd1 vccd1 vccd1 _12264_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14002_ _14395_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14002_/X sky130_fd_sc_hd__or2_1
X_11214_ hold4347/X _11103_/A _11213_/X vssd1 vssd1 vccd1 vccd1 _11214_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12194_ hold2512/X _17222_/Q _13796_/S vssd1 vssd1 vccd1 vccd1 _12195_/B sky130_fd_sc_hd__mux2_1
Xoutput73 _13137_/A vssd1 vssd1 vccd1 vccd1 output73/X sky130_fd_sc_hd__buf_6
XTAP_6030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11145_ hold3508/X _11049_/A _11144_/X vssd1 vssd1 vccd1 vccd1 _11145_/Y sky130_fd_sc_hd__a21oi_1
Xoutput84 _13217_/A vssd1 vssd1 vccd1 vccd1 output84/X sky130_fd_sc_hd__buf_6
XFILLER_0_222_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput95 _13297_/A vssd1 vssd1 vccd1 vccd1 output95/X sky130_fd_sc_hd__buf_6
XTAP_6052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15953_ _17300_/CLK _15953_/D vssd1 vssd1 vccd1 vccd1 hold861/A sky130_fd_sc_hd__dfxtp_1
X_11076_ _11655_/A _11076_/B vssd1 vssd1 vccd1 vccd1 _11076_/X sky130_fd_sc_hd__or2_1
XTAP_6096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10027_ _11203_/A _10027_/B vssd1 vssd1 vccd1 vccd1 _10027_/Y sky130_fd_sc_hd__nor2_1
XTAP_5373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14904_ _14974_/A _14910_/B vssd1 vssd1 vccd1 vccd1 _14904_/X sky130_fd_sc_hd__or2_1
XFILLER_0_204_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ _17561_/CLK _15884_/D vssd1 vssd1 vccd1 vccd1 _15884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17623_ _17720_/CLK _17623_/D vssd1 vssd1 vccd1 vccd1 _17623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14835_ hold2865/X _14826_/B _14834_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _14835_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _18229_/CLK _17554_/D vssd1 vssd1 vccd1 vccd1 _17554_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14766_ _15213_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14766_/X sky130_fd_sc_hd__or2_1
X_11978_ hold955/X hold5773/X _12362_/C vssd1 vssd1 vccd1 vccd1 _11979_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16505_ _18386_/CLK _16505_/D vssd1 vssd1 vccd1 vccd1 _16505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10929_ _11121_/A _10929_/B vssd1 vssd1 vccd1 vccd1 _10929_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13717_ hold4841/X _13811_/B _13716_/X _12822_/A vssd1 vssd1 vccd1 vccd1 _13717_/X
+ sky130_fd_sc_hd__o211a_1
X_14697_ hold1209/X _14720_/B _14696_/X _14697_/C1 vssd1 vssd1 vccd1 vccd1 _14697_/X
+ sky130_fd_sc_hd__o211a_1
X_17485_ _17486_/CLK _17485_/D vssd1 vssd1 vccd1 vccd1 _17485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16436_ _18381_/CLK _16436_/D vssd1 vssd1 vccd1 vccd1 _16436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13648_ hold5289/X _13856_/B _13647_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13648_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16367_ _18376_/CLK _16367_/D vssd1 vssd1 vccd1 vccd1 _16367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13579_ hold4003/X _13795_/A2 _13578_/X _13729_/C1 vssd1 vssd1 vccd1 vccd1 _13579_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18106_ _18106_/CLK hold960/X vssd1 vssd1 vccd1 vccd1 hold959/A sky130_fd_sc_hd__dfxtp_1
X_15318_ hold487/X _15484_/A2 _09392_/D hold839/X vssd1 vssd1 vccd1 vccd1 _15318_/X
+ sky130_fd_sc_hd__a22o_1
X_16298_ _18460_/CLK _16298_/D vssd1 vssd1 vccd1 vccd1 _16298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5508 _13405_/X vssd1 vssd1 vccd1 vccd1 _17588_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5519 _17611_/Q vssd1 vssd1 vccd1 vccd1 hold5519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18037_ _18061_/CLK _18037_/D vssd1 vssd1 vccd1 vccd1 _18037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15249_ hold689/X _15485_/A2 _15488_/A2 hold844/X _15248_/X vssd1 vssd1 vccd1 vccd1
+ _15252_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_169_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4807 _16898_/Q vssd1 vssd1 vccd1 vccd1 hold4807/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4818 _10936_/X vssd1 vssd1 vccd1 vccd1 _16802_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4829 _16437_/Q vssd1 vssd1 vccd1 vccd1 hold4829/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_238_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09810_ _09912_/A _09810_/B vssd1 vssd1 vccd1 vccd1 _09810_/X sky130_fd_sc_hd__or2_1
Xfanout307 _09984_/A vssd1 vssd1 vccd1 vccd1 _09933_/A sky130_fd_sc_hd__buf_4
Xfanout318 _11088_/A vssd1 vssd1 vccd1 vccd1 _11121_/A sky130_fd_sc_hd__buf_4
XFILLER_0_22_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout329 fanout335/A vssd1 vssd1 vccd1 vccd1 _10386_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_201_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09741_ _09933_/A _09741_/B vssd1 vssd1 vccd1 vccd1 _09741_/X sky130_fd_sc_hd__or2_1
XFILLER_0_185_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09672_ _09954_/A _09672_/B vssd1 vssd1 vccd1 vccd1 _09672_/X sky130_fd_sc_hd__or2_1
XFILLER_0_207_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_4_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_4_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08623_ hold77/X hold751/X _08623_/S vssd1 vssd1 vccd1 vccd1 hold752/A sky130_fd_sc_hd__mux2_1
XFILLER_0_179_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ hold163/X hold281/X _08592_/S vssd1 vssd1 vccd1 vccd1 hold282/A sky130_fd_sc_hd__mux2_1
XFILLER_0_210_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08485_ hold2343/X _08488_/B _08484_/Y _08143_/A vssd1 vssd1 vccd1 vccd1 _08485_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09106_ _15547_/A _09106_/B vssd1 vssd1 vccd1 vccd1 _09106_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_45_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09037_ _15314_/A _09037_/B vssd1 vssd1 vccd1 vccd1 _16135_/D sky130_fd_sc_hd__and2_1
XFILLER_0_143_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold350 hold350/A vssd1 vssd1 vccd1 vccd1 hold350/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold361 hold361/A vssd1 vssd1 vccd1 vccd1 hold361/X sky130_fd_sc_hd__clkbuf_2
Xhold372 input18/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__buf_1
Xhold383 input44/X vssd1 vssd1 vccd1 vccd1 hold383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 input32/X vssd1 vssd1 vccd1 vccd1 hold394/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout830 fanout843/X vssd1 vssd1 vccd1 vccd1 _14863_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout841 _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14877_/C1 sky130_fd_sc_hd__buf_4
Xfanout852 _17754_/Q vssd1 vssd1 vccd1 vccd1 _11203_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09939_ _09981_/A _09939_/B vssd1 vssd1 vccd1 vccd1 _09939_/X sky130_fd_sc_hd__or2_1
Xfanout863 _15161_/A vssd1 vssd1 vccd1 vccd1 _15541_/A sky130_fd_sc_hd__buf_12
Xfanout874 _07780_/Y vssd1 vssd1 vccd1 vccd1 _14952_/A sky130_fd_sc_hd__buf_12
Xfanout885 _15195_/A vssd1 vssd1 vccd1 vccd1 _15521_/A sky130_fd_sc_hd__clkbuf_16
X_12950_ hold4015/X _12949_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12951_/B sky130_fd_sc_hd__mux2_1
Xfanout896 _14974_/A vssd1 vssd1 vccd1 vccd1 _15515_/A sky130_fd_sc_hd__clkbuf_16
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1050 _08296_/X vssd1 vssd1 vccd1 vccd1 _15781_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1061 _14883_/X vssd1 vssd1 vccd1 vccd1 _18230_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ _13797_/A _11901_/B vssd1 vssd1 vccd1 vccd1 _11901_/X sky130_fd_sc_hd__or2_1
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1072 _18277_/Q vssd1 vssd1 vccd1 vccd1 hold1072/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1083 _07901_/X vssd1 vssd1 vccd1 vccd1 _15594_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ hold3152/X _12880_/X _12905_/S vssd1 vssd1 vccd1 vccd1 _12881_/X sky130_fd_sc_hd__mux2_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1094 _13940_/X vssd1 vssd1 vccd1 vccd1 _13941_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_375_wb_clk_i clkbuf_6_32_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17728_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14620_ _15229_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14620_/X sky130_fd_sc_hd__or2_1
X_11832_ _12216_/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11832_/X sky130_fd_sc_hd__or2_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_304_wb_clk_i clkbuf_6_44_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17832_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14551_ _15231_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14551_/X sky130_fd_sc_hd__or2_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11763_ hold4393/X _12243_/A _11762_/X vssd1 vssd1 vccd1 vccd1 _11763_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ hold5551/X _11213_/B _10713_/X _14342_/A vssd1 vssd1 vccd1 vccd1 _10714_/X
+ sky130_fd_sc_hd__o211a_1
X_13502_ hold2340/X _17621_/Q _13877_/C vssd1 vssd1 vccd1 vccd1 _13503_/B sky130_fd_sc_hd__mux2_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14482_ hold2693/X _14481_/B _14481_/Y _14350_/A vssd1 vssd1 vccd1 vccd1 _14482_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ _17270_/CLK _17270_/D vssd1 vssd1 vccd1 vccd1 _17270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11694_ _11694_/A _11694_/B vssd1 vssd1 vccd1 vccd1 _11694_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13433_ hold1052/X _17598_/Q _13766_/S vssd1 vssd1 vccd1 vccd1 _13434_/B sky130_fd_sc_hd__mux2_1
X_16221_ _17452_/CLK _16221_/D vssd1 vssd1 vccd1 vccd1 _16221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10645_ _11218_/A _10645_/B vssd1 vssd1 vccd1 vccd1 _10645_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_125_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16152_ _17492_/CLK _16152_/D vssd1 vssd1 vccd1 vccd1 _16152_/Q sky130_fd_sc_hd__dfxtp_1
X_13364_ hold1430/X hold4303/X _13886_/C vssd1 vssd1 vccd1 vccd1 _13365_/B sky130_fd_sc_hd__mux2_1
X_10576_ _11206_/A _10576_/B vssd1 vssd1 vccd1 vccd1 _16682_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_224_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15103_ _15103_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15103_/X sky130_fd_sc_hd__or2_1
X_12315_ hold4267/X _13482_/A _12314_/X vssd1 vssd1 vccd1 vccd1 _12315_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_210_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16083_ _17291_/CLK _16083_/D vssd1 vssd1 vccd1 vccd1 hold807/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_239_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13295_ _13311_/A1 _13293_/X _13294_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13295_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15034_ _15473_/A _15034_/B vssd1 vssd1 vccd1 vccd1 _18302_/D sky130_fd_sc_hd__and2_1
XFILLER_0_121_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12246_ _12273_/A _12246_/B vssd1 vssd1 vccd1 vccd1 _12246_/X sky130_fd_sc_hd__or2_1
XFILLER_0_224_1278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_91_wb_clk_i clkbuf_6_17_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18404_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_139_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12177_ _13407_/A _12177_/B vssd1 vssd1 vccd1 vccd1 _12177_/X sky130_fd_sc_hd__or2_1
XFILLER_0_208_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_wb_clk_i clkbuf_6_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17468_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11128_ hold4807/X _11222_/B _11127_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _11128_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16985_ _17894_/CLK _16985_/D vssd1 vssd1 vccd1 vccd1 _16985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15936_ _17345_/CLK _15936_/D vssd1 vssd1 vccd1 vccd1 _15936_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11059_ hold4889/X _11153_/B _11058_/X _14354_/A vssd1 vssd1 vccd1 vccd1 _11059_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15867_ _17738_/CLK _15867_/D vssd1 vssd1 vccd1 vccd1 _15867_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_231_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17606_ _17606_/CLK _17606_/D vssd1 vssd1 vccd1 vccd1 _17606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14818_ _15103_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14818_/X sky130_fd_sc_hd__or2_1
XFILLER_0_231_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15798_ _17697_/CLK _15798_/D vssd1 vssd1 vccd1 vccd1 _15798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17537_ _18372_/CLK _17537_/D vssd1 vssd1 vccd1 vccd1 _17537_/Q sky130_fd_sc_hd__dfxtp_1
X_14749_ hold1839/X _14772_/B _14748_/X _14853_/C1 vssd1 vssd1 vccd1 vccd1 _14749_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08270_ _15549_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08270_/X sky130_fd_sc_hd__or2_1
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17468_ _17468_/CLK _17468_/D vssd1 vssd1 vccd1 vccd1 _17468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16419_ _18390_/CLK _16419_/D vssd1 vssd1 vccd1 vccd1 _16419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17399_ _18451_/CLK _17399_/D vssd1 vssd1 vccd1 vccd1 _17399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6006 _17548_/Q vssd1 vssd1 vccd1 vccd1 hold6006/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6017 _17537_/Q vssd1 vssd1 vccd1 vccd1 hold6017/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6028 _17534_/Q vssd1 vssd1 vccd1 vccd1 hold6028/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6039 data_in[26] vssd1 vssd1 vccd1 vccd1 hold312/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5305 _17185_/Q vssd1 vssd1 vccd1 vccd1 hold5305/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5316 _11548_/X vssd1 vssd1 vccd1 vccd1 _17006_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5327 _16806_/Q vssd1 vssd1 vccd1 vccd1 hold5327/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5338 _13594_/X vssd1 vssd1 vccd1 vccd1 _17651_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4604 _16394_/Q vssd1 vssd1 vccd1 vccd1 hold4604/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5349 _16987_/Q vssd1 vssd1 vccd1 vccd1 hold5349/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4615 _10945_/X vssd1 vssd1 vccd1 vccd1 _16805_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4626 _16673_/Q vssd1 vssd1 vccd1 vccd1 hold4626/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4637 _11736_/Y vssd1 vssd1 vccd1 vccd1 _11737_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3903 _16416_/Q vssd1 vssd1 vccd1 vccd1 hold3903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4648 _16500_/Q vssd1 vssd1 vccd1 vccd1 hold4648/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3914 _10210_/X vssd1 vssd1 vccd1 vccd1 _16560_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4659 _13699_/X vssd1 vssd1 vccd1 vccd1 _17686_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3925 _16384_/Q vssd1 vssd1 vccd1 vccd1 hold3925/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3936 _11926_/X vssd1 vssd1 vccd1 vccd1 _17132_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_240_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3947 _09553_/X vssd1 vssd1 vccd1 vccd1 _16341_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3958 _16866_/Q vssd1 vssd1 vccd1 vccd1 hold3958/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3969 _17411_/Q vssd1 vssd1 vccd1 vccd1 hold3969/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout148 _12812_/S vssd1 vssd1 vccd1 vccd1 _12839_/S sky130_fd_sc_hd__buf_6
Xfanout159 hold2272/X vssd1 vssd1 vccd1 vccd1 _12905_/S sky130_fd_sc_hd__buf_4
X_07985_ hold2453/X _07978_/B _07984_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _07985_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09724_ hold5821/X _10022_/B _09723_/X _15202_/C1 vssd1 vssd1 vccd1 vccd1 _09724_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_241_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_236_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09655_ hold3860/X _10049_/B _09654_/X _15146_/C1 vssd1 vssd1 vccd1 vccd1 _09655_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08606_ _09440_/B hold887/X vssd1 vssd1 vccd1 vccd1 _15925_/D sky130_fd_sc_hd__and2_1
XFILLER_0_167_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09586_ hold3925/X _10568_/B _09585_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _09586_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08537_ _15314_/A hold736/X vssd1 vssd1 vccd1 vccd1 _15892_/D sky130_fd_sc_hd__and2_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08468_ _14413_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08468_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_231_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08399_ _15513_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08399_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10430_ hold1265/X _16634_/Q _10640_/C vssd1 vssd1 vccd1 vccd1 _10431_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10361_ hold2743/X hold3326/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10362_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12100_ hold4803/X _12308_/B _12099_/X _08167_/A vssd1 vssd1 vccd1 vccd1 _12100_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5850 output91/X vssd1 vssd1 vccd1 vccd1 data_out[27] sky130_fd_sc_hd__buf_12
X_13080_ _13073_/X _13079_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17528_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_104_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5861 hold6014/X vssd1 vssd1 vccd1 vccd1 _13153_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10292_ hold1986/X _16588_/Q _10625_/C vssd1 vssd1 vccd1 vccd1 _10293_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5872 output73/X vssd1 vssd1 vccd1 vccd1 data_out[10] sky130_fd_sc_hd__buf_12
XFILLER_0_237_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5883 hold6026/X vssd1 vssd1 vccd1 vccd1 _13209_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5894 output83/X vssd1 vssd1 vccd1 vccd1 data_out[1] sky130_fd_sc_hd__buf_12
XFILLER_0_44_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12031_ hold5295/X _12317_/B _12030_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _12031_/X
+ sky130_fd_sc_hd__o211a_1
Xhold180 hold11/X vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold191 hold676/X vssd1 vssd1 vccd1 vccd1 hold677/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_218_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout660 _12588_/A vssd1 vssd1 vccd1 vccd1 _15506_/A sky130_fd_sc_hd__buf_4
Xfanout671 _08351_/A vssd1 vssd1 vccd1 vccd1 _13795_/C1 sky130_fd_sc_hd__buf_2
XFILLER_0_232_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout682 fanout689/X vssd1 vssd1 vccd1 vccd1 _14356_/A sky130_fd_sc_hd__buf_2
X_16770_ _18005_/CLK _16770_/D vssd1 vssd1 vccd1 vccd1 _16770_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout693 _15284_/A vssd1 vssd1 vccd1 vccd1 _15244_/A sky130_fd_sc_hd__clkbuf_4
X_13982_ _15163_/A _13986_/B vssd1 vssd1 vccd1 vccd1 _13982_/Y sky130_fd_sc_hd__nand2_1
X_15721_ _17190_/CLK _15721_/D vssd1 vssd1 vccd1 vccd1 _15721_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ _12987_/A _12933_/B vssd1 vssd1 vccd1 vccd1 _17487_/D sky130_fd_sc_hd__and2_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_35_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_35_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_18440_ _18455_/CLK _18440_/D vssd1 vssd1 vccd1 vccd1 _18440_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _17259_/CLK _15652_/D vssd1 vssd1 vccd1 vccd1 _15652_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _12864_/A _12864_/B vssd1 vssd1 vccd1 vccd1 _17464_/D sky130_fd_sc_hd__and2_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ hold1976/X _14610_/B _14602_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14603_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ _18371_/CLK _18371_/D vssd1 vssd1 vccd1 vccd1 _18371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11815_ hold5099/X _12293_/B _11814_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _11815_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12795_ _12798_/A _12795_/B vssd1 vssd1 vccd1 vccd1 _17441_/D sky130_fd_sc_hd__and2_1
X_15583_ _17749_/CLK _15583_/D vssd1 vssd1 vccd1 vccd1 _15583_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _17322_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 _17322_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14534_ hold2086/X _14537_/B _14533_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _14534_/X
+ sky130_fd_sc_hd__o211a_1
X_11746_ _12301_/A _11746_/B vssd1 vssd1 vccd1 vccd1 _17072_/D sky130_fd_sc_hd__nor2_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17253_ _17264_/CLK _17253_/D vssd1 vssd1 vccd1 vccd1 _17253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14465_ _15199_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14465_/X sky130_fd_sc_hd__or2_1
X_11677_ hold5701/X _11771_/B _11676_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _11677_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16204_ _17435_/CLK _16204_/D vssd1 vssd1 vccd1 vccd1 _16204_/Q sky130_fd_sc_hd__dfxtp_1
X_10628_ _16700_/Q _10628_/B _10628_/C vssd1 vssd1 vccd1 vccd1 _10628_/X sky130_fd_sc_hd__and3_1
X_13416_ _13800_/A _13416_/B vssd1 vssd1 vccd1 vccd1 _13416_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14396_ hold1927/X _14446_/A2 _14395_/X _14462_/C1 vssd1 vssd1 vccd1 vccd1 _14396_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17184_ _17280_/CLK _17184_/D vssd1 vssd1 vccd1 vccd1 _17184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16135_ _16139_/CLK _16135_/D vssd1 vssd1 vccd1 vccd1 hold760/A sky130_fd_sc_hd__dfxtp_1
X_13347_ _13737_/A _13347_/B vssd1 vssd1 vccd1 vccd1 _13347_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10559_ hold1829/X hold3243/X _10601_/C vssd1 vssd1 vccd1 vccd1 _10560_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_52_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13278_ _13278_/A _13294_/B vssd1 vssd1 vccd1 vccd1 _13278_/X sky130_fd_sc_hd__or2_1
X_16066_ _18417_/CLK _16066_/D vssd1 vssd1 vccd1 vccd1 hold561/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15017_ hold6084/X _15004_/B hold200/X _15212_/C1 vssd1 vssd1 vccd1 vccd1 hold201/A
+ sky130_fd_sc_hd__o211a_1
X_12229_ _12323_/A _12356_/B _12228_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _12229_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2509 _15657_/Q vssd1 vssd1 vccd1 vccd1 hold2509/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1808 _09409_/X vssd1 vssd1 vccd1 vccd1 _16290_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1819 _15867_/Q vssd1 vssd1 vccd1 vccd1 hold1819/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_297_wb_clk_i clkbuf_6_39_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17862_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_224_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16968_ _18429_/CLK _16968_/D vssd1 vssd1 vccd1 vccd1 _16968_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_226_wb_clk_i clkbuf_6_63_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18125_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15919_ _16086_/CLK _15919_/D vssd1 vssd1 vccd1 vccd1 hold599/A sky130_fd_sc_hd__dfxtp_1
X_16899_ _18070_/CLK _16899_/D vssd1 vssd1 vccd1 vccd1 _16899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09440_ _18463_/A _09440_/B vssd1 vssd1 vccd1 vccd1 _09484_/B sky130_fd_sc_hd__and2_1
XFILLER_0_204_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09371_ hold863/X _15486_/B1 _09386_/D hold694/X _09370_/X vssd1 vssd1 vccd1 vccd1
+ _09375_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_149_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08322_ hold2357/X _08323_/B _08321_/Y _12738_/A vssd1 vssd1 vccd1 vccd1 _08322_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08253_ hold1404/X _08262_/B _08252_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _08253_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08184_ hold2322/X _08209_/B _08183_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _08184_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5102 _13384_/X vssd1 vssd1 vccd1 vccd1 _17581_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_1362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5113 _17043_/Q vssd1 vssd1 vccd1 vccd1 hold5113/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5124 _12121_/X vssd1 vssd1 vccd1 vccd1 _17197_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5135 _17074_/Q vssd1 vssd1 vccd1 vccd1 hold5135/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5146 _16554_/Q vssd1 vssd1 vccd1 vccd1 hold5146/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4401 _11209_/Y vssd1 vssd1 vccd1 vccd1 _16893_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5157 _16819_/Q vssd1 vssd1 vccd1 vccd1 hold5157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4412 _11796_/Y vssd1 vssd1 vccd1 vccd1 _11797_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4423 _13855_/Y vssd1 vssd1 vccd1 vccd1 _17738_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5168 _12178_/X vssd1 vssd1 vccd1 vccd1 _17216_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4434 _12336_/Y vssd1 vssd1 vccd1 vccd1 _12337_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3700 _16571_/Q vssd1 vssd1 vccd1 vccd1 hold3700/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5179 _17176_/Q vssd1 vssd1 vccd1 vccd1 hold5179/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4445 _17486_/Q vssd1 vssd1 vccd1 vccd1 hold4445/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3711 _10528_/X vssd1 vssd1 vccd1 vccd1 _16666_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4456 _16604_/Q vssd1 vssd1 vccd1 vccd1 hold4456/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4467 _17490_/Q vssd1 vssd1 vccd1 vccd1 hold4467/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3722 _17412_/Q vssd1 vssd1 vccd1 vccd1 hold3722/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3733 _09883_/X vssd1 vssd1 vccd1 vccd1 _16451_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4478 _12518_/X vssd1 vssd1 vccd1 vccd1 _12519_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3744 _16448_/Q vssd1 vssd1 vccd1 vccd1 hold3744/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4489 _13884_/Y vssd1 vssd1 vccd1 vccd1 _13885_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3755 _16440_/Q vssd1 vssd1 vccd1 vccd1 hold3755/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3766 _10513_/X vssd1 vssd1 vccd1 vccd1 _16661_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3777 _16423_/Q vssd1 vssd1 vccd1 vccd1 hold3777/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3788 _16925_/Q vssd1 vssd1 vccd1 vccd1 hold3788/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3799 _16573_/Q vssd1 vssd1 vccd1 vccd1 hold3799/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07968_ _15537_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07968_/X sky130_fd_sc_hd__or2_1
X_09707_ hold2561/X hold3694/X _10004_/C vssd1 vssd1 vccd1 vccd1 _09708_/B sky130_fd_sc_hd__mux2_1
X_07899_ hold2537/X _07924_/B _07898_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _07899_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09638_ hold2187/X _16370_/Q _11171_/C vssd1 vssd1 vccd1 vccd1 _09639_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09569_ hold2875/X _16347_/Q _10475_/S vssd1 vssd1 vccd1 vccd1 _09570_/B sky130_fd_sc_hd__mux2_1
X_11600_ hold2167/X _17024_/Q _12335_/C vssd1 vssd1 vccd1 vccd1 _11601_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_183_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12580_ hold2159/X hold3365/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12580_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11531_ hold3012/X hold5368/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11532_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14250_ _15199_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14250_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11462_ hold2324/X _16978_/Q _11753_/C vssd1 vssd1 vccd1 vccd1 _11463_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_163_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13201_ _13201_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13201_/X sky130_fd_sc_hd__and2_1
XFILLER_0_208_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10413_ _10413_/A _10413_/B vssd1 vssd1 vccd1 vccd1 _10413_/X sky130_fd_sc_hd__or2_1
XFILLER_0_184_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14181_ hold2248/X _14202_/B _14180_/X _14346_/A vssd1 vssd1 vccd1 vccd1 _14181_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11393_ hold2639/X hold5138/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11394_/B sky130_fd_sc_hd__mux2_1
X_13132_ hold4281/X _13131_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13132_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_103_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10344_ _10536_/A _10344_/B vssd1 vssd1 vccd1 vccd1 _10344_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13063_ _13199_/A1 _13061_/X _13062_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13063_/X
+ sky130_fd_sc_hd__o211a_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5680 _11581_/X vssd1 vssd1 vccd1 vccd1 _17017_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17940_ _18069_/CLK _17940_/D vssd1 vssd1 vccd1 vccd1 _17940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10275_ _10530_/A _10275_/B vssd1 vssd1 vccd1 vccd1 _10275_/X sky130_fd_sc_hd__or2_1
Xhold5691 _16936_/Q vssd1 vssd1 vccd1 vccd1 hold5691/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12014_ hold1303/X hold4787/X _12293_/C vssd1 vssd1 vccd1 vccd1 _12015_/B sky130_fd_sc_hd__mux2_1
Xhold4990 _11473_/X vssd1 vssd1 vccd1 vccd1 _16981_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17871_ _17871_/CLK _17871_/D vssd1 vssd1 vccd1 vccd1 _17871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_219_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_390_wb_clk_i clkbuf_6_38_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17107_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16822_ _17929_/CLK _16822_/D vssd1 vssd1 vccd1 vccd1 _16822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_217_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout490 _09992_/C vssd1 vssd1 vccd1 vccd1 _10022_/C sky130_fd_sc_hd__clkbuf_8
X_16753_ _17967_/CLK _16753_/D vssd1 vssd1 vccd1 vccd1 _16753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13965_ hold3059/X _13995_/A2 _13964_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _13965_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_232_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15704_ _17154_/CLK _15704_/D vssd1 vssd1 vccd1 vccd1 _15704_/Q sky130_fd_sc_hd__dfxtp_1
X_12916_ hold1626/X _17483_/Q _12916_/S vssd1 vssd1 vccd1 vccd1 _12916_/X sky130_fd_sc_hd__mux2_1
X_16684_ _18146_/CLK _16684_/D vssd1 vssd1 vccd1 vccd1 _16684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13896_ _14970_/A hold2055/X hold297/X vssd1 vssd1 vccd1 vccd1 _13897_/B sky130_fd_sc_hd__mux2_1
X_18423_ _18423_/CLK _18423_/D vssd1 vssd1 vccd1 vccd1 _18423_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_201_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15635_ _17899_/CLK _15635_/D vssd1 vssd1 vccd1 vccd1 _15635_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ hold1622/X hold3149/X _12850_/S vssd1 vssd1 vccd1 vccd1 _12847_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_158_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _18380_/CLK _18354_/D vssd1 vssd1 vccd1 vccd1 _18354_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ _17262_/CLK _15566_/D vssd1 vssd1 vccd1 vccd1 _15566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12778_ hold3000/X hold4036/X _12838_/S vssd1 vssd1 vccd1 vccd1 _12778_/X sky130_fd_sc_hd__mux2_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _17320_/CLK _17305_/D vssd1 vssd1 vccd1 vccd1 hold410/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14517_ _14517_/A _14543_/B vssd1 vssd1 vccd1 vccd1 _14517_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18285_ _18387_/CLK _18285_/D vssd1 vssd1 vccd1 vccd1 _18285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11729_ _17067_/Q _11732_/B _11732_/C vssd1 vssd1 vccd1 vccd1 _11729_/X sky130_fd_sc_hd__and3_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15497_ _14972_/A hold1710/X _15505_/S vssd1 vssd1 vccd1 vccd1 _15497_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17236_ _17236_/CLK _17236_/D vssd1 vssd1 vccd1 vccd1 _17236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14448_ _15128_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14479_/B sky130_fd_sc_hd__or2_4
XFILLER_0_181_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17167_ _17167_/CLK _17167_/D vssd1 vssd1 vccd1 vccd1 _17167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold905 hold905/A vssd1 vssd1 vccd1 vccd1 hold905/X sky130_fd_sc_hd__buf_1
XFILLER_0_25_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14379_ hold97/X _17989_/Q _14381_/S vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__mux2_1
Xhold916 hold916/A vssd1 vssd1 vccd1 vccd1 hold916/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold927 hold927/A vssd1 vssd1 vccd1 vccd1 hold927/X sky130_fd_sc_hd__buf_12
X_16118_ _17341_/CLK _16118_/D vssd1 vssd1 vccd1 vccd1 _16118_/Q sky130_fd_sc_hd__dfxtp_1
Xhold938 hold938/A vssd1 vssd1 vccd1 vccd1 hold938/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold949 hold965/X vssd1 vssd1 vccd1 vccd1 hold966/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17098_ _17127_/CLK _17098_/D vssd1 vssd1 vccd1 vccd1 _17098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3007 _14183_/X vssd1 vssd1 vccd1 vccd1 _17894_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16049_ _16129_/CLK _16049_/D vssd1 vssd1 vccd1 vccd1 _16049_/Q sky130_fd_sc_hd__dfxtp_1
X_08940_ _12412_/A hold664/X vssd1 vssd1 vccd1 vccd1 _16087_/D sky130_fd_sc_hd__and2_1
Xhold3018 _14536_/X vssd1 vssd1 vccd1 vccd1 _18064_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3029 _16270_/Q vssd1 vssd1 vccd1 vccd1 hold3029/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2306 _18393_/Q vssd1 vssd1 vccd1 vccd1 hold2306/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_407_wb_clk_i clkbuf_6_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17867_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08871_ _15244_/A hold648/X vssd1 vssd1 vccd1 vccd1 _16053_/D sky130_fd_sc_hd__and2_1
Xhold2317 _14512_/X vssd1 vssd1 vccd1 vccd1 _18052_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2328 _18026_/Q vssd1 vssd1 vccd1 vccd1 hold2328/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2339 _08028_/X vssd1 vssd1 vccd1 vccd1 _15655_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1605 _07987_/X vssd1 vssd1 vccd1 vccd1 _15636_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07822_ hold235/X hold220/X vssd1 vssd1 vccd1 vccd1 _09496_/A sky130_fd_sc_hd__or2_1
Xhold1616 _18060_/Q vssd1 vssd1 vccd1 vccd1 hold1616/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1627 _09173_/X vssd1 vssd1 vccd1 vccd1 _16199_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1638 _08508_/X vssd1 vssd1 vccd1 vccd1 _15881_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1649 _15126_/X vssd1 vssd1 vccd1 vccd1 _18347_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09423_ _07804_/A _09463_/A _08851_/A _09422_/X vssd1 vssd1 vccd1 vccd1 _09423_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09354_ _09366_/A _09366_/B _09361_/C vssd1 vssd1 vccd1 vccd1 _09354_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_192_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08305_ _15203_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08305_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09285_ hold406/X hold363/A vssd1 vssd1 vccd1 vccd1 _09285_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_75_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08236_ _14850_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08236_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08167_ _08167_/A _08167_/B vssd1 vssd1 vccd1 vccd1 _15721_/D sky130_fd_sc_hd__and2_1
XFILLER_0_15_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08098_ _15557_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08098_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4220 _15433_/X vssd1 vssd1 vccd1 vccd1 _15434_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4231 _13827_/Y vssd1 vssd1 vccd1 vccd1 _13828_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4242 _17567_/Q vssd1 vssd1 vccd1 vccd1 hold4242/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4253 _11173_/Y vssd1 vssd1 vccd1 vccd1 _16881_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4264 _16341_/Q vssd1 vssd1 vccd1 vccd1 _13198_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_148_wb_clk_i clkbuf_6_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18398_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold3530 _17435_/Q vssd1 vssd1 vccd1 vccd1 hold3530/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4275 _12355_/Y vssd1 vssd1 vccd1 vccd1 _17275_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3541 _16511_/Q vssd1 vssd1 vccd1 vccd1 hold3541/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10060_ _11206_/A _10060_/B vssd1 vssd1 vccd1 vccd1 _10060_/Y sky130_fd_sc_hd__nor2_1
Xhold4286 _11164_/Y vssd1 vssd1 vccd1 vccd1 _16878_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3552 _16383_/Q vssd1 vssd1 vccd1 vccd1 hold3552/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4297 _11800_/Y vssd1 vssd1 vccd1 vccd1 _17090_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3563 _09670_/X vssd1 vssd1 vccd1 vccd1 _16380_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3574 _16461_/Q vssd1 vssd1 vccd1 vccd1 hold3574/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3585 _09691_/X vssd1 vssd1 vccd1 vccd1 _16387_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2840 _15596_/Q vssd1 vssd1 vccd1 vccd1 hold2840/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3596 _10078_/X vssd1 vssd1 vccd1 vccd1 _16516_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2851 _14321_/X vssd1 vssd1 vccd1 vccd1 _17960_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2862 _08255_/X vssd1 vssd1 vccd1 vccd1 _15762_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2873 _17813_/Q vssd1 vssd1 vccd1 vccd1 hold2873/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2884 _17836_/Q vssd1 vssd1 vccd1 vccd1 hold2884/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2895 _15870_/Q vssd1 vssd1 vccd1 vccd1 hold2895/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10962_ _11136_/A _10962_/B vssd1 vssd1 vccd1 vccd1 _10962_/X sky130_fd_sc_hd__or2_1
X_13750_ hold5478/X _12374_/B _13749_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _13750_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12701_ hold3793/X _12700_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12701_/X sky130_fd_sc_hd__mux2_1
X_10893_ _11091_/A _10893_/B vssd1 vssd1 vccd1 vccd1 _10893_/X sky130_fd_sc_hd__or2_1
X_13681_ hold5378/X _13871_/B _13680_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13681_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15420_ _15983_/Q _09365_/B _09362_/D hold665/X _15418_/X vssd1 vssd1 vccd1 vccd1
+ _15422_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_128_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12632_ hold3139/X _12631_/X _12851_/S vssd1 vssd1 vccd1 vccd1 _12632_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_167_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15351_ _16299_/Q _09362_/A _09392_/B hold663/X _15350_/X vssd1 vssd1 vccd1 vccd1
+ _15352_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_148_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12563_ hold4999/X _12562_/X _12929_/S vssd1 vssd1 vccd1 vccd1 _12564_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_136_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14302_ hold933/X _14338_/B vssd1 vssd1 vccd1 vccd1 _14302_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ _11697_/A _11514_/B vssd1 vssd1 vccd1 vccd1 _11514_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_227_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18070_ _18070_/CLK _18070_/D vssd1 vssd1 vccd1 vccd1 _18070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12494_ _17340_/Q _12506_/B vssd1 vssd1 vccd1 vccd1 _12494_/X sky130_fd_sc_hd__or2_1
X_15282_ _15489_/A _15282_/B _15282_/C _15282_/D vssd1 vssd1 vccd1 vccd1 _15282_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_124_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17021_ _17901_/CLK _17021_/D vssd1 vssd1 vccd1 vccd1 _17021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11445_ _11637_/A _11445_/B vssd1 vssd1 vccd1 vccd1 _11445_/X sky130_fd_sc_hd__or2_1
X_14233_ hold406/X _14502_/B vssd1 vssd1 vccd1 vccd1 _14282_/B sky130_fd_sc_hd__or2_4
XFILLER_0_123_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14164_ _14164_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14164_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11376_ _11670_/A _11376_/B vssd1 vssd1 vccd1 vccd1 _11376_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10327_ hold3308/X _10637_/B _10326_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _10327_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13115_ _13114_/X hold4345/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13115_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_238_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14095_ hold2555/X _14094_/B _14094_/Y _13897_/A vssd1 vssd1 vccd1 vccd1 _14095_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_237_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _17523_/Q hold907/X _13046_/C _13046_/D vssd1 vssd1 vccd1 vccd1 _13046_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_221_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17923_ _18039_/CLK hold652/X vssd1 vssd1 vccd1 vccd1 hold651/A sky130_fd_sc_hd__dfxtp_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ hold4594/X _10646_/B _10257_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10258_/X
+ sky130_fd_sc_hd__o211a_1
X_17854_ _17886_/CLK _17854_/D vssd1 vssd1 vccd1 vccd1 _17854_/Q sky130_fd_sc_hd__dfxtp_1
X_10189_ hold3292/X _10571_/B _10188_/X _14769_/C1 vssd1 vssd1 vccd1 vccd1 _10189_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16805_ _18072_/CLK _16805_/D vssd1 vssd1 vccd1 vccd1 _16805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17785_ _18432_/CLK _17785_/D vssd1 vssd1 vccd1 vccd1 _17785_/Q sky130_fd_sc_hd__dfxtp_1
X_14997_ hold1827/X _15004_/B _14996_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _14997_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16736_ _18067_/CLK _16736_/D vssd1 vssd1 vccd1 vccd1 _16736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13948_ _14164_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13948_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16667_ _18225_/CLK _16667_/D vssd1 vssd1 vccd1 vccd1 _16667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13879_ _13888_/A _13879_/B vssd1 vssd1 vccd1 vccd1 _13879_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_53_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_234_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18406_ _18406_/CLK _18406_/D vssd1 vssd1 vccd1 vccd1 _18406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15618_ _17278_/CLK _15618_/D vssd1 vssd1 vccd1 vccd1 _15618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16598_ _18188_/CLK _16598_/D vssd1 vssd1 vccd1 vccd1 _16598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18337_ _18373_/CLK hold643/X vssd1 vssd1 vccd1 vccd1 _18337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15549_ _15549_/A _15549_/B vssd1 vssd1 vccd1 vccd1 _15549_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09070_ _15511_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09070_/X sky130_fd_sc_hd__or2_1
X_18268_ _18298_/CLK hold409/X vssd1 vssd1 vccd1 vccd1 _18268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08021_ _09313_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08021_/X sky130_fd_sc_hd__or2_1
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17219_ _17749_/CLK _17219_/D vssd1 vssd1 vccd1 vccd1 _17219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18199_ _18218_/CLK _18199_/D vssd1 vssd1 vccd1 vccd1 _18199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold702 hold702/A vssd1 vssd1 vccd1 vccd1 hold702/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 input70/X vssd1 vssd1 vccd1 vccd1 hold713/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold724 hold724/A vssd1 vssd1 vccd1 vccd1 hold724/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 hold735/A vssd1 vssd1 vccd1 vccd1 hold735/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 hold746/A vssd1 vssd1 vccd1 vccd1 hold746/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold757 hold757/A vssd1 vssd1 vccd1 vccd1 hold757/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold768 hold768/A vssd1 vssd1 vccd1 vccd1 hold768/X sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ _10560_/A _09972_/B vssd1 vssd1 vccd1 vccd1 _09972_/X sky130_fd_sc_hd__or2_1
Xhold779 hold779/A vssd1 vssd1 vccd1 vccd1 hold779/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_241_wb_clk_i clkbuf_6_60_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18172_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08923_ _09440_/B _08923_/B vssd1 vssd1 vccd1 vccd1 _16079_/D sky130_fd_sc_hd__and2_1
Xhold2103 hold2227/X vssd1 vssd1 vccd1 vccd1 hold2103/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2114 _14683_/X vssd1 vssd1 vccd1 vccd1 _18133_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2125 _17914_/Q vssd1 vssd1 vccd1 vccd1 hold2125/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_239_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2136 _14741_/X vssd1 vssd1 vccd1 vccd1 _18161_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1402 _17939_/Q vssd1 vssd1 vccd1 vccd1 hold1402/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2147 _17854_/Q vssd1 vssd1 vccd1 vccd1 hold2147/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08854_ hold438/X hold515/X _08866_/S vssd1 vssd1 vccd1 vccd1 _08855_/B sky130_fd_sc_hd__mux2_1
Xhold2158 _15156_/X vssd1 vssd1 vccd1 vccd1 _18361_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1413 _17768_/Q vssd1 vssd1 vccd1 vccd1 hold1413/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1424 _15043_/X vssd1 vssd1 vccd1 vccd1 _15044_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2169 _18211_/Q vssd1 vssd1 vccd1 vccd1 hold2169/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1435 _15208_/X vssd1 vssd1 vccd1 vccd1 _18386_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07805_ _07805_/A vssd1 vssd1 vccd1 vccd1 _07805_/Y sky130_fd_sc_hd__inv_2
Xhold1446 _16160_/Q vssd1 vssd1 vccd1 vccd1 hold1446/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08785_ hold82/X hold154/X _08793_/S vssd1 vssd1 vccd1 vccd1 hold155/A sky130_fd_sc_hd__mux2_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1457 _17804_/Q vssd1 vssd1 vccd1 vccd1 hold1457/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1468 _16175_/Q vssd1 vssd1 vccd1 vccd1 _07788_/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_79_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1479 _18349_/Q vssd1 vssd1 vccd1 vccd1 hold1479/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09406_ _09438_/B _16289_/Q vssd1 vssd1 vccd1 vccd1 _09406_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09337_ _15559_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09337_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09268_ _09272_/A hold598/X vssd1 vssd1 vccd1 vccd1 _16245_/D sky130_fd_sc_hd__and2_1
XFILLER_0_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08219_ _14726_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08219_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09199_ hold6056/X _09214_/B _09198_/X _12810_/A vssd1 vssd1 vccd1 vccd1 hold968/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_329_wb_clk_i clkbuf_6_44_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17247_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11230_ hold4111/X _12305_/B _11229_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11230_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11161_ _11203_/A _11161_/B vssd1 vssd1 vccd1 vccd1 _11161_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_101_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4050 _16996_/Q vssd1 vssd1 vccd1 vccd1 hold4050/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10112_ hold2441/X hold3468/X _10634_/C vssd1 vssd1 vccd1 vccd1 _10113_/B sky130_fd_sc_hd__mux2_1
Xhold4061 _17198_/Q vssd1 vssd1 vccd1 vccd1 hold4061/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4072 _17153_/Q vssd1 vssd1 vccd1 vccd1 hold4072/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11092_ hold4897/X _11186_/B _11091_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _11092_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4083 _17029_/Q vssd1 vssd1 vccd1 vccd1 hold4083/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4094 _11611_/X vssd1 vssd1 vccd1 vccd1 _17027_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3360 _17463_/Q vssd1 vssd1 vccd1 vccd1 hold3360/X sky130_fd_sc_hd__dlygate4sd3_1
X_10043_ _16505_/Q _10049_/B _10385_/S vssd1 vssd1 vccd1 vccd1 _10043_/X sky130_fd_sc_hd__and3_1
XFILLER_0_234_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14920_ _15189_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14920_/X sky130_fd_sc_hd__or2_1
Xhold3371 _12638_/X vssd1 vssd1 vccd1 vccd1 _12639_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3382 _12548_/X vssd1 vssd1 vccd1 vccd1 _12549_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3393 _12797_/X vssd1 vssd1 vccd1 vccd1 _12798_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__buf_2
XTAP_5577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2670 _08318_/X vssd1 vssd1 vccd1 vccd1 _15792_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2681 _18117_/Q vssd1 vssd1 vccd1 vccd1 hold2681/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14851_ hold2727/X hold332/X _14850_/X _15019_/C1 vssd1 vssd1 vccd1 vccd1 _14851_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2692 _07947_/X vssd1 vssd1 vccd1 vccd1 _15616_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13802_ _17721_/Q _13814_/B _13817_/C vssd1 vssd1 vccd1 vccd1 _13802_/X sky130_fd_sc_hd__and3_1
XFILLER_0_215_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1980 _18222_/Q vssd1 vssd1 vccd1 vccd1 hold1980/X sky130_fd_sc_hd__dlygate4sd3_1
X_17570_ _17630_/CLK _17570_/D vssd1 vssd1 vccd1 vccd1 _17570_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14782_ _15229_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14782_/X sky130_fd_sc_hd__or2_1
Xhold1991 _09306_/X vssd1 vssd1 vccd1 vccd1 _16263_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11994_ _13407_/A _11994_/B vssd1 vssd1 vccd1 vccd1 _11994_/X sky130_fd_sc_hd__or2_1
X_16521_ _18206_/CLK _16521_/D vssd1 vssd1 vccd1 vccd1 _16521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13733_ hold2733/X hold4569/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13734_/B sky130_fd_sc_hd__mux2_1
X_10945_ hold4614/X _11153_/B _10944_/X _14552_/C1 vssd1 vssd1 vccd1 vccd1 _10945_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_45_wb_clk_i clkbuf_6_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17949_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16452_ _18379_/CLK _16452_/D vssd1 vssd1 vccd1 vccd1 _16452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13664_ hold2946/X _17675_/Q _13871_/C vssd1 vssd1 vccd1 vccd1 _13665_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10876_ hold4845/X _11162_/B _10875_/X _14372_/A vssd1 vssd1 vccd1 vccd1 _10876_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_213_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15403_ _15490_/A1 _15395_/X _15402_/X _15481_/B1 hold5923/A vssd1 vssd1 vccd1 vccd1
+ _15403_/X sky130_fd_sc_hd__a32o_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12615_ _12924_/A _12615_/B vssd1 vssd1 vccd1 vccd1 _17381_/D sky130_fd_sc_hd__and2_1
X_16383_ _18296_/CLK _16383_/D vssd1 vssd1 vccd1 vccd1 _16383_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13595_ hold2897/X _17652_/Q _13883_/C vssd1 vssd1 vccd1 vccd1 _13596_/B sky130_fd_sc_hd__mux2_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18122_ _18220_/CLK _18122_/D vssd1 vssd1 vccd1 vccd1 _18122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15334_ _15414_/A _15334_/B vssd1 vssd1 vccd1 vccd1 _18409_/D sky130_fd_sc_hd__and2_1
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12546_ _12924_/A _12546_/B vssd1 vssd1 vccd1 vccd1 _17358_/D sky130_fd_sc_hd__and2_1
XFILLER_0_13_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18053_ _18053_/CLK _18053_/D vssd1 vssd1 vccd1 vccd1 _18053_/Q sky130_fd_sc_hd__dfxtp_1
X_15265_ hold325/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15265_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12477_ hold11/X _12445_/A _12445_/B _12476_/X _12438_/A vssd1 vssd1 vccd1 vccd1
+ hold12/A sky130_fd_sc_hd__o311a_1
XFILLER_0_112_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_4 _13068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17004_ _17884_/CLK _17004_/D vssd1 vssd1 vccd1 vccd1 _17004_/Q sky130_fd_sc_hd__dfxtp_1
X_14216_ _14897_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14216_/Y sky130_fd_sc_hd__nor2_2
X_11428_ hold4165/X _11717_/B _11427_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11428_/X
+ sky130_fd_sc_hd__o211a_1
X_15196_ hold1857/X _15219_/B _15195_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _15196_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14147_ hold2553/X _14148_/B _14146_/Y _14147_/C1 vssd1 vssd1 vccd1 vccd1 _14147_/X
+ sky130_fd_sc_hd__o211a_1
X_11359_ hold5565/X _11741_/B _11358_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11359_/X
+ sky130_fd_sc_hd__o211a_1
X_14078_ _15531_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14078_/X sky130_fd_sc_hd__or2_1
XFILLER_0_238_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13029_ hold935/X _13029_/B vssd1 vssd1 vccd1 vccd1 hold936/A sky130_fd_sc_hd__or2_1
XFILLER_0_219_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17906_ _17906_/CLK _17906_/D vssd1 vssd1 vccd1 vccd1 _17906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17837_ _17891_/CLK _17837_/D vssd1 vssd1 vccd1 vccd1 _17837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08570_ hold215/X hold582/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08571_/B sky130_fd_sc_hd__mux2_1
X_17768_ _17874_/CLK _17768_/D vssd1 vssd1 vccd1 vccd1 _17768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16719_ _18019_/CLK _16719_/D vssd1 vssd1 vccd1 vccd1 _16719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17699_ _17731_/CLK _17699_/D vssd1 vssd1 vccd1 vccd1 _17699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09122_ _09122_/A _09400_/B vssd1 vssd1 vccd1 vccd1 _09122_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_130_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ _12412_/A _09053_/B vssd1 vssd1 vccd1 vccd1 _16143_/D sky130_fd_sc_hd__and2_1
XFILLER_0_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08004_ hold2449/X _08033_/B _08003_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _08004_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_422_wb_clk_i clkbuf_6_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17264_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold510 hold510/A vssd1 vssd1 vccd1 vccd1 hold510/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold521 hold521/A vssd1 vssd1 vccd1 vccd1 hold521/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 hold532/A vssd1 vssd1 vccd1 vccd1 hold532/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 hold543/A vssd1 vssd1 vccd1 vccd1 hold543/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold554 hold554/A vssd1 vssd1 vccd1 vccd1 hold554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 hold565/A vssd1 vssd1 vccd1 vccd1 hold565/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 hold576/A vssd1 vssd1 vccd1 vccd1 hold576/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 hold587/A vssd1 vssd1 vccd1 vccd1 hold587/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 hold598/A vssd1 vssd1 vccd1 vccd1 hold598/X sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ hold3588/X _10049_/B _09954_/X _15212_/C1 vssd1 vssd1 vccd1 vccd1 _09955_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_217_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08906_ hold245/X hold501/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08907_/B sky130_fd_sc_hd__mux2_1
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ hold5839/X _10022_/B _09885_/X _15202_/C1 vssd1 vssd1 vccd1 vccd1 _09886_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 _14697_/X vssd1 vssd1 vccd1 vccd1 _18140_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 _14733_/X vssd1 vssd1 vccd1 vccd1 _18158_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1232 _14205_/X vssd1 vssd1 vccd1 vccd1 _17905_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08837_ _15254_/A hold662/X vssd1 vssd1 vccd1 vccd1 _16037_/D sky130_fd_sc_hd__and2_1
Xhold1243 _09290_/X vssd1 vssd1 vccd1 vccd1 _16255_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1254 _14604_/A vssd1 vssd1 vccd1 vccd1 _14194_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_212_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1265 _18192_/Q vssd1 vssd1 vccd1 vccd1 hold1265/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1276 _08077_/X vssd1 vssd1 vccd1 vccd1 _15678_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1287 _15683_/Q vssd1 vssd1 vccd1 vccd1 hold1287/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _15394_/A _08768_/B vssd1 vssd1 vccd1 vccd1 _16004_/D sky130_fd_sc_hd__and2_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1298 _09338_/X vssd1 vssd1 vccd1 vccd1 _16279_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ hold254/X hold263/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08700_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10730_ hold2435/X hold3512/X _11210_/C vssd1 vssd1 vccd1 vccd1 _10731_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_48_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10661_ hold2125/X hold3442/X _11144_/C vssd1 vssd1 vccd1 vccd1 _10662_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_36_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12400_ _15254_/A hold811/X vssd1 vssd1 vccd1 vccd1 _17293_/D sky130_fd_sc_hd__and2_1
XFILLER_0_193_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13380_ _13752_/A _13380_/B vssd1 vssd1 vccd1 vccd1 _13380_/X sky130_fd_sc_hd__or2_1
X_10592_ _16688_/Q _10598_/B _10634_/C vssd1 vssd1 vccd1 vccd1 _10592_/X sky130_fd_sc_hd__and3_1
XFILLER_0_134_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12331_ _12331_/A _12331_/B vssd1 vssd1 vccd1 vccd1 _12331_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_163_wb_clk_i clkbuf_6_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18373_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_161_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15050_ _15050_/A _15050_/B vssd1 vssd1 vccd1 vccd1 _18310_/D sky130_fd_sc_hd__and2_1
X_12262_ hold5301/X _12356_/B _12261_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _12262_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11213_ _16895_/Q _11213_/B _11213_/C vssd1 vssd1 vccd1 vccd1 _11213_/X sky130_fd_sc_hd__and3_1
X_14001_ _14681_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14052_/B sky130_fd_sc_hd__or2_4
XFILLER_0_181_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12193_ hold5076/X _12353_/B _12192_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _12193_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11144_ _16872_/Q _11144_/B _11144_/C vssd1 vssd1 vccd1 vccd1 _11144_/X sky130_fd_sc_hd__and3_1
XFILLER_0_43_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput74 _13145_/A vssd1 vssd1 vccd1 vccd1 output74/X sky130_fd_sc_hd__buf_6
XTAP_6031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput85 _13225_/A vssd1 vssd1 vccd1 vccd1 output85/X sky130_fd_sc_hd__buf_6
XTAP_6042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput96 _13305_/A vssd1 vssd1 vccd1 vccd1 output96/X sky130_fd_sc_hd__buf_6
XTAP_6053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15952_ _17299_/CLK _15952_/D vssd1 vssd1 vccd1 vccd1 hold868/A sky130_fd_sc_hd__dfxtp_1
X_11075_ hold2316/X hold4997/X _11654_/S vssd1 vssd1 vccd1 vccd1 _11076_/B sky130_fd_sc_hd__mux2_1
XTAP_6075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3190 _10054_/Y vssd1 vssd1 vccd1 vccd1 _16508_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10026_ _13182_/A _09912_/A _10025_/X vssd1 vssd1 vccd1 vccd1 _10026_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14903_ hold1913/X _14896_/Y _14902_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _14903_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15883_ _17561_/CLK _15883_/D vssd1 vssd1 vccd1 vccd1 _15883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17622_ _17686_/CLK _17622_/D vssd1 vssd1 vccd1 vccd1 _17622_/Q sky130_fd_sc_hd__dfxtp_1
X_14834_ _15227_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14834_/X sky130_fd_sc_hd__or2_1
XFILLER_0_192_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17553_ _18229_/CLK _17553_/D vssd1 vssd1 vccd1 vccd1 _17553_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ hold1785/X _14772_/B _14764_/X _14769_/C1 vssd1 vssd1 vccd1 vccd1 _14765_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ hold4585/X _12332_/B _11976_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _11977_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16504_ _18385_/CLK _16504_/D vssd1 vssd1 vccd1 vccd1 _16504_/Q sky130_fd_sc_hd__dfxtp_1
X_13716_ _13716_/A _13716_/B vssd1 vssd1 vccd1 vccd1 _13716_/X sky130_fd_sc_hd__or2_1
XFILLER_0_58_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10928_ hold994/X _16800_/Q _11216_/C vssd1 vssd1 vccd1 vccd1 _10929_/B sky130_fd_sc_hd__mux2_1
X_17484_ _17484_/CLK _17484_/D vssd1 vssd1 vccd1 vccd1 _17484_/Q sky130_fd_sc_hd__dfxtp_1
X_14696_ _15197_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14696_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16435_ _18372_/CLK _16435_/D vssd1 vssd1 vccd1 vccd1 _16435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13647_ _13773_/A _13647_/B vssd1 vssd1 vccd1 vccd1 _13647_/X sky130_fd_sc_hd__or2_1
X_10859_ hold2593/X hold3985/X _11144_/C vssd1 vssd1 vccd1 vccd1 _10860_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_184_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _18357_/CLK _16366_/D vssd1 vssd1 vccd1 vccd1 _16366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _13794_/A _13578_/B vssd1 vssd1 vccd1 vccd1 _13578_/X sky130_fd_sc_hd__or2_1
X_18105_ _18181_/CLK _18105_/D vssd1 vssd1 vccd1 vccd1 _18105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15317_ hold138/X _15487_/A2 _15484_/B1 _17315_/Q _15316_/X vssd1 vssd1 vccd1 vccd1
+ _15322_/B sky130_fd_sc_hd__a221o_1
X_12529_ hold1062/X _17354_/Q _12925_/S vssd1 vssd1 vccd1 vccd1 _12529_/X sky130_fd_sc_hd__mux2_1
X_16297_ _16315_/CLK _16297_/D vssd1 vssd1 vccd1 vccd1 _16297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5509 _17137_/Q vssd1 vssd1 vccd1 vccd1 hold5509/X sky130_fd_sc_hd__dlygate4sd3_1
X_18036_ _18036_/CLK _18036_/D vssd1 vssd1 vccd1 vccd1 _18036_/Q sky130_fd_sc_hd__dfxtp_1
X_15248_ _15938_/Q _15484_/A2 _09392_/D hold808/X vssd1 vssd1 vccd1 vccd1 _15248_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4808 _11128_/X vssd1 vssd1 vccd1 vccd1 _16866_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4819 _16796_/Q vssd1 vssd1 vccd1 vccd1 hold4819/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_238_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15179_ _15233_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15179_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout308 _11061_/A vssd1 vssd1 vccd1 vccd1 _09984_/A sky130_fd_sc_hd__buf_4
XFILLER_0_205_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout319 _10539_/A vssd1 vssd1 vccd1 vccd1 _11088_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09740_ hold1470/X hold4545/X _10028_/C vssd1 vssd1 vccd1 vccd1 _09741_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_201_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
.ends

