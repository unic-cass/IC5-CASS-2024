* NGSPICE file created from ascon_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt ascon_wrapper clk io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_oeb[0]
+ io_oeb[10] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[1] io_out[2] rst vccd1 vssd1
XFILLER_0_94_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18869_ _18951_/A _18873_/B vssd1 vssd1 vccd1 vccd1 _18871_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20900_ _26300_/Q _20731_/X hold503/X vssd1 vssd1 vccd1 vccd1 _20903_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21880_ _21880_/A _21880_/B vssd1 vssd1 vccd1 vccd1 _21880_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_179_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20831_ _20831_/A _25898_/Q vssd1 vssd1 vccd1 vccd1 _20836_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_76_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20762_ _21677_/B vssd1 vssd1 vccd1 vccd1 _21676_/B sky130_fd_sc_hd__inv_2
X_23550_ _24942_/S hold449/A _23549_/X vssd1 vssd1 vccd1 vccd1 _23550_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22501_ _22653_/A _22501_/B vssd1 vssd1 vccd1 vccd1 _22501_/X sky130_fd_sc_hd__or2_1
X_23481_ _23469_/X _23480_/X _24949_/S vssd1 vssd1 vccd1 vccd1 _23481_/X sky130_fd_sc_hd__mux2_4
XFILLER_0_169_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20693_ _26294_/Q hold760/X vssd1 vssd1 vccd1 vccd1 _20693_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_64_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22432_ _22561_/A _22432_/B vssd1 vssd1 vccd1 vccd1 _22432_/Y sky130_fd_sc_hd__nand2_1
X_25220_ _25807_/CLK hold712/X vssd1 vssd1 vccd1 vccd1 hold710/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22363_ _22561_/A _22363_/B vssd1 vssd1 vccd1 vccd1 _22363_/Y sky130_fd_sc_hd__nand2_1
X_25151_ _26236_/CLK hold565/X vssd1 vssd1 vccd1 vccd1 hold563/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24102_ hold2226/X hold2124/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24103_/A sky130_fd_sc_hd__mux2_1
X_21314_ _21314_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21314_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_115_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25082_ _26167_/CLK hold980/X vssd1 vssd1 vccd1 vccd1 hold979/A sky130_fd_sc_hd__dfxtp_1
X_22294_ _22292_/X _15839_/B _22293_/Y _14860_/A _21725_/X vssd1 vssd1 vccd1 vccd1
+ _22295_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_20_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24033_ _24033_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24034_/A sky130_fd_sc_hd__and2_1
Xhold340 hold340/A vssd1 vssd1 vccd1 vccd1 hold340/X sky130_fd_sc_hd__dlygate4sd3_1
X_21245_ _21245_/A _21245_/B vssd1 vssd1 vccd1 vccd1 _21675_/C sky130_fd_sc_hd__nand2_2
Xhold351 hold351/A vssd1 vssd1 vccd1 vccd1 hold351/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold362 hold362/A vssd1 vssd1 vccd1 vccd1 hold362/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold373 hold373/A vssd1 vssd1 vccd1 vccd1 hold373/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 hold384/A vssd1 vssd1 vccd1 vccd1 hold384/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21176_ _26310_/Q hold488/X vssd1 vssd1 vccd1 vccd1 _21176_/Y sky130_fd_sc_hd__nand2_1
Xhold395 hold395/A vssd1 vssd1 vccd1 vccd1 hold395/X sky130_fd_sc_hd__dlygate4sd3_1
X_20127_ _20127_/A _20127_/B vssd1 vssd1 vccd1 vccd1 _20128_/A sky130_fd_sc_hd__nand2_1
X_25984_ _26001_/CLK _25984_/D vssd1 vssd1 vccd1 vccd1 _25984_/Q sky130_fd_sc_hd__dfxtp_1
X_24935_ _16168_/B _16177_/Y _24944_/S vssd1 vssd1 vccd1 vccd1 _24935_/X sky130_fd_sc_hd__mux2_1
X_20058_ _25878_/Q _20058_/B _20058_/C vssd1 vssd1 vccd1 vccd1 _20062_/B sky130_fd_sc_hd__nand3b_1
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1040 _12757_/X vssd1 vssd1 vccd1 vccd1 _25003_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 _25527_/Q vssd1 vssd1 vccd1 vccd1 _16539_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1062 _13328_/X vssd1 vssd1 vccd1 vccd1 _25106_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24866_ _24863_/X _24865_/Y _24946_/A vssd1 vssd1 vccd1 vccd1 _24866_/X sky130_fd_sc_hd__mux2_1
Xhold1073 _25124_/Q vssd1 vssd1 vccd1 vccd1 _19047_/B sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ _12840_/X _12878_/X _12827_/X _12879_/X vssd1 vssd1 vccd1 vccd1 _12880_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1084 _16744_/Y vssd1 vssd1 vccd1 vccd1 _25545_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 _25066_/Q vssd1 vssd1 vccd1 vccd1 _17819_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23817_ _23817_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23818_/A sky130_fd_sc_hd__and2_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24797_ _24797_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24798_/A sky130_fd_sc_hd__and2_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14550_ _14548_/Y hold345/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold346/A sky130_fd_sc_hd__a21oi_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23748_ _14752_/B _14761_/B _23754_/S vssd1 vssd1 vccd1 vccd1 _23749_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_56_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13501_ _26218_/Q _13426_/X _13468_/X _13500_/Y vssd1 vssd1 vccd1 vccd1 _13502_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _14479_/Y hold198/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold199/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_181_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23679_ _23679_/A vssd1 vssd1 vccd1 vccd1 _25965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16220_ hold957/X vssd1 vssd1 vccd1 vccd1 _16224_/B sky130_fd_sc_hd__inv_2
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25418_ _25418_/CLK _25418_/D vssd1 vssd1 vccd1 vccd1 _25418_/Q sky130_fd_sc_hd__dfxtp_1
X_13432_ _13522_/A _13430_/X _23629_/B _13431_/X vssd1 vssd1 vccd1 vccd1 _13432_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16151_ _16156_/B _16152_/A vssd1 vssd1 vccd1 vccd1 _16151_/X sky130_fd_sc_hd__or2_1
X_25349_ _26301_/CLK hold307/X vssd1 vssd1 vccd1 vccd1 hold305/A sky130_fd_sc_hd__dfxtp_1
X_13363_ _18961_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13363_/X sky130_fd_sc_hd__or2_1
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15102_ _15089_/A _15084_/A _15084_/B vssd1 vssd1 vccd1 vccd1 _15104_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_133_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16082_ _16097_/B _16082_/B vssd1 vssd1 vccd1 vccd1 _16103_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_134_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13294_ _13207_/X _13292_/X _13192_/X _13293_/X vssd1 vssd1 vccd1 vccd1 _13294_/X
+ sky130_fd_sc_hd__o211a_1
X_15033_ _15033_/A _15033_/B vssd1 vssd1 vccd1 vccd1 _15037_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19910_ _20043_/A _22692_/B _25644_/Q vssd1 vssd1 vccd1 vccd1 _20048_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_32_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19841_ _26264_/Q hold521/X vssd1 vssd1 vccd1 vccd1 _19841_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16984_ _20023_/B _25838_/Q _25774_/Q vssd1 vssd1 vccd1 vccd1 _16985_/B sky130_fd_sc_hd__mux2_2
X_19772_ _19771_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19773_/B
+ sky130_fd_sc_hd__a211o_1
X_15935_ _15940_/B _15936_/A vssd1 vssd1 vccd1 vccd1 _15935_/X sky130_fd_sc_hd__or2_1
XFILLER_0_155_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18723_ _18721_/Y _18722_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25680_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18654_ _20370_/B _22350_/A vssd1 vssd1 vccd1 vccd1 _20361_/A sky130_fd_sc_hd__nand2_2
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15866_ _15866_/A _15866_/B vssd1 vssd1 vccd1 vccd1 _15867_/B sky130_fd_sc_hd__nand2_1
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14817_ _22144_/B _15778_/B vssd1 vssd1 vccd1 vccd1 _14818_/A sky130_fd_sc_hd__nand2_1
X_17605_ _17605_/A _17605_/B vssd1 vssd1 vccd1 vccd1 _17605_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_87_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18585_ _18585_/A _18585_/B vssd1 vssd1 vccd1 vccd1 _22266_/A sky130_fd_sc_hd__nand2_1
X_15797_ hold902/X vssd1 vssd1 vccd1 vccd1 _15799_/A sky130_fd_sc_hd__inv_2
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17536_ _17624_/A _17536_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17536_/X sky130_fd_sc_hd__and3_1
X_14748_ _25843_/Q _13466_/A _14747_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14749_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17467_ _17467_/A _17467_/B vssd1 vssd1 vccd1 vccd1 _17467_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_104_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14679_ _14688_/A hold350/X vssd1 vssd1 vccd1 vccd1 hold351/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16418_ _16394_/A _16440_/B _16417_/Y vssd1 vssd1 vccd1 vccd1 _16420_/A sky130_fd_sc_hd__a21bo_1
X_19206_ _19206_/A _20468_/B vssd1 vssd1 vccd1 vccd1 _19206_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_89_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17398_ _25619_/Q vssd1 vssd1 vccd1 vccd1 _21265_/B sky130_fd_sc_hd__inv_2
XFILLER_0_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19137_ _19137_/A vssd1 vssd1 vccd1 vccd1 _19138_/C sky130_fd_sc_hd__inv_2
X_16349_ _16331_/B _16331_/A _16341_/C vssd1 vssd1 vccd1 vccd1 _16351_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19068_ _19082_/A _19068_/B _22786_/A vssd1 vssd1 vccd1 vccd1 _19068_/X sky130_fd_sc_hd__and3_1
XFILLER_0_11_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18019_ _18019_/A _18019_/B vssd1 vssd1 vccd1 vccd1 _18020_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_125_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21030_ _21548_/B vssd1 vssd1 vccd1 vccd1 _21545_/C sky130_fd_sc_hd__inv_2
XFILLER_0_61_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22981_ _26071_/Q vssd1 vssd1 vccd1 vccd1 _22982_/A sky130_fd_sc_hd__inv_2
X_24720_ _24720_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24721_/A sky130_fd_sc_hd__and2_1
X_21932_ _21930_/Y _21931_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _21932_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24651_ hold1945/X _26280_/Q _24664_/S vssd1 vssd1 vccd1 vccd1 _24651_/X sky130_fd_sc_hd__mux2_1
X_21863_ _21861_/Y _21862_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21863_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_171_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23602_ _23602_/A vssd1 vssd1 vccd1 vccd1 _23920_/S sky130_fd_sc_hd__buf_4
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20814_ _20814_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _20814_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21794_ _21792_/Y _21793_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21794_/Y sky130_fd_sc_hd__a21oi_1
X_24582_ _24582_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24583_/A sky130_fd_sc_hd__and2_1
XFILLER_0_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26321_ _26325_/CLK _26321_/D vssd1 vssd1 vccd1 vccd1 _26321_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_65_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23533_ hold158/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23533_/X sky130_fd_sc_hd__or2b_1
X_20745_ _20745_/A _21734_/B _20745_/C vssd1 vssd1 vccd1 vccd1 _20748_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26252_ _26252_/CLK _26252_/D vssd1 vssd1 vccd1 vccd1 _26252_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_135_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20676_ _23085_/B vssd1 vssd1 vccd1 vccd1 _22544_/B sky130_fd_sc_hd__inv_2
X_23464_ hold53/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23464_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25203_ _25783_/CLK hold538/X vssd1 vssd1 vccd1 vccd1 hold536/A sky130_fd_sc_hd__dfxtp_1
X_22415_ _22992_/B vssd1 vssd1 vccd1 vccd1 _22991_/B sky130_fd_sc_hd__inv_2
XFILLER_0_18_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26183_ _26184_/CLK _26183_/D vssd1 vssd1 vccd1 vccd1 _26183_/Q sky130_fd_sc_hd__dfxtp_1
X_23395_ _23388_/X _23394_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _23395_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_162_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25134_ _26122_/CLK hold767/X vssd1 vssd1 vccd1 vccd1 hold766/A sky130_fd_sc_hd__dfxtp_1
X_22346_ _22346_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _22346_/X sky130_fd_sc_hd__and2_1
XFILLER_0_27_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22277_ _22277_/A _25855_/Q vssd1 vssd1 vccd1 vccd1 _22277_/Y sky130_fd_sc_hd__nand2_1
X_25065_ _26151_/CLK _25065_/D vssd1 vssd1 vccd1 vccd1 _25065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24016_ _24016_/A vssd1 vssd1 vccd1 vccd1 _26073_/D sky130_fd_sc_hd__clkbuf_1
X_21228_ _21228_/A vssd1 vssd1 vccd1 vccd1 _21228_/X sky130_fd_sc_hd__buf_4
Xhold170 hold170/A vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold181 hold181/A vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 hold192/A vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
X_21159_ _21159_/A _25871_/Q vssd1 vssd1 vccd1 vccd1 _21164_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25967_ _26042_/CLK _25967_/D vssd1 vssd1 vccd1 vccd1 _25967_/Q sky130_fd_sc_hd__dfxtp_1
X_13981_ _14170_/A vssd1 vssd1 vccd1 vccd1 _13981_/X sky130_fd_sc_hd__clkbuf_16
X_15720_ _15701_/A _15763_/A _15719_/X vssd1 vssd1 vccd1 vccd1 _15720_/X sky130_fd_sc_hd__a21bo_1
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24918_ _24946_/A _24915_/X _24958_/B _24917_/Y vssd1 vssd1 vccd1 vccd1 _24918_/X
+ sky130_fd_sc_hd__a211o_1
X_12932_ _12891_/X _14397_/A _12909_/X _25617_/Q vssd1 vssd1 vccd1 vccd1 _12932_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25898_ _25898_/CLK _25898_/D vssd1 vssd1 vccd1 vccd1 _25898_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15651_ _23044_/B _15776_/B vssd1 vssd1 vccd1 vccd1 _16571_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_73_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24849_ _15341_/A _15356_/B _24863_/S vssd1 vssd1 vccd1 vccd1 _24849_/X sky130_fd_sc_hd__mux2_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _26107_/Q _12748_/X _12862_/X vssd1 vssd1 vccd1 vccd1 _12863_/X sky130_fd_sc_hd__a21o_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14602_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14602_/Y sky130_fd_sc_hd__nand2_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18370_ _18370_/A _21183_/A vssd1 vssd1 vccd1 vccd1 _18718_/A sky130_fd_sc_hd__xor2_4
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15582_ _15582_/A _15810_/B vssd1 vssd1 vccd1 vccd1 _15583_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_29_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12726_/B _14316_/A _12752_/X _25591_/Q vssd1 vssd1 vccd1 vccd1 _12794_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _17520_/A _17321_/B vssd1 vssd1 vccd1 vccd1 _17321_/X sky130_fd_sc_hd__xor2_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14533_ _14533_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14533_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_55_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17252_ _20752_/B _25896_/Q _25832_/Q vssd1 vssd1 vccd1 vccd1 _17253_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_55_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14464_ _14464_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14464_/Y sky130_fd_sc_hd__nand2_1
X_16203_ _16676_/A _16203_/B vssd1 vssd1 vccd1 vccd1 _16205_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13415_ _13220_/A _14663_/A _13242_/X _19816_/A vssd1 vssd1 vccd1 vccd1 _13415_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17183_ _20558_/B _25891_/Q _25827_/Q vssd1 vssd1 vccd1 vccd1 _17184_/B sky130_fd_sc_hd__mux2_2
X_14395_ _14404_/A hold353/X vssd1 vssd1 vccd1 vccd1 hold354/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16134_ _16134_/A _16134_/B vssd1 vssd1 vccd1 vccd1 _16157_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_144_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13346_ _13315_/X _13344_/X _13300_/X _13345_/X vssd1 vssd1 vccd1 vccd1 _13346_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16065_ _16063_/Y hold801/X _15805_/X vssd1 vssd1 vccd1 vccd1 hold802/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13277_ _13277_/A vssd1 vssd1 vccd1 vccd1 _19504_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15016_ _14997_/B _15015_/A _15007_/B vssd1 vssd1 vccd1 vccd1 _15016_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_166_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19824_ _19975_/A _19824_/B vssd1 vssd1 vccd1 vccd1 _19824_/Y sky130_fd_sc_hd__nand2_1
Xhold1809 _22364_/Y vssd1 vssd1 vccd1 vccd1 _25858_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19755_ _26258_/Q hold524/X vssd1 vssd1 vccd1 vccd1 _19755_/Y sky130_fd_sc_hd__nand2_1
X_16967_ _16967_/A _16967_/B vssd1 vssd1 vccd1 vccd1 _16967_/Y sky130_fd_sc_hd__nand2_1
X_18706_ _20479_/B _19758_/A vssd1 vssd1 vccd1 vccd1 _18707_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15918_ _15918_/A _15918_/B vssd1 vssd1 vccd1 vccd1 _15919_/B sky130_fd_sc_hd__nand2_1
X_16898_ _16896_/X _16711_/X _16897_/Y _25889_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16899_/A sky130_fd_sc_hd__a32o_1
X_19686_ _19683_/Y _19686_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19686_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15849_ _15846_/B _15869_/B _15848_/Y vssd1 vssd1 vccd1 vccd1 _15849_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_149_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18637_ _18637_/A _18637_/B vssd1 vssd1 vccd1 vccd1 _18637_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_176_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18568_ _18793_/A _25754_/Q _18894_/C vssd1 vssd1 vccd1 vccd1 _18569_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_176_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17519_ _17519_/A _17570_/A vssd1 vssd1 vccd1 vccd1 _17520_/B sky130_fd_sc_hd__xnor2_1
X_18499_ _18497_/Y _18498_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25669_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20530_ _21578_/A _21305_/B vssd1 vssd1 vccd1 vccd1 _20531_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_156_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20461_ _21042_/A _20461_/B _20460_/X vssd1 vssd1 vccd1 vccd1 _20462_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_55_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22200_ _22177_/X _22199_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _22200_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23180_ _23171_/Y _23179_/Y _19199_/A vssd1 vssd1 vccd1 vccd1 _23180_/X sky130_fd_sc_hd__a21o_1
X_20392_ _20392_/A _25848_/Q vssd1 vssd1 vccd1 vccd1 _20397_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22131_ _25786_/Q _22131_/B vssd1 vssd1 vccd1 vccd1 _22131_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22062_ _22060_/X _15839_/B _22061_/Y _14795_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _22063_/A sky130_fd_sc_hd__a32o_1
X_21013_ _26304_/Q _20731_/X hold371/X vssd1 vssd1 vccd1 vccd1 _21016_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25821_ _25822_/CLK _25821_/D vssd1 vssd1 vccd1 vccd1 _25821_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25752_ _25752_/CLK _25752_/D vssd1 vssd1 vccd1 vccd1 _25752_/Q sky130_fd_sc_hd__dfxtp_1
X_22964_ _26070_/Q vssd1 vssd1 vccd1 vccd1 _22965_/A sky130_fd_sc_hd__inv_2
XFILLER_0_168_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24703_ _24703_/A vssd1 vssd1 vccd1 vccd1 _26296_/D sky130_fd_sc_hd__clkbuf_1
X_21915_ _21915_/A _21915_/B vssd1 vssd1 vccd1 vccd1 _21915_/Y sky130_fd_sc_hd__nand2_1
X_25683_ _25687_/CLK _25683_/D vssd1 vssd1 vccd1 vccd1 _25683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22895_ _26066_/Q vssd1 vssd1 vccd1 vccd1 _22896_/A sky130_fd_sc_hd__inv_2
XFILLER_0_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24634_ _24634_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24635_/A sky130_fd_sc_hd__and2_1
XFILLER_0_167_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21846_ _21846_/A _21846_/B vssd1 vssd1 vccd1 vccd1 _21846_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24565_ _24565_/A vssd1 vssd1 vccd1 vccd1 _26251_/D sky130_fd_sc_hd__clkbuf_1
X_21777_ _25867_/Q _21778_/A vssd1 vssd1 vccd1 vccd1 _21779_/A sky130_fd_sc_hd__or2_1
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26304_ _26306_/CLK _26304_/D vssd1 vssd1 vccd1 vccd1 _26304_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23516_ hold161/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23516_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_135_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20728_ _20728_/A _21338_/B _20728_/C vssd1 vssd1 vccd1 vccd1 _20729_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24496_ _24496_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24497_/A sky130_fd_sc_hd__and2_1
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26235_ _26235_/CLK _26235_/D vssd1 vssd1 vccd1 vccd1 _26235_/Q sky130_fd_sc_hd__dfxtp_2
X_23447_ _24922_/S hold137/A _23446_/X vssd1 vssd1 vccd1 vccd1 _23447_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20659_ _20659_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _20659_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_18_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ _13109_/X _13198_/X _13192_/X _13199_/X vssd1 vssd1 vccd1 vccd1 _13200_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14180_ _14180_/A _14180_/B vssd1 vssd1 vccd1 vccd1 _14180_/Y sky130_fd_sc_hd__nand2_1
X_26166_ _26297_/CLK _26166_/D vssd1 vssd1 vccd1 vccd1 _26166_/Q sky130_fd_sc_hd__dfxtp_1
X_23378_ _23378_/A vssd1 vssd1 vccd1 vccd1 _25938_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25117_ _26198_/CLK _25117_/D vssd1 vssd1 vccd1 vccd1 _25117_/Q sky130_fd_sc_hd__dfxtp_1
X_13131_ _13049_/X _14518_/A _13067_/X _25655_/Q vssd1 vssd1 vccd1 vccd1 _13131_/X
+ sky130_fd_sc_hd__a22o_1
X_22329_ _22329_/A _22329_/B vssd1 vssd1 vccd1 vccd1 _22329_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26097_ _26103_/CLK _26097_/D vssd1 vssd1 vccd1 vccd1 _26097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25048_ _26130_/CLK _25048_/D vssd1 vssd1 vccd1 vccd1 _25048_/Q sky130_fd_sc_hd__dfxtp_1
X_13062_ _26145_/Q _12907_/X _13061_/X vssd1 vssd1 vccd1 vccd1 _13062_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17870_ _25648_/Q vssd1 vssd1 vccd1 vccd1 _21821_/A sky130_fd_sc_hd__inv_2
XFILLER_0_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16821_ _16819_/Y _16820_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16821_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16752_ _16980_/A _16757_/B vssd1 vssd1 vccd1 vccd1 _16754_/B sky130_fd_sc_hd__nand2_1
X_19540_ _19723_/A _19540_/B vssd1 vssd1 vccd1 vccd1 _19540_/Y sky130_fd_sc_hd__nand2_1
X_13964_ _18035_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13964_/Y sky130_fd_sc_hd__nor2_1
X_15703_ _15703_/A vssd1 vssd1 vccd1 vccd1 _15712_/B sky130_fd_sc_hd__inv_2
X_12915_ _12891_/X _14388_/A _12909_/X _25614_/Q vssd1 vssd1 vccd1 vccd1 _12915_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16683_ _16683_/A _16683_/B vssd1 vssd1 vccd1 vccd1 _16685_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_159_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19471_ _19470_/Y _19272_/X _19131_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19472_/B
+ sky130_fd_sc_hd__a211o_1
X_13895_ _20197_/B vssd1 vssd1 vccd1 vccd1 _17976_/B sky130_fd_sc_hd__inv_2
XFILLER_0_115_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15634_ _15634_/A _15810_/B vssd1 vssd1 vccd1 vccd1 _15635_/B sky130_fd_sc_hd__nand2_1
X_18422_ _21265_/B _19560_/A vssd1 vssd1 vccd1 vccd1 _18423_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_158_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12846_ _26232_/Q _25601_/Q vssd1 vssd1 vccd1 vccd1 _14348_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18353_ _18535_/A hold979/X _18393_/C vssd1 vssd1 vccd1 vccd1 _18353_/X sky130_fd_sc_hd__and3_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15565_ _15565_/A _15810_/B vssd1 vssd1 vccd1 vccd1 _15566_/B sky130_fd_sc_hd__nand2_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12777_ _12746_/X hold993/X _14910_/B _12776_/X vssd1 vssd1 vccd1 vccd1 hold994/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _25644_/Q vssd1 vssd1 vccd1 vccd1 _20044_/B sky130_fd_sc_hd__inv_2
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14516_ _14525_/A hold179/X vssd1 vssd1 vccd1 vccd1 hold180/A sky130_fd_sc_hd__nand2_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18284_ _18528_/A vssd1 vssd1 vccd1 vccd1 _18951_/A sky130_fd_sc_hd__buf_12
X_15496_ _15496_/A _15496_/B vssd1 vssd1 vccd1 vccd1 _15502_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17235_ _25639_/Q vssd1 vssd1 vccd1 vccd1 _20712_/B sky130_fd_sc_hd__inv_2
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14447_ _14465_/A hold272/X vssd1 vssd1 vccd1 vccd1 hold273/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17166_ _25600_/Q vssd1 vssd1 vccd1 vccd1 _20702_/B sky130_fd_sc_hd__inv_2
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14378_ _14376_/Y hold243/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold244/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold906 hold906/A vssd1 vssd1 vccd1 vccd1 hold906/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16117_ _16133_/A _16133_/B _16134_/A _16116_/Y vssd1 vssd1 vccd1 vccd1 _16117_/X
+ sky130_fd_sc_hd__a31o_1
Xhold917 hold917/A vssd1 vssd1 vccd1 vccd1 hold917/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold928 hold928/A vssd1 vssd1 vccd1 vccd1 hold928/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13329_ _13329_/A vssd1 vssd1 vccd1 vccd1 _19616_/A sky130_fd_sc_hd__clkbuf_8
X_17097_ _17095_/Y _17096_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _17097_/Y sky130_fd_sc_hd__a21oi_1
Xhold939 hold939/A vssd1 vssd1 vccd1 vccd1 hold939/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16048_ _16049_/B _16049_/A vssd1 vssd1 vccd1 vccd1 _16071_/B sky130_fd_sc_hd__or2_1
XFILLER_0_161_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2307 _26118_/Q vssd1 vssd1 vccd1 vccd1 hold2307/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2318 _26140_/Q vssd1 vssd1 vccd1 vccd1 hold2318/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2329 _26262_/Q vssd1 vssd1 vccd1 vccd1 hold2329/X sky130_fd_sc_hd__dlygate4sd3_1
X_19807_ _19807_/A _19807_/B vssd1 vssd1 vccd1 vccd1 _19807_/Y sky130_fd_sc_hd__nand2_1
Xhold1606 _25811_/Q vssd1 vssd1 vccd1 vccd1 _21288_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1617 _17287_/Y vssd1 vssd1 vccd1 vccd1 _25601_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1628 _25834_/Q vssd1 vssd1 vccd1 vccd1 _21671_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17999_ _18612_/A _19424_/B _18083_/C vssd1 vssd1 vccd1 vccd1 _18000_/C sky130_fd_sc_hd__nand3_1
Xhold1639 _25617_/Q vssd1 vssd1 vccd1 vccd1 _17453_/B sky130_fd_sc_hd__dlygate4sd3_1
X_19738_ _19975_/A _19738_/B vssd1 vssd1 vccd1 vccd1 _19738_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_159_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19669_ _26252_/Q _19483_/X hold542/X vssd1 vssd1 vccd1 vccd1 _19669_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21700_ _21716_/A _21700_/B _21699_/X vssd1 vssd1 vccd1 vccd1 _21701_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_35_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22680_ _22680_/A vssd1 vssd1 vccd1 vccd1 _22680_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_176_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21631_ _21631_/A _21631_/B vssd1 vssd1 vccd1 vccd1 _21632_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24350_ hold2016/X _26182_/Q _24356_/S vssd1 vssd1 vccd1 vccd1 _24350_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21562_ _21562_/A _21611_/A vssd1 vssd1 vccd1 vccd1 _21564_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23301_ _23301_/A hold985/X vssd1 vssd1 vccd1 vccd1 hold986/A sky130_fd_sc_hd__nand2_1
X_20513_ _20513_/A _20513_/B vssd1 vssd1 vccd1 vccd1 _20515_/A sky130_fd_sc_hd__nand2_1
X_21493_ _23245_/A vssd1 vssd1 vccd1 vccd1 _21493_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24281_ _24281_/A vssd1 vssd1 vccd1 vccd1 _26159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26020_ _26032_/CLK _26020_/D vssd1 vssd1 vccd1 vccd1 _26020_/Q sky130_fd_sc_hd__dfxtp_1
X_23232_ _23232_/A vssd1 vssd1 vccd1 vccd1 _24958_/B sky130_fd_sc_hd__buf_12
X_20444_ _20447_/A _20447_/C vssd1 vssd1 vccd1 vccd1 _20446_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23163_ _23163_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _23163_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20375_ _20375_/A _20375_/B _21114_/C vssd1 vssd1 vccd1 vccd1 _20379_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_113_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22114_ _22112_/Y _22113_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _22114_/Y sky130_fd_sc_hd__a21oi_1
X_23094_ _26078_/Q vssd1 vssd1 vccd1 vccd1 _23095_/A sky130_fd_sc_hd__inv_2
XFILLER_0_100_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22045_ _22045_/A _22772_/B vssd1 vssd1 vccd1 vccd1 _22046_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25804_ _25808_/CLK _25804_/D vssd1 vssd1 vccd1 vccd1 _25804_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_98_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23996_ _23996_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23997_/A sky130_fd_sc_hd__and2_1
XFILLER_0_138_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25735_ _25740_/CLK _25735_/D vssd1 vssd1 vccd1 vccd1 _25735_/Q sky130_fd_sc_hd__dfxtp_1
X_22947_ _26069_/Q vssd1 vssd1 vccd1 vccd1 _22948_/A sky130_fd_sc_hd__inv_2
XFILLER_0_168_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12700_ _12713_/B _12700_/B vssd1 vssd1 vccd1 vccd1 _12701_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_70_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25666_ _26297_/CLK _25666_/D vssd1 vssd1 vccd1 vccd1 _25666_/Q sky130_fd_sc_hd__dfxtp_1
X_13680_ hold546/X _13678_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold547/A sky130_fd_sc_hd__a21oi_1
X_22878_ _22878_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22878_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12631_ _12631_/A vssd1 vssd1 vccd1 vccd1 _24979_/D sky130_fd_sc_hd__clkbuf_1
X_24617_ _24617_/A vssd1 vssd1 vccd1 vccd1 _26268_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21829_ _21827_/Y _21828_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21829_/Y sky130_fd_sc_hd__a21oi_1
X_25597_ _26109_/CLK _25597_/D vssd1 vssd1 vccd1 vccd1 _25597_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_66_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15350_ _15350_/A _15776_/B vssd1 vssd1 vccd1 vccd1 _15351_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_164_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12562_ _12562_/A vssd1 vssd1 vccd1 vccd1 _23597_/C sky130_fd_sc_hd__inv_4
X_24548_ _24548_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24549_/A sky130_fd_sc_hd__and2_1
XFILLER_0_109_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14301_ _14301_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14301_/Y sky130_fd_sc_hd__nand2_1
X_15281_ _25445_/Q vssd1 vssd1 vccd1 vccd1 _15290_/B sky130_fd_sc_hd__inv_2
X_12493_ _24999_/Q vssd1 vssd1 vccd1 vccd1 _13220_/A sky130_fd_sc_hd__clkbuf_16
X_24479_ _24479_/A vssd1 vssd1 vccd1 vccd1 _26223_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17020_ _17867_/B _17020_/B vssd1 vssd1 vccd1 vccd1 _17616_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_149_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26218_ _26219_/CLK _26218_/D vssd1 vssd1 vccd1 vccd1 _26218_/Q sky130_fd_sc_hd__dfxtp_2
X_14232_ _18854_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14232_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_22_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26149_ _26151_/CLK _26149_/D vssd1 vssd1 vccd1 vccd1 _26149_/Q sky130_fd_sc_hd__dfxtp_1
X_14163_ _14236_/A hold839/X vssd1 vssd1 vccd1 vccd1 _14163_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_145_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13114_ _13109_/X _13112_/X _13096_/X _13113_/X vssd1 vssd1 vccd1 vccd1 _13114_/X
+ sky130_fd_sc_hd__o211a_1
X_14094_ _14118_/A hold539/X vssd1 vssd1 vccd1 vccd1 hold540/A sky130_fd_sc_hd__nand2_1
X_18971_ _18971_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _18971_/Y sky130_fd_sc_hd__nand2_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_2__f_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_2__f_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _25841_/Q vssd1 vssd1 vccd1 vccd1 _20144_/A sky130_fd_sc_hd__inv_2
X_13045_ _12891_/X _14469_/A _12909_/X _25639_/Q vssd1 vssd1 vccd1 vccd1 _13045_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17853_ _25849_/Q _17853_/B _17853_/C vssd1 vssd1 vccd1 vccd1 _17861_/A sky130_fd_sc_hd__or3_2
XFILLER_0_79_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16804_ _16802_/X _16711_/X _16803_/Y _25875_/Q _14170_/X vssd1 vssd1 vccd1 vccd1
+ _16805_/A sky130_fd_sc_hd__a32o_1
X_14996_ _14996_/A _14996_/B vssd1 vssd1 vccd1 vccd1 _14997_/B sky130_fd_sc_hd__nand2_1
X_17784_ _17784_/A _17784_/B vssd1 vssd1 vccd1 vccd1 _18119_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_89_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19523_ _19523_/A _19523_/B vssd1 vssd1 vccd1 vccd1 _19523_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_163_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16735_ _16735_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16735_/Y sky130_fd_sc_hd__nand2_1
X_13947_ _26289_/Q _13801_/X _13793_/X _13946_/Y vssd1 vssd1 vccd1 vccd1 _13948_/B
+ sky130_fd_sc_hd__a22o_1
X_16666_ _16667_/B _16667_/A vssd1 vssd1 vccd1 vccd1 _16668_/A sky130_fd_sc_hd__or2_1
X_19454_ _26237_/Q _12537_/B hold491/X vssd1 vssd1 vccd1 vccd1 _19454_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13878_ _13941_/A _13878_/B vssd1 vssd1 vccd1 vccd1 _13878_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_9_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15617_ _26033_/Q _25969_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15618_/A sky130_fd_sc_hd__mux2_1
X_18405_ _18405_/A _25810_/Q _18405_/C vssd1 vssd1 vccd1 vccd1 _21243_/B sky130_fd_sc_hd__nand3_1
X_12829_ _12746_/X _12826_/X _12827_/X _12828_/X vssd1 vssd1 vccd1 vccd1 _12829_/X
+ sky130_fd_sc_hd__o211a_1
X_16597_ _16597_/A _16597_/B vssd1 vssd1 vccd1 vccd1 _16598_/A sky130_fd_sc_hd__nand2_1
X_19385_ _26232_/Q hold590/X vssd1 vssd1 vccd1 vccd1 _19385_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15548_ _15548_/A _15548_/B vssd1 vssd1 vccd1 vccd1 _15549_/A sky130_fd_sc_hd__nor2_1
X_18336_ _18641_/A _19244_/A vssd1 vssd1 vccd1 vccd1 _18336_/Y sky130_fd_sc_hd__nand2_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18267_ _18474_/A _18617_/A vssd1 vssd1 vccd1 vccd1 _18268_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15479_ _15479_/A vssd1 vssd1 vccd1 vccd1 _16848_/A sky130_fd_sc_hd__inv_2
XFILLER_0_112_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_150_clk clkbuf_4_11__f_clk/X vssd1 vssd1 vccd1 vccd1 _26181_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17218_ _17216_/Y _17217_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _17218_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18198_ _18445_/A _18202_/B vssd1 vssd1 vccd1 vccd1 _18200_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_170_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold703 hold703/A vssd1 vssd1 vccd1 vccd1 hold703/X sky130_fd_sc_hd__dlygate4sd3_1
X_17149_ _17147_/X _23187_/B _17148_/X vssd1 vssd1 vccd1 vccd1 _17150_/A sky130_fd_sc_hd__a21o_1
Xhold714 hold714/A vssd1 vssd1 vccd1 vccd1 hold714/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold725 hold725/A vssd1 vssd1 vccd1 vccd1 hold725/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 hold736/A vssd1 vssd1 vccd1 vccd1 hold736/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold747 hold747/A vssd1 vssd1 vccd1 vccd1 hold747/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20160_ _20660_/A _20160_/B vssd1 vssd1 vccd1 vccd1 _20160_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold758 hold758/A vssd1 vssd1 vccd1 vccd1 hold758/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold769 hold769/A vssd1 vssd1 vccd1 vccd1 hold769/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20091_ _20091_/A _22723_/B vssd1 vssd1 vccd1 vccd1 _20095_/B sky130_fd_sc_hd__nand2_1
Xhold2104 _24725_/X vssd1 vssd1 vccd1 vccd1 _24726_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2115 _25433_/Q vssd1 vssd1 vccd1 vccd1 _15076_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2126 _26046_/Q vssd1 vssd1 vccd1 vccd1 hold2126/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2137 _25918_/Q vssd1 vssd1 vccd1 vccd1 _23278_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold2148 _15089_/Y vssd1 vssd1 vccd1 vccd1 hold2148/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1403 _25403_/Q vssd1 vssd1 vccd1 vccd1 _14831_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1414 _23070_/Y vssd1 vssd1 vccd1 vccd1 _25893_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2159 _26128_/Q vssd1 vssd1 vccd1 vccd1 hold2159/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1425 _25722_/Q vssd1 vssd1 vccd1 vccd1 _19297_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1436 _13352_/X vssd1 vssd1 vccd1 vccd1 _25110_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23850_ hold1928/X _26021_/Q _23907_/S vssd1 vssd1 vccd1 vccd1 _23850_/X sky130_fd_sc_hd__mux2_1
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1447 _25739_/Q vssd1 vssd1 vccd1 vccd1 _19540_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1458 _20198_/Y vssd1 vssd1 vccd1 vccd1 _25778_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1469 _25837_/Q vssd1 vssd1 vccd1 vccd1 _21719_/B sky130_fd_sc_hd__dlygate4sd3_1
X_22801_ _22801_/A _23001_/B _22801_/C vssd1 vssd1 vccd1 vccd1 _22801_/X sky130_fd_sc_hd__and3_1
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23781_ _23781_/A vssd1 vssd1 vccd1 vccd1 _25998_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20993_ _20993_/A _22006_/B vssd1 vssd1 vccd1 vccd1 _20994_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_170_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25520_ _25534_/CLK hold867/X vssd1 vssd1 vccd1 vccd1 hold866/A sky130_fd_sc_hd__dfxtp_1
X_22732_ _15317_/B _22680_/X _14273_/X vssd1 vssd1 vccd1 vccd1 _22732_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25451_ _26057_/CLK _25451_/D vssd1 vssd1 vccd1 vccd1 _25451_/Q sky130_fd_sc_hd__dfxtp_1
X_22663_ _22661_/X _22662_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22663_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24402_ _24402_/A vssd1 vssd1 vccd1 vccd1 _26198_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21614_ _21614_/A _21614_/B vssd1 vssd1 vccd1 vccd1 _21616_/A sky130_fd_sc_hd__nand2_1
X_25382_ _26205_/CLK hold64/X vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22594_ _22595_/B _22595_/A vssd1 vssd1 vccd1 vccd1 _22596_/A sky130_fd_sc_hd__or2_1
XFILLER_0_30_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24333_ _24333_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24334_/A sky130_fd_sc_hd__and2_1
XFILLER_0_62_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21545_ _21545_/A _21545_/B _21545_/C vssd1 vssd1 vccd1 vccd1 _21549_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_168_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_141_clk clkbuf_4_11__f_clk/X vssd1 vssd1 vccd1 vccd1 _25807_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24264_ hold2235/X hold2221/X _24279_/S vssd1 vssd1 vccd1 vccd1 _24265_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_161_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21476_ _21573_/A _21476_/B vssd1 vssd1 vccd1 vccd1 _21476_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26003_ _26047_/CLK _26003_/D vssd1 vssd1 vccd1 vccd1 _26003_/Q sky130_fd_sc_hd__dfxtp_1
X_23215_ _23215_/A vssd1 vssd1 vccd1 vccd1 _24863_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_160_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20427_ _20425_/Y _20426_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _20427_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24195_ _24195_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24196_/A sky130_fd_sc_hd__and2_1
X_23146_ _16963_/B _22421_/A _23140_/X _23141_/Y _23145_/X vssd1 vssd1 vccd1 vccd1
+ _23147_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_140_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20358_ _20358_/A _20358_/B _20358_/C vssd1 vssd1 vccd1 vccd1 _20359_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23077_ _15684_/B _22893_/A _22829_/X vssd1 vssd1 vccd1 vccd1 _23077_/Y sky130_fd_sc_hd__a21oi_1
X_20289_ _20291_/B _20291_/C vssd1 vssd1 vccd1 vccd1 _20290_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_140_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22028_ _22028_/A _22028_/B vssd1 vssd1 vccd1 vccd1 _23026_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_175_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2660 _26238_/Q vssd1 vssd1 vccd1 vccd1 hold2660/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2671 _25457_/Q vssd1 vssd1 vccd1 vccd1 _15486_/A sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ _14900_/A _14852_/A vssd1 vssd1 vccd1 vccd1 _14850_/Y sky130_fd_sc_hd__nand2_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2682 _15821_/Y vssd1 vssd1 vccd1 vccd1 _25475_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2693 _26331_/Q vssd1 vssd1 vccd1 vccd1 hold2693/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ _14262_/B vssd1 vssd1 vccd1 vccd1 _13801_/X sky130_fd_sc_hd__buf_12
XFILLER_0_98_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1970 _12582_/Y vssd1 vssd1 vccd1 vccd1 _12583_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold1981 _26341_/Q vssd1 vssd1 vccd1 vccd1 hold1981/X sky130_fd_sc_hd__dlygate4sd3_1
X_14781_ _22035_/B _15778_/B vssd1 vssd1 vccd1 vccd1 _14782_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1992 _23622_/X vssd1 vssd1 vccd1 vccd1 _23623_/A sky130_fd_sc_hd__dlygate4sd3_1
X_23979_ _23979_/A vssd1 vssd1 vccd1 vccd1 _26061_/D sky130_fd_sc_hd__clkbuf_1
X_16520_ _16676_/A _16520_/B vssd1 vssd1 vccd1 vccd1 _16522_/A sky130_fd_sc_hd__or2_1
XFILLER_0_168_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25718_ _26244_/CLK hold924/X vssd1 vssd1 vccd1 vccd1 hold922/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_10__f_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_10__f_clk/X
+ sky130_fd_sc_hd__clkbuf_16
X_13732_ _18529_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13732_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_98_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16451_ _16451_/A hold935/X _16691_/B vssd1 vssd1 vccd1 vccd1 _16452_/B sky130_fd_sc_hd__and3_1
XFILLER_0_183_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25649_ _26152_/CLK _25649_/D vssd1 vssd1 vccd1 vccd1 _25649_/Q sky130_fd_sc_hd__dfxtp_1
X_13663_ hold981/A vssd1 vssd1 vccd1 vccd1 _18307_/B sky130_fd_sc_hd__inv_2
XFILLER_0_38_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15402_ _15403_/B _16824_/A vssd1 vssd1 vccd1 vccd1 _15404_/A sky130_fd_sc_hd__nor2_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12614_ _12614_/A _24836_/B _12618_/A vssd1 vssd1 vccd1 vccd1 _12614_/X sky130_fd_sc_hd__and3_1
X_19170_ _19186_/A hold815/X vssd1 vssd1 vccd1 vccd1 hold816/A sky130_fd_sc_hd__nand2_1
X_16382_ _16490_/A _16382_/B vssd1 vssd1 vccd1 vccd1 _16393_/A sky130_fd_sc_hd__nand2_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13594_ _17957_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13594_/Y sky130_fd_sc_hd__nor2_1
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18121_ _18121_/A hold937/A vssd1 vssd1 vccd1 vccd1 _18125_/A sky130_fd_sc_hd__nand2_2
X_15333_ _26017_/Q _25953_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15334_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12545_ _14267_/A vssd1 vssd1 vccd1 vccd1 _20957_/A sky130_fd_sc_hd__inv_8
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_132_clk clkbuf_leaf_82_clk/A vssd1 vssd1 vccd1 vccd1 _26340_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_124_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18052_ _18793_/A _18052_/B _18891_/C vssd1 vssd1 vccd1 vccd1 _18053_/C sky130_fd_sc_hd__nand3_1
X_15264_ _15264_/A _15264_/B vssd1 vssd1 vccd1 vccd1 _15265_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17003_ _19082_/A vssd1 vssd1 vccd1 vccd1 _17393_/A sky130_fd_sc_hd__buf_6
X_14215_ _26332_/Q _13518_/B _14170_/X _14214_/Y vssd1 vssd1 vccd1 vccd1 _14216_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA_5 _22228_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ hold927/X _15197_/A vssd1 vssd1 vccd1 vccd1 _15199_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_105_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14146_ _18572_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14146_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18954_ _18954_/A _25773_/Q vssd1 vssd1 vccd1 vccd1 _18956_/A sky130_fd_sc_hd__nand2_1
X_14077_ _25807_/Q vssd1 vssd1 vccd1 vccd1 _18348_/B sky130_fd_sc_hd__inv_2
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17905_ _18612_/A _25729_/Q _18083_/C vssd1 vssd1 vccd1 vccd1 _17906_/C sky130_fd_sc_hd__nand3_1
X_13028_ _13018_/X _13026_/X _13005_/X _13027_/X vssd1 vssd1 vccd1 vccd1 _13028_/X
+ sky130_fd_sc_hd__o211a_1
X_18885_ _25706_/Q _20829_/B vssd1 vssd1 vccd1 vccd1 _18888_/A sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_199_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _25604_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_174_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17836_ _17836_/A _19093_/A vssd1 vssd1 vccd1 vccd1 _19025_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_89_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17767_ _17766_/B _17767_/B vssd1 vssd1 vccd1 vccd1 _17781_/C sky130_fd_sc_hd__nand2b_1
X_14979_ _14980_/B _14980_/A vssd1 vssd1 vccd1 vccd1 _14981_/A sky130_fd_sc_hd__or2_1
XFILLER_0_117_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19506_ _21156_/A _19504_/Y _21160_/C vssd1 vssd1 vccd1 vccd1 _19593_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_159_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16718_ _16719_/B _16719_/A vssd1 vssd1 vccd1 vccd1 _16718_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17698_ _17698_/A _17725_/B vssd1 vssd1 vccd1 vccd1 _17705_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_159_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19437_ _19429_/X _19436_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19437_/Y sky130_fd_sc_hd__o21ai_1
X_16649_ _16649_/A _16649_/B vssd1 vssd1 vccd1 vccd1 _16650_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19368_ _19366_/Y _19367_/Y _19086_/X vssd1 vssd1 vccd1 vccd1 _19368_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18319_ _21878_/B _25614_/Q vssd1 vssd1 vccd1 vccd1 _18321_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_123_clk clkbuf_4_11__f_clk/X vssd1 vssd1 vccd1 vccd1 _26325_/CLK sky130_fd_sc_hd__clkbuf_16
X_19299_ _26226_/Q _12537_/B hold581/X vssd1 vssd1 vccd1 vccd1 _19299_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21330_ _21330_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21330_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_143_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21261_ _22586_/A vssd1 vssd1 vccd1 vccd1 _21573_/A sky130_fd_sc_hd__clkbuf_8
Xhold500 hold500/A vssd1 vssd1 vccd1 vccd1 hold500/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 hold511/A vssd1 vssd1 vccd1 vccd1 hold511/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold522 hold522/A vssd1 vssd1 vccd1 vccd1 hold522/X sky130_fd_sc_hd__dlygate4sd3_1
X_23000_ _22999_/A _22849_/X _22999_/B vssd1 vssd1 vccd1 vccd1 _23001_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold533 hold533/A vssd1 vssd1 vccd1 vccd1 hold533/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20212_ _20214_/A _20214_/C vssd1 vssd1 vccd1 vccd1 _20213_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21192_ _21643_/C vssd1 vssd1 vccd1 vccd1 _21646_/B sky130_fd_sc_hd__inv_2
Xhold544 hold544/A vssd1 vssd1 vccd1 vccd1 hold544/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 hold555/A vssd1 vssd1 vccd1 vccd1 hold555/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 hold566/A vssd1 vssd1 vccd1 vccd1 hold566/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold577 hold577/A vssd1 vssd1 vccd1 vccd1 hold577/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20143_ _20143_/A _20143_/B vssd1 vssd1 vccd1 vccd1 _20144_/B sky130_fd_sc_hd__nand2_1
Xhold588 hold588/A vssd1 vssd1 vccd1 vccd1 hold588/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold599 hold599/A vssd1 vssd1 vccd1 vccd1 hold599/X sky130_fd_sc_hd__dlygate4sd3_1
X_24951_ hold948/X hold920/X _24956_/S vssd1 vssd1 vccd1 vccd1 _24951_/X sky130_fd_sc_hd__mux2_1
X_20074_ _21693_/A _21386_/A vssd1 vssd1 vccd1 vccd1 _20075_/C sky130_fd_sc_hd__nand2_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1200 _19597_/Y vssd1 vssd1 vccd1 vccd1 _25743_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1211 _25750_/Q vssd1 vssd1 vccd1 vccd1 _19695_/B sky130_fd_sc_hd__dlygate4sd3_1
X_23902_ _23902_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23903_/A sky130_fd_sc_hd__and2_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1222 _19710_/Y vssd1 vssd1 vccd1 vccd1 _25751_/D sky130_fd_sc_hd__dlygate4sd3_1
X_24882_ hold964/A hold861/A _24956_/S vssd1 vssd1 vccd1 vccd1 _24883_/B sky130_fd_sc_hd__mux2_1
Xhold1233 _16934_/Y vssd1 vssd1 vccd1 vccd1 _25573_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1244 _25710_/Q vssd1 vssd1 vccd1 vccd1 _19112_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1255 _16765_/Y vssd1 vssd1 vccd1 vccd1 _25548_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1266 _25790_/Q vssd1 vssd1 vccd1 vccd1 _20660_/B sky130_fd_sc_hd__clkdlybuf4s25_1
X_23833_ _23833_/A vssd1 vssd1 vccd1 vccd1 _26015_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1277 _16737_/Y vssd1 vssd1 vccd1 vccd1 _25544_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1288 _25086_/Q vssd1 vssd1 vccd1 vccd1 _18435_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 _12975_/X vssd1 vssd1 vccd1 vccd1 _25045_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23764_ _14797_/B _25993_/Q _23831_/S vssd1 vssd1 vccd1 vccd1 _23764_/X sky130_fd_sc_hd__mux2_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20976_ _21513_/C vssd1 vssd1 vccd1 vccd1 _21516_/B sky130_fd_sc_hd__inv_2
XFILLER_0_170_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25503_ _25510_/CLK hold913/X vssd1 vssd1 vccd1 vccd1 hold912/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22715_ _22937_/A _22715_/B vssd1 vssd1 vccd1 vccd1 _22715_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23695_ _23695_/A vssd1 vssd1 vccd1 vccd1 _25970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25434_ _26002_/CLK _25434_/D vssd1 vssd1 vccd1 vccd1 _25434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22646_ _22646_/A _22646_/B vssd1 vssd1 vccd1 vccd1 _23136_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25365_ _26193_/CLK hold316/X vssd1 vssd1 vccd1 vccd1 hold314/A sky130_fd_sc_hd__dfxtp_1
X_22577_ _22653_/A _22577_/B vssd1 vssd1 vccd1 vccd1 _22577_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_114_clk clkbuf_4_14__f_clk/X vssd1 vssd1 vccd1 vccd1 _26334_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_180_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24316_ _24316_/A vssd1 vssd1 vccd1 vccd1 _26170_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21528_ _21530_/A _21579_/A vssd1 vssd1 vccd1 vccd1 _21529_/B sky130_fd_sc_hd__nand2_1
X_25296_ _26249_/CLK hold286/X vssd1 vssd1 vccd1 vccd1 hold284/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24247_ _24247_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24248_/A sky130_fd_sc_hd__and2_1
XFILLER_0_133_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21459_ _21459_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21459_/Y sky130_fd_sc_hd__nand2_1
X_14000_ _14000_/A hold554/X vssd1 vssd1 vccd1 vccd1 hold555/A sky130_fd_sc_hd__nand2_1
XFILLER_0_181_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24178_ hold2157/X _26126_/Q _24203_/S vssd1 vssd1 vccd1 vccd1 _24178_/X sky130_fd_sc_hd__mux2_1
X_23129_ _23129_/A _23193_/B _23129_/C vssd1 vssd1 vccd1 vccd1 _23129_/X sky130_fd_sc_hd__and3_1
XFILLER_0_101_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15951_ _15951_/A _15951_/B vssd1 vssd1 vccd1 vccd1 _15952_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14902_ _14903_/B _14903_/A vssd1 vssd1 vccd1 vccd1 _14902_/Y sky130_fd_sc_hd__nor2_1
X_15882_ _15882_/A _15882_/B vssd1 vssd1 vccd1 vccd1 _15894_/B sky130_fd_sc_hd__nand2_1
X_18670_ _18952_/A _19824_/B _18891_/C vssd1 vssd1 vccd1 vccd1 _18671_/C sky130_fd_sc_hd__nand3_1
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2490 _15646_/Y vssd1 vssd1 vccd1 vccd1 _25465_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ _17619_/Y _17620_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _17621_/Y sky130_fd_sc_hd__a21oi_1
X_14833_ _15839_/A _25996_/Q vssd1 vssd1 vccd1 vccd1 _22204_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14764_ _14764_/A vssd1 vssd1 vccd1 vccd1 _14955_/A sky130_fd_sc_hd__inv_2
X_17552_ _17552_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17552_/Y sky130_fd_sc_hd__nand2_1
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16503_ _16524_/A _16503_/B vssd1 vssd1 vccd1 vccd1 _16513_/A sky130_fd_sc_hd__or2_1
X_13715_ _26252_/Q _13612_/X _13605_/X _13714_/Y vssd1 vssd1 vccd1 vccd1 _13716_/B
+ sky130_fd_sc_hd__a22o_1
X_17483_ _17481_/Y _17482_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _25621_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14695_ _22680_/A vssd1 vssd1 vccd1 vccd1 _22893_/A sky130_fd_sc_hd__buf_8
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19222_ _20957_/A vssd1 vssd1 vccd1 vccd1 _19222_/X sky130_fd_sc_hd__buf_12
X_16434_ hold866/X vssd1 vssd1 vccd1 vccd1 _16437_/B sky130_fd_sc_hd__inv_2
XFILLER_0_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13646_ _26241_/Q _13612_/X _13605_/X _13645_/Y vssd1 vssd1 vccd1 vccd1 _13647_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _16365_/A _16378_/A vssd1 vssd1 vccd1 vccd1 _16374_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19153_ _26216_/Q hold413/X vssd1 vssd1 vccd1 vccd1 _19153_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_82_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_105_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _25491_/CLK sky130_fd_sc_hd__clkbuf_16
X_13577_ _13583_/A _13577_/B vssd1 vssd1 vccd1 vccd1 _13577_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15316_ _15316_/A _15776_/B vssd1 vssd1 vccd1 vccd1 _15317_/B sky130_fd_sc_hd__nand2_2
X_18104_ _18104_/A _20882_/A vssd1 vssd1 vccd1 vccd1 _18494_/A sky130_fd_sc_hd__xor2_4
X_12528_ _22829_/A _12535_/A vssd1 vssd1 vccd1 vccd1 _17008_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_48_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16296_ _16296_/A vssd1 vssd1 vccd1 vccd1 _16309_/B sky130_fd_sc_hd__inv_2
XFILLER_0_82_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19084_ _19084_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _19084_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_87_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15247_ _16761_/A _15247_/B vssd1 vssd1 vccd1 vccd1 _15248_/B sky130_fd_sc_hd__and2_1
XFILLER_0_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18035_ _18035_/A _18035_/B _18035_/C vssd1 vssd1 vccd1 vccd1 _22221_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15178_ _15178_/A _15178_/B vssd1 vssd1 vccd1 vccd1 _15184_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_140_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14129_ _26318_/Q _13988_/X _13981_/X _14128_/Y vssd1 vssd1 vccd1 vccd1 _14130_/B
+ sky130_fd_sc_hd__a22o_1
X_19986_ _22586_/A vssd1 vssd1 vccd1 vccd1 _20660_/A sky130_fd_sc_hd__buf_8
XFILLER_0_123_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18937_ _20050_/B _22694_/A vssd1 vssd1 vccd1 vccd1 _20043_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_185_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18868_ _25897_/Q _22614_/A vssd1 vssd1 vccd1 vccd1 _18876_/A sky130_fd_sc_hd__or2_2
XFILLER_0_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17819_ _18535_/A _17819_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _17819_/X sky130_fd_sc_hd__and3_1
XFILLER_0_59_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18799_ _19026_/A _18799_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18799_/X sky130_fd_sc_hd__and3_1
XFILLER_0_90_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20830_ _20833_/A _20833_/C vssd1 vssd1 vccd1 vccd1 _20831_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20761_ _21400_/C _21677_/B vssd1 vssd1 vccd1 vccd1 _20764_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_187_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22500_ _22500_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _22500_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23480_ _23474_/X _23479_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _23480_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_92_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20692_ _26294_/Q _20078_/X hold760/X vssd1 vssd1 vccd1 vccd1 _20695_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22431_ _22420_/Y _22429_/Y _23197_/A vssd1 vssd1 vccd1 vccd1 _22431_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25150_ _26234_/CLK hold457/X vssd1 vssd1 vccd1 vccd1 hold455/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22362_ _22346_/X _22361_/Y _17229_/B vssd1 vssd1 vccd1 vccd1 _22362_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24101_ _24101_/A vssd1 vssd1 vccd1 vccd1 _26100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21313_ _21313_/A _21313_/B vssd1 vssd1 vccd1 vccd1 _21314_/A sky130_fd_sc_hd__nand2_1
X_25081_ _26164_/CLK _25081_/D vssd1 vssd1 vccd1 vccd1 _25081_/Q sky130_fd_sc_hd__dfxtp_1
X_22293_ _22293_/A _22387_/B vssd1 vssd1 vccd1 vccd1 _22293_/Y sky130_fd_sc_hd__nand2_1
X_24032_ hold2494/X hold2389/X _24047_/S vssd1 vssd1 vccd1 vccd1 _24033_/A sky130_fd_sc_hd__mux2_1
Xhold330 hold330/A vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__dlygate4sd3_1
X_21244_ _21243_/B _21244_/B _21244_/C vssd1 vssd1 vccd1 vccd1 _21245_/B sky130_fd_sc_hd__nand3b_1
Xhold341 hold341/A vssd1 vssd1 vccd1 vccd1 hold341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 hold352/A vssd1 vssd1 vccd1 vccd1 hold352/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 hold363/A vssd1 vssd1 vccd1 vccd1 hold363/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold374 hold374/A vssd1 vssd1 vccd1 vccd1 hold374/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 hold385/A vssd1 vssd1 vccd1 vccd1 hold385/X sky130_fd_sc_hd__dlygate4sd3_1
X_21175_ _26310_/Q _20731_/X hold488/X vssd1 vssd1 vccd1 vccd1 _21178_/B sky130_fd_sc_hd__a21oi_1
Xhold396 hold396/A vssd1 vssd1 vccd1 vccd1 hold396/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20126_ _21042_/A _20126_/B _20125_/X vssd1 vssd1 vccd1 vccd1 _20127_/B sky130_fd_sc_hd__or3b_1
X_25983_ _26004_/CLK _25983_/D vssd1 vssd1 vccd1 vccd1 _25983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24934_ _24946_/A _24934_/B vssd1 vssd1 vccd1 vccd1 _24934_/Y sky130_fd_sc_hd__nor2_1
X_20057_ _20057_/A _22821_/B vssd1 vssd1 vccd1 vccd1 _20062_/A sky130_fd_sc_hd__nand2_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1030 _16751_/Y vssd1 vssd1 vccd1 vccd1 _25546_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1041 _25016_/Q vssd1 vssd1 vccd1 vccd1 _17214_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1052 _16540_/Y vssd1 vssd1 vccd1 vccd1 _25527_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24865_ _24944_/S _25460_/Q _24864_/Y vssd1 vssd1 vccd1 vccd1 _24865_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1063 _25036_/Q vssd1 vssd1 vccd1 vccd1 _17442_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1074 _13437_/X vssd1 vssd1 vccd1 vccd1 _25124_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1085 _25564_/Q vssd1 vssd1 vccd1 vccd1 _16872_/B sky130_fd_sc_hd__buf_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23816_ _24560_/A vssd1 vssd1 vccd1 vccd1 _23905_/B sky130_fd_sc_hd__buf_6
Xhold1096 _13087_/X vssd1 vssd1 vccd1 vccd1 _25066_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24796_ hold2691/X _26327_/Q _24817_/S vssd1 vssd1 vccd1 vccd1 _24796_/X sky130_fd_sc_hd__mux2_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23747_ _23747_/A vssd1 vssd1 vccd1 vccd1 _25987_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20959_ _21042_/A _20959_/B _20958_/X vssd1 vssd1 vccd1 vccd1 _20960_/B sky130_fd_sc_hd__or3b_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13500_ _13500_/A _13518_/B vssd1 vssd1 vccd1 vccd1 _13500_/Y sky130_fd_sc_hd__nor2_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14525_/A hold197/X vssd1 vssd1 vccd1 vccd1 hold198/A sky130_fd_sc_hd__nand2_1
X_23678_ _23678_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23679_/A sky130_fd_sc_hd__and2_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25417_ _25418_/CLK _25417_/D vssd1 vssd1 vccd1 vccd1 _25417_/Q sky130_fd_sc_hd__dfxtp_1
X_13431_ _19040_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13431_/X sky130_fd_sc_hd__or2_1
X_22629_ _15242_/B _22387_/B _14273_/X vssd1 vssd1 vccd1 vccd1 _22629_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16150_ _16150_/A _16150_/B vssd1 vssd1 vccd1 vccd1 _16152_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13362_ _26195_/Q _13239_/X _13361_/X vssd1 vssd1 vccd1 vccd1 _13362_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_24_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25348_ _26175_/CLK hold163/X vssd1 vssd1 vccd1 vccd1 hold161/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15101_ _15101_/A _15101_/B vssd1 vssd1 vccd1 vccd1 _15106_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_122_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16081_ _16081_/A _16081_/B vssd1 vssd1 vccd1 vccd1 _16082_/B sky130_fd_sc_hd__nand2_1
X_25279_ _26232_/CLK hold340/X vssd1 vssd1 vccd1 vccd1 hold338/A sky130_fd_sc_hd__dfxtp_1
X_13293_ _18739_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13293_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15032_ _15032_/A _15032_/B _15032_/C vssd1 vssd1 vccd1 vccd1 _15033_/B sky130_fd_sc_hd__and3_1
XFILLER_0_107_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19840_ _26264_/Q _19134_/X hold521/X vssd1 vssd1 vccd1 vccd1 _19840_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19771_ _26259_/Q hold500/X vssd1 vssd1 vccd1 vccd1 _19771_/Y sky130_fd_sc_hd__nand2_1
X_16983_ _23191_/B _16773_/A hold1226/X _16982_/Y _14345_/A vssd1 vssd1 vccd1 vccd1
+ _16983_/Y sky130_fd_sc_hd__a221oi_1
X_18722_ _18986_/A _19518_/A vssd1 vssd1 vccd1 vccd1 _18722_/Y sky130_fd_sc_hd__nand2_1
X_15934_ _15934_/A _15934_/B vssd1 vssd1 vccd1 vccd1 _15936_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18653_ _18653_/A _18653_/B _18653_/C vssd1 vssd1 vccd1 vccd1 _22350_/A sky130_fd_sc_hd__nand3_2
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15865_ _15866_/B _15866_/A vssd1 vssd1 vccd1 vccd1 _15884_/C sky130_fd_sc_hd__or2_1
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17604_ _17604_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _17604_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_153_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14816_ _14822_/B _22145_/A vssd1 vssd1 vccd1 vccd1 _22144_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_189_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18584_ _20236_/B _19673_/A vssd1 vssd1 vccd1 vccd1 _18585_/B sky130_fd_sc_hd__nand2_1
X_15796_ hold902/X _15798_/A vssd1 vssd1 vccd1 vccd1 _15800_/A sky130_fd_sc_hd__nor2_1
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17535_ _17535_/A _17535_/B vssd1 vssd1 vccd1 vccd1 _17535_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_98_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14747_ _25843_/Q _12527_/A _14938_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14747_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14678_ _14678_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _14678_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17466_ _17466_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17466_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_67_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19205_ _19205_/A _19980_/B _19205_/C vssd1 vssd1 vccd1 vccd1 _19205_/X sky130_fd_sc_hd__and3_1
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16417_ _16403_/A _16389_/A _16402_/B vssd1 vssd1 vccd1 vccd1 _16417_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_144_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13629_ hold495/X _13628_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold496/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_183_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17397_ _17395_/Y _17396_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _17397_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19136_ _19136_/A _23195_/B _19136_/C vssd1 vssd1 vccd1 vccd1 _19136_/X sky130_fd_sc_hd__and3_1
X_16348_ _16361_/B vssd1 vssd1 vccd1 vccd1 _16351_/B sky130_fd_sc_hd__inv_2
XFILLER_0_54_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16279_ _16279_/A _16279_/B vssd1 vssd1 vccd1 vccd1 _16490_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19067_ _19067_/A _19067_/B vssd1 vssd1 vccd1 vccd1 _19067_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18018_ _17761_/B _17760_/B _17973_/B vssd1 vssd1 vccd1 vccd1 _18019_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_120_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19969_ _19969_/A _19980_/B _19969_/C vssd1 vssd1 vccd1 vccd1 _19969_/X sky130_fd_sc_hd__and3_1
X_22980_ _15583_/B _22680_/X _22829_/X vssd1 vssd1 vccd1 vccd1 _22980_/Y sky130_fd_sc_hd__a21oi_1
X_21931_ _22058_/A _21931_/B vssd1 vssd1 vccd1 vccd1 _21931_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24650_ _24650_/A vssd1 vssd1 vccd1 vccd1 _26279_/D sky130_fd_sc_hd__clkbuf_1
X_21862_ _22058_/A _21862_/B vssd1 vssd1 vccd1 vccd1 _21862_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23601_ _23599_/B _23598_/B _23599_/Y _23600_/X _12515_/X vssd1 vssd1 vccd1 vccd1
+ _23602_/A sky130_fd_sc_hd__a221o_4
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20813_ _20813_/A _20813_/B vssd1 vssd1 vccd1 vccd1 _20814_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24581_ hold2707/X hold2701/X _24587_/S vssd1 vssd1 vccd1 vccd1 _24582_/A sky130_fd_sc_hd__mux2_1
X_21793_ _22058_/A _21793_/B vssd1 vssd1 vccd1 vccd1 _21793_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_78_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26320_ _26325_/CLK _26320_/D vssd1 vssd1 vccd1 vccd1 _26320_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23532_ _23508_/X _23531_/X _25912_/Q vssd1 vssd1 vccd1 vccd1 _23532_/X sky130_fd_sc_hd__mux2_2
X_20744_ _25857_/Q vssd1 vssd1 vccd1 vccd1 _21734_/B sky130_fd_sc_hd__inv_2
XFILLER_0_33_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26251_ _26251_/CLK _26251_/D vssd1 vssd1 vccd1 vccd1 _26251_/Q sky130_fd_sc_hd__dfxtp_2
X_23463_ _23460_/Y _23462_/Y _24957_/S vssd1 vssd1 vccd1 vccd1 _23463_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_161_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20675_ _20675_/A _25894_/Q vssd1 vssd1 vccd1 vccd1 _20681_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_163_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25202_ _26239_/CLK hold391/X vssd1 vssd1 vccd1 vccd1 hold389/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22414_ _22414_/A _22414_/B vssd1 vssd1 vccd1 vccd1 _22992_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_18_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26182_ _26184_/CLK _26182_/D vssd1 vssd1 vccd1 vccd1 _26182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23394_ _23390_/Y _23393_/Y _24858_/S vssd1 vssd1 vccd1 vccd1 _23394_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25133_ _25135_/CLK hold415/X vssd1 vssd1 vccd1 vccd1 hold413/A sky130_fd_sc_hd__dfxtp_1
X_22345_ _22343_/X _15839_/B _22344_/Y _14882_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _22346_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_131_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25064_ _25712_/CLK _25064_/D vssd1 vssd1 vccd1 vccd1 _25064_/Q sky130_fd_sc_hd__dfxtp_1
X_22276_ _22743_/A _22890_/B vssd1 vssd1 vccd1 vccd1 _22287_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24015_ _24015_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24016_/A sky130_fd_sc_hd__and2_1
Xhold160 hold160/A vssd1 vssd1 vccd1 vccd1 hold160/X sky130_fd_sc_hd__dlygate4sd3_1
X_21227_ _21227_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _21233_/A sky130_fd_sc_hd__nand2_1
Xhold171 hold171/A vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 hold182/A vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 hold193/A vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
X_21158_ _21160_/B _21160_/C vssd1 vssd1 vccd1 vccd1 _21159_/A sky130_fd_sc_hd__nand2_1
X_20109_ _21402_/A vssd1 vssd1 vccd1 vccd1 _21401_/A sky130_fd_sc_hd__inv_2
X_13980_ _14000_/A hold718/X vssd1 vssd1 vccd1 vccd1 hold719/A sky130_fd_sc_hd__nand2_1
X_25966_ _26042_/CLK _25966_/D vssd1 vssd1 vccd1 vccd1 _25966_/Q sky130_fd_sc_hd__dfxtp_1
X_21089_ _21089_/A _21089_/B _21089_/C vssd1 vssd1 vccd1 vccd1 _21090_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_137_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12931_ _26248_/Q _25617_/Q vssd1 vssd1 vccd1 vccd1 _14397_/A sky130_fd_sc_hd__xor2_1
X_24917_ _24946_/A _24917_/B vssd1 vssd1 vccd1 vccd1 _24917_/Y sky130_fd_sc_hd__nor2_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25897_ _26080_/CLK _25897_/D vssd1 vssd1 vccd1 vccd1 _25897_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ _23047_/B _15650_/B vssd1 vssd1 vccd1 vccd1 _23044_/B sky130_fd_sc_hd__xor2_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ _12726_/B _14358_/A _12752_/X _25604_/Q vssd1 vssd1 vccd1 vccd1 _12862_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24848_ _15373_/B _15387_/B _24860_/S vssd1 vssd1 vccd1 vccd1 _24848_/X sky130_fd_sc_hd__mux2_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _14599_/Y hold369/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold370/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15581_ _26031_/Q _25967_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15582_/A sky130_fd_sc_hd__mux2_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _26222_/Q _25591_/Q vssd1 vssd1 vccd1 vccd1 _14316_/A sky130_fd_sc_hd__xor2_2
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24779_ _24779_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24780_/A sky130_fd_sc_hd__and2_1
XFILLER_0_185_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14532_ _14529_/Y hold228/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold229/A sky130_fd_sc_hd__a21oi_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _17571_/A _17651_/A vssd1 vssd1 vccd1 vccd1 _17321_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14463_ _14461_/Y hold30/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__a21oi_1
X_17251_ _25640_/Q vssd1 vssd1 vccd1 vccd1 _20752_/B sky130_fd_sc_hd__inv_2
XFILLER_0_126_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16202_ _16200_/X _16201_/Y _16076_/X vssd1 vssd1 vccd1 vccd1 _25502_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13414_ _26332_/Q _19816_/A vssd1 vssd1 vccd1 vccd1 _14663_/A sky130_fd_sc_hd__xor2_1
X_17182_ _25635_/Q vssd1 vssd1 vccd1 vccd1 _20558_/B sky130_fd_sc_hd__inv_2
X_14394_ _14394_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14394_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_180_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16133_ _16133_/A _16133_/B vssd1 vssd1 vccd1 vccd1 _16135_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_141_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13345_ _18900_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13345_/X sky130_fd_sc_hd__or2_1
XFILLER_0_148_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16064_ _16212_/A hold800/X vssd1 vssd1 vccd1 vccd1 hold801/A sky130_fd_sc_hd__nand2_1
XFILLER_0_122_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13276_ _13207_/X _13274_/X _13192_/X _13275_/X vssd1 vssd1 vccd1 vccd1 _13276_/X
+ sky130_fd_sc_hd__o211a_1
X_15015_ _15015_/A _15015_/B vssd1 vssd1 vccd1 vccd1 _15030_/A sky130_fd_sc_hd__nor2_1
X_19823_ _19815_/X _19822_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19823_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19754_ _26258_/Q _19134_/X hold524/X vssd1 vssd1 vccd1 vccd1 _19754_/Y sky130_fd_sc_hd__a21oi_1
X_16966_ _16967_/B _16967_/A vssd1 vssd1 vccd1 vccd1 _16966_/X sky130_fd_sc_hd__or2_1
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18705_ _22408_/B _25633_/Q vssd1 vssd1 vccd1 vccd1 _18707_/A sky130_fd_sc_hd__nand2_1
X_15917_ _15918_/B _15918_/A vssd1 vssd1 vccd1 vccd1 _15934_/B sky130_fd_sc_hd__or2_1
XFILLER_0_189_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19685_ _19684_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19686_/B
+ sky130_fd_sc_hd__a211o_1
X_16897_ _16897_/A _16897_/B vssd1 vssd1 vccd1 vccd1 _16897_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_182_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18636_ _18838_/A _18966_/A vssd1 vssd1 vccd1 vccd1 _18637_/B sky130_fd_sc_hd__xnor2_1
X_15848_ _15857_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _15848_/Y sky130_fd_sc_hd__nand2_1
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18567_ _18792_/A _18571_/B vssd1 vssd1 vccd1 vccd1 _18569_/A sky130_fd_sc_hd__nand2_1
X_15779_ _15780_/B _16967_/A vssd1 vssd1 vccd1 vccd1 _15781_/A sky130_fd_sc_hd__or2_1
XFILLER_0_74_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17518_ _17516_/Y _17517_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _17518_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18498_ _18641_/A _19359_/A vssd1 vssd1 vccd1 vccd1 _18498_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17449_ _17624_/A _17449_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17449_/X sky130_fd_sc_hd__and3_1
XFILLER_0_89_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20460_ _20459_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20460_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_172_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19119_ _19961_/B _19220_/A vssd1 vssd1 vccd1 vccd1 _19120_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20391_ _20394_/A _20394_/C vssd1 vssd1 vccd1 vccd1 _20392_/A sky130_fd_sc_hd__nand2_1
X_22130_ _22130_/A _25850_/Q vssd1 vssd1 vccd1 vccd1 _22130_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_112_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22061_ _22061_/A _22145_/B vssd1 vssd1 vccd1 vccd1 _22061_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21012_ _21012_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _21017_/A sky130_fd_sc_hd__nand2_1
X_25820_ _25822_/CLK _25820_/D vssd1 vssd1 vccd1 vccd1 _25820_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25751_ _25752_/CLK _25751_/D vssd1 vssd1 vccd1 vccd1 _25751_/Q sky130_fd_sc_hd__dfxtp_1
X_22963_ _15566_/B _22680_/X _22829_/X vssd1 vssd1 vccd1 vccd1 _22963_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_94_clk clkbuf_leaf_95_clk/A vssd1 vssd1 vccd1 vccd1 _26002_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24702_ _24702_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24703_/A sky130_fd_sc_hd__and2_1
X_21914_ _18350_/A _25807_/Q _21912_/Y _21913_/Y vssd1 vssd1 vccd1 vccd1 _21915_/B
+ sky130_fd_sc_hd__a31o_1
X_25682_ _25687_/CLK _25682_/D vssd1 vssd1 vccd1 vccd1 _25682_/Q sky130_fd_sc_hd__dfxtp_1
X_22894_ _15490_/B _16980_/A _14273_/X vssd1 vssd1 vccd1 vccd1 _22894_/Y sky130_fd_sc_hd__a21oi_1
X_24633_ hold2733/X hold2720/X _24664_/S vssd1 vssd1 vccd1 vccd1 _24634_/A sky130_fd_sc_hd__mux2_1
X_21845_ _18310_/A _21844_/A _21843_/Y _21844_/Y vssd1 vssd1 vccd1 vccd1 _21846_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24564_ _24564_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24565_/A sky130_fd_sc_hd__and2_1
XFILLER_0_65_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21776_ _19444_/A _21775_/A _21775_/Y vssd1 vssd1 vccd1 vccd1 _21778_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23515_ _24944_/S hold374/A _23514_/X vssd1 vssd1 vccd1 vccd1 _23515_/Y sky130_fd_sc_hd__o21ai_1
X_26303_ _26303_/CLK _26303_/D vssd1 vssd1 vccd1 vccd1 _26303_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_135_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20727_ _21387_/B _21661_/B vssd1 vssd1 vccd1 vccd1 _20728_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_135_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24495_ hold2600/X _26229_/Q _24510_/S vssd1 vssd1 vccd1 vccd1 _24495_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26234_ _26234_/CLK _26234_/D vssd1 vssd1 vccd1 vccd1 _26234_/Q sky130_fd_sc_hd__dfxtp_1
X_23446_ hold14/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23446_/X sky130_fd_sc_hd__or2b_1
X_20658_ _20658_/A _20658_/B vssd1 vssd1 vccd1 vccd1 _20659_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_151_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26165_ _26297_/CLK _26165_/D vssd1 vssd1 vccd1 vccd1 _26165_/Q sky130_fd_sc_hd__dfxtp_1
X_23377_ _23377_/A _23377_/B _23380_/A vssd1 vssd1 vccd1 vccd1 _23377_/X sky130_fd_sc_hd__and3_1
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20589_ _25853_/Q vssd1 vssd1 vccd1 vccd1 _22224_/B sky130_fd_sc_hd__inv_2
XFILLER_0_34_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25116_ _26200_/CLK _25116_/D vssd1 vssd1 vccd1 vccd1 _25116_/Q sky130_fd_sc_hd__dfxtp_1
X_13130_ _26286_/Q _25655_/Q vssd1 vssd1 vccd1 vccd1 _14518_/A sky130_fd_sc_hd__xor2_2
X_22328_ _18635_/A _25821_/Q _22326_/Y _22327_/Y vssd1 vssd1 vccd1 vccd1 _22329_/B
+ sky130_fd_sc_hd__a31o_1
X_26096_ _26096_/CLK _26096_/D vssd1 vssd1 vccd1 vccd1 _26096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25047_ _26135_/CLK hold901/X vssd1 vssd1 vccd1 vccd1 _25047_/Q sky130_fd_sc_hd__dfxtp_1
X_13061_ _13049_/X _14479_/A _12909_/X _25642_/Q vssd1 vssd1 vccd1 vccd1 _13061_/X
+ sky130_fd_sc_hd__a22o_1
X_22259_ _22235_/X _22258_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _22259_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16820_ _16858_/A _16820_/B vssd1 vssd1 vccd1 vccd1 _16820_/Y sky130_fd_sc_hd__nand2_1
X_16751_ _16749_/Y _16750_/Y _16594_/X vssd1 vssd1 vccd1 vccd1 _16751_/Y sky130_fd_sc_hd__a21oi_1
X_25949_ _26014_/CLK _25949_/D vssd1 vssd1 vccd1 vccd1 _25949_/Q sky130_fd_sc_hd__dfxtp_1
X_13963_ _25789_/Q vssd1 vssd1 vccd1 vccd1 _18035_/B sky130_fd_sc_hd__inv_2
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_85_clk clkbuf_leaf_95_clk/A vssd1 vssd1 vccd1 vccd1 _25875_/CLK sky130_fd_sc_hd__clkbuf_16
X_15702_ _15700_/X hold2444/X _15464_/X vssd1 vssd1 vccd1 vccd1 _15702_/Y sky130_fd_sc_hd__a21oi_1
X_19470_ _26238_/Q hold494/X vssd1 vssd1 vccd1 vccd1 _19470_/Y sky130_fd_sc_hd__nand2_1
X_12914_ _26245_/Q _25614_/Q vssd1 vssd1 vccd1 vccd1 _14388_/A sky130_fd_sc_hd__xor2_1
X_16682_ _16670_/B _16680_/A _16668_/A vssd1 vssd1 vccd1 vccd1 _16683_/B sky130_fd_sc_hd__o21a_1
X_13894_ _14000_/A hold557/X vssd1 vssd1 vccd1 vccd1 hold558/A sky130_fd_sc_hd__nand2_1
X_18421_ _22040_/B _25619_/Q vssd1 vssd1 vccd1 vccd1 _18423_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_159_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15633_ _26034_/Q _25970_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15634_/A sky130_fd_sc_hd__mux2_1
X_12845_ _12840_/X _12843_/X _12827_/X _12844_/X vssd1 vssd1 vccd1 vccd1 _12845_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _19080_/A _18352_/B vssd1 vssd1 vccd1 vccd1 _18352_/X sky130_fd_sc_hd__xor2_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15564_ _26030_/Q _25966_/Q _15773_/S vssd1 vssd1 vccd1 vccd1 _15565_/A sky130_fd_sc_hd__mux2_1
X_12776_ _25007_/Q _14264_/A vssd1 vssd1 vccd1 vccd1 _12776_/X sky130_fd_sc_hd__or2_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _19430_/A _17303_/B vssd1 vssd1 vccd1 vccd1 _17563_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_167_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14515_ _14515_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14515_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15495_ _16855_/A _15495_/B vssd1 vssd1 vccd1 vccd1 _15496_/B sky130_fd_sc_hd__and2_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18283_ _18283_/A _25804_/Q _18283_/C vssd1 vssd1 vccd1 vccd1 _21080_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_72_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17234_ _19359_/A _17234_/B vssd1 vssd1 vccd1 vccd1 _17527_/A sky130_fd_sc_hd__xor2_4
X_14446_ _14446_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14446_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17165_ _17163_/Y _17164_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _25592_/D sky130_fd_sc_hd__a21oi_1
X_14377_ _14404_/A hold242/X vssd1 vssd1 vccd1 vccd1 hold243/A sky130_fd_sc_hd__nand2_1
XFILLER_0_80_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold907 hold907/A vssd1 vssd1 vccd1 vccd1 hold907/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold918 hold918/A vssd1 vssd1 vccd1 vccd1 hold918/X sky130_fd_sc_hd__dlygate4sd3_1
X_16116_ _16125_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16116_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13328_ _13315_/X _13325_/X _13300_/X _13327_/X vssd1 vssd1 vccd1 vccd1 _13328_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold929 hold929/A vssd1 vssd1 vccd1 vccd1 hold929/X sky130_fd_sc_hd__dlygate4sd3_1
X_17096_ _17272_/A _17096_/B vssd1 vssd1 vccd1 vccd1 _17096_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_51_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16047_ _22232_/B _16691_/B vssd1 vssd1 vccd1 vccd1 _16049_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_122_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13259_ _13259_/A vssd1 vssd1 vccd1 vccd1 _19458_/A sky130_fd_sc_hd__buf_4
XFILLER_0_23_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2308 _24157_/X vssd1 vssd1 vccd1 vccd1 _24158_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2319 _25661_/Q vssd1 vssd1 vccd1 vccd1 _13164_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19806_ _19807_/B _19807_/A vssd1 vssd1 vccd1 vccd1 _19806_/X sky130_fd_sc_hd__or2_1
Xhold1607 _21289_/Y vssd1 vssd1 vccd1 vccd1 _25811_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1618 _25824_/Q vssd1 vssd1 vccd1 vccd1 _21509_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17998_ _18611_/A _18002_/B vssd1 vssd1 vccd1 vccd1 _18000_/A sky130_fd_sc_hd__nand2_1
Xhold1629 _21672_/Y vssd1 vssd1 vccd1 vccd1 _25834_/D sky130_fd_sc_hd__dlygate4sd3_1
X_19737_ _22586_/A vssd1 vssd1 vccd1 vccd1 _19975_/A sky130_fd_sc_hd__buf_6
X_16949_ _16977_/A _16949_/B vssd1 vssd1 vccd1 vccd1 _16949_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_76_clk clkbuf_leaf_82_clk/A vssd1 vssd1 vccd1 vccd1 _25838_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19668_ _19666_/Y _19667_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19668_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18619_ _18617_/X _18269_/X _18618_/X vssd1 vssd1 vccd1 vccd1 _18620_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_177_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19599_ _26247_/Q hold614/X vssd1 vssd1 vccd1 vccd1 _19599_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_176_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21630_ _21630_/A _21630_/B _21630_/C vssd1 vssd1 vccd1 vccd1 _21631_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21561_ _21561_/A _21561_/B _21561_/C vssd1 vssd1 vccd1 vccd1 _21565_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_129_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23300_ _23300_/A vssd1 vssd1 vccd1 vccd1 _25922_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20512_ _20514_/B _20514_/C vssd1 vssd1 vccd1 vccd1 _20513_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24280_ _24280_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24281_/A sky130_fd_sc_hd__and2_1
XFILLER_0_51_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21492_ _21573_/A _21492_/B vssd1 vssd1 vccd1 vccd1 _21492_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_105_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23231_ _23231_/A _24867_/S vssd1 vssd1 vccd1 vccd1 _23234_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_117_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20443_ _20443_/A _22396_/B _20443_/C vssd1 vssd1 vccd1 vccd1 _20447_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_16_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23162_ _16970_/B _22421_/A _23156_/X _23157_/Y _23161_/X vssd1 vssd1 vccd1 vccd1
+ _23163_/A sky130_fd_sc_hd__a221o_1
X_20374_ _21514_/A _21195_/C vssd1 vssd1 vccd1 vccd1 _20375_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22113_ _22561_/A _22113_/B vssd1 vssd1 vccd1 vccd1 _22113_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_113_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23093_ _15707_/B _22893_/A _22829_/X vssd1 vssd1 vccd1 vccd1 _23093_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22044_ _22772_/B _22045_/A vssd1 vssd1 vccd1 vccd1 _22046_/A sky130_fd_sc_hd__or2_1
XFILLER_0_167_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25803_ _25803_/CLK _25803_/D vssd1 vssd1 vccd1 vccd1 _25803_/Q sky130_fd_sc_hd__dfxtp_1
X_23995_ _26066_/Q hold2478/X _24001_/S vssd1 vssd1 vccd1 vccd1 _23995_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_67_clk _25472_/CLK vssd1 vssd1 vccd1 vccd1 _25877_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22946_ _15540_/B _22680_/X _22829_/X vssd1 vssd1 vccd1 vccd1 _22946_/Y sky130_fd_sc_hd__a21oi_1
X_25734_ _25796_/CLK _25734_/D vssd1 vssd1 vccd1 vccd1 _25734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22877_ _23026_/A _22877_/B vssd1 vssd1 vccd1 vccd1 _22878_/A sky130_fd_sc_hd__xor2_1
X_25665_ _26296_/CLK _25665_/D vssd1 vssd1 vccd1 vccd1 _25665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12630_ _12630_/A _24836_/B _12635_/A vssd1 vssd1 vccd1 vccd1 _12630_/X sky130_fd_sc_hd__and3_1
XFILLER_0_78_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21828_ _22058_/A _21828_/B vssd1 vssd1 vccd1 vccd1 _21828_/Y sky130_fd_sc_hd__nand2_1
X_24616_ _24616_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24617_/A sky130_fd_sc_hd__and2_1
XFILLER_0_183_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25596_ _25596_/CLK _25596_/D vssd1 vssd1 vccd1 vccd1 _25596_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12561_ _12561_/A vssd1 vssd1 vccd1 vccd1 _24965_/D sky130_fd_sc_hd__clkbuf_1
X_24547_ hold2647/X hold2642/X _24587_/S vssd1 vssd1 vccd1 vccd1 _24548_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_164_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21759_ _22893_/A _21759_/B vssd1 vssd1 vccd1 vccd1 _21759_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14300_ _14298_/Y hold183/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold184/A sky130_fd_sc_hd__a21oi_1
X_15280_ _15278_/X _15279_/Y _15090_/X vssd1 vssd1 vccd1 vccd1 _25444_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12492_ _23193_/B vssd1 vssd1 vccd1 vccd1 _23001_/B sky130_fd_sc_hd__buf_8
X_24478_ _24478_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24479_/A sky130_fd_sc_hd__and2_1
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14231_ _25832_/Q vssd1 vssd1 vccd1 vccd1 _18854_/B sky130_fd_sc_hd__inv_2
XFILLER_0_184_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26217_ _26219_/CLK _26217_/D vssd1 vssd1 vccd1 vccd1 _26217_/Q sky130_fd_sc_hd__dfxtp_2
X_23429_ _23426_/Y _23428_/Y _24858_/S vssd1 vssd1 vccd1 vccd1 _23429_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_163_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26148_ _26148_/CLK _26148_/D vssd1 vssd1 vccd1 vccd1 _26148_/Q sky130_fd_sc_hd__dfxtp_1
X_14162_ hold648/X _14161_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold649/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13113_ _18058_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13113_/X sky130_fd_sc_hd__or2_1
X_26079_ _26079_/CLK _26079_/D vssd1 vssd1 vccd1 vccd1 _26079_/Q sky130_fd_sc_hd__dfxtp_1
X_14093_ hold570/X _14092_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold571/A sky130_fd_sc_hd__a21oi_1
X_18970_ _21791_/A vssd1 vssd1 vccd1 vccd1 _19126_/B sky130_fd_sc_hd__buf_8
XFILLER_0_104_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17921_ _21855_/A _25585_/Q vssd1 vssd1 vccd1 vccd1 _17923_/B sky130_fd_sc_hd__nand2_1
X_13044_ _26270_/Q _25639_/Q vssd1 vssd1 vccd1 vccd1 _14469_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17852_ _25593_/Q _22106_/A vssd1 vssd1 vccd1 vccd1 _17853_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_156_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16803_ _16803_/A _16803_/B vssd1 vssd1 vccd1 vccd1 _16803_/Y sky130_fd_sc_hd__nand2_1
X_17783_ _17781_/B _17783_/B _17783_/C vssd1 vssd1 vccd1 vccd1 _17784_/B sky130_fd_sc_hd__nand3b_2
Xclkbuf_leaf_58_clk _25472_/CLK vssd1 vssd1 vccd1 vccd1 _25534_/CLK sky130_fd_sc_hd__clkbuf_16
X_14995_ _14996_/B _14996_/A vssd1 vssd1 vccd1 vccd1 _14997_/A sky130_fd_sc_hd__or2_1
X_19522_ _19523_/B _19523_/A vssd1 vssd1 vccd1 vccd1 _19522_/X sky130_fd_sc_hd__or2_1
X_16734_ _16732_/X _16711_/X _16733_/Y _25865_/Q _14170_/X vssd1 vssd1 vccd1 vccd1
+ _16735_/A sky130_fd_sc_hd__a32o_1
X_13946_ _17896_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13946_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19453_ _19451_/Y _19452_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19453_/Y sky130_fd_sc_hd__a21oi_1
X_16665_ _16665_/A _16691_/B vssd1 vssd1 vccd1 vccd1 _16667_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13877_ _26278_/Q _13801_/X _13793_/X _13876_/Y vssd1 vssd1 vccd1 vccd1 _13878_/B
+ sky130_fd_sc_hd__a22o_1
X_18404_ _18446_/A _25746_/Q _21716_/A vssd1 vssd1 vccd1 vccd1 _18405_/C sky130_fd_sc_hd__nand3_1
X_15616_ _25569_/Q vssd1 vssd1 vccd1 vccd1 _23015_/B sky130_fd_sc_hd__inv_2
XFILLER_0_29_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12828_ _17227_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12828_/X sky130_fd_sc_hd__or2_1
X_19384_ _26232_/Q _12537_/B hold590/X vssd1 vssd1 vccd1 vccd1 _19384_/Y sky130_fd_sc_hd__a21oi_1
X_16596_ _16596_/A _16596_/B vssd1 vssd1 vccd1 vccd1 _16597_/B sky130_fd_sc_hd__and2_1
XFILLER_0_118_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18335_ _18335_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18335_/Y sky130_fd_sc_hd__nand2_1
X_15547_ _15547_/A vssd1 vssd1 vccd1 vccd1 _15548_/B sky130_fd_sc_hd__inv_2
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12759_ _12726_/B _14295_/A _12752_/X _25584_/Q vssd1 vssd1 vccd1 vccd1 _12759_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18266_ _18266_/A _21047_/A vssd1 vssd1 vccd1 vccd1 _18617_/A sky130_fd_sc_hd__xor2_4
X_15478_ hold916/X vssd1 vssd1 vccd1 vccd1 _15480_/A sky130_fd_sc_hd__inv_2
XFILLER_0_155_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17217_ _17272_/A _17217_/B vssd1 vssd1 vccd1 vccd1 _17217_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_13_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14429_ _14465_/A hold239/X vssd1 vssd1 vccd1 vccd1 hold240/A sky130_fd_sc_hd__nand2_1
XFILLER_0_181_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18197_ _25864_/Q _21971_/A vssd1 vssd1 vccd1 vccd1 _18205_/A sky130_fd_sc_hd__or2_2
XFILLER_0_181_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold704 hold704/A vssd1 vssd1 vccd1 vccd1 hold704/X sky130_fd_sc_hd__dlygate4sd3_1
X_17148_ _17393_/A _17148_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17148_/X sky130_fd_sc_hd__and3_1
XFILLER_0_80_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold715 hold715/A vssd1 vssd1 vccd1 vccd1 hold715/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold726 hold726/A vssd1 vssd1 vccd1 vccd1 hold726/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 hold737/A vssd1 vssd1 vccd1 vccd1 hold737/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold748 hold748/A vssd1 vssd1 vccd1 vccd1 hold748/X sky130_fd_sc_hd__dlygate4sd3_1
X_17079_ _17079_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17079_/Y sky130_fd_sc_hd__nand2_1
Xhold759 hold759/A vssd1 vssd1 vccd1 vccd1 hold759/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20090_ _23197_/B vssd1 vssd1 vccd1 vccd1 _22723_/B sky130_fd_sc_hd__inv_2
XFILLER_0_23_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2105 _26010_/Q vssd1 vssd1 vccd1 vccd1 hold2105/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2116 _15080_/Y vssd1 vssd1 vccd1 vccd1 hold2116/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2127 _23935_/X vssd1 vssd1 vccd1 vccd1 _23936_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2138 _23277_/X vssd1 vssd1 vccd1 vccd1 _23279_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1404 _14832_/Y vssd1 vssd1 vccd1 vccd1 _25403_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2149 _15091_/Y vssd1 vssd1 vccd1 vccd1 _25434_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1415 _25720_/Q vssd1 vssd1 vccd1 vccd1 _19268_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1426 _19298_/Y vssd1 vssd1 vccd1 vccd1 _25722_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1437 _25558_/Q vssd1 vssd1 vccd1 vccd1 _16834_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1448 _19541_/Y vssd1 vssd1 vccd1 vccd1 _25739_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_49_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _26021_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1459 _25107_/Q vssd1 vssd1 vccd1 vccd1 _18859_/B sky130_fd_sc_hd__dlygate4sd3_1
X_22800_ _22799_/A _22454_/X _22799_/B vssd1 vssd1 vccd1 vccd1 _22801_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23780_ _23780_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23781_/A sky130_fd_sc_hd__and2_1
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20992_ _20990_/Y _20991_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _20992_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22731_ _23188_/A _22731_/B vssd1 vssd1 vccd1 vccd1 _22731_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25450_ _25450_/CLK _25450_/D vssd1 vssd1 vccd1 vccd1 _25450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22662_ _22937_/A _22662_/B vssd1 vssd1 vccd1 vccd1 _22662_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24401_ _24401_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24402_/A sky130_fd_sc_hd__and2_1
XFILLER_0_164_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21613_ _21613_/A _21613_/B _21613_/C vssd1 vssd1 vccd1 vccd1 _21614_/B sky130_fd_sc_hd__nand3_1
X_25381_ _26205_/CLK hold223/X vssd1 vssd1 vccd1 vccd1 hold221/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22593_ _25704_/Q _22592_/A _22592_/Y vssd1 vssd1 vccd1 vccd1 _22595_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24332_ hold1891/X _26176_/Q _24356_/S vssd1 vssd1 vccd1 vccd1 _24332_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21544_ _21595_/A _21547_/A vssd1 vssd1 vccd1 vccd1 _21545_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24263_ _24263_/A vssd1 vssd1 vccd1 vccd1 _26153_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21475_ _21475_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21475_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26002_ _26002_/CLK _26002_/D vssd1 vssd1 vccd1 vccd1 _26002_/Q sky130_fd_sc_hd__dfxtp_1
X_23214_ _12518_/Y _16980_/A _12533_/X input1/X vssd1 vssd1 vccd1 vccd1 _25907_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20426_ _20660_/A _20426_/B vssd1 vssd1 vccd1 vccd1 _20426_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24194_ hold899/X hold1831/X _24203_/S vssd1 vssd1 vccd1 vccd1 _24195_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23145_ _23145_/A _23193_/B _23145_/C vssd1 vssd1 vccd1 vccd1 _23145_/X sky130_fd_sc_hd__and3_1
X_20357_ _20357_/A vssd1 vssd1 vccd1 vccd1 _20358_/B sky130_fd_sc_hd__inv_2
XFILLER_0_30_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23076_ _23188_/A _23076_/B vssd1 vssd1 vccd1 vccd1 _23076_/X sky130_fd_sc_hd__or2_1
X_20288_ _25845_/Q _20288_/B _20288_/C vssd1 vssd1 vccd1 vccd1 _20291_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22027_ _18158_/B _17138_/B _18160_/A vssd1 vssd1 vccd1 vccd1 _22028_/B sky130_fd_sc_hd__o21ai_2
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2650 _15217_/X vssd1 vssd1 vccd1 vccd1 hold2650/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2661 _26277_/Q vssd1 vssd1 vccd1 vccd1 hold2661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2672 _15499_/X vssd1 vssd1 vccd1 vccd1 hold2672/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2683 _26234_/Q vssd1 vssd1 vccd1 vccd1 hold2683/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2694 _24808_/X vssd1 vssd1 vccd1 vccd1 _24809_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1960 _24731_/X vssd1 vssd1 vccd1 vccd1 _24732_/A sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ _13880_/A hold617/X vssd1 vssd1 vccd1 vccd1 hold618/A sky130_fd_sc_hd__nand2_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
X_14780_ _14786_/B _22036_/A vssd1 vssd1 vccd1 vccd1 _22035_/B sky130_fd_sc_hd__xnor2_2
Xhold1971 _12583_/Y vssd1 vssd1 vccd1 vccd1 _12584_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1982 _24962_/Y vssd1 vssd1 vccd1 vccd1 hold1982/X sky130_fd_sc_hd__dlygate4sd3_1
X_23978_ _23978_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23979_/A sky130_fd_sc_hd__and2_1
Xhold1993 _25960_/Q vssd1 vssd1 vccd1 vccd1 hold1993/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25717_ _26154_/CLK hold939/X vssd1 vssd1 vccd1 vccd1 hold937/A sky130_fd_sc_hd__dfxtp_1
X_13731_ _25752_/Q vssd1 vssd1 vccd1 vccd1 _18529_/B sky130_fd_sc_hd__inv_2
XFILLER_0_97_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22929_ _15524_/B _22680_/X _22829_/X vssd1 vssd1 vccd1 vccd1 _22929_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16450_ _16451_/A _16691_/B hold935/X vssd1 vssd1 vccd1 vccd1 _16452_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13662_ _13760_/A hold674/X vssd1 vssd1 vccd1 vccd1 hold675/A sky130_fd_sc_hd__nand2_1
X_25648_ _26152_/CLK _25648_/D vssd1 vssd1 vccd1 vccd1 _25648_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_39_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _16387_/A _16711_/A vssd1 vssd1 vccd1 vccd1 _16824_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12613_ _12613_/A _12613_/B vssd1 vssd1 vccd1 vccd1 _12613_/Y sky130_fd_sc_hd__nand2_1
X_16381_ _16489_/A vssd1 vssd1 vccd1 vccd1 _16382_/B sky130_fd_sc_hd__inv_2
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13593_ _25730_/Q vssd1 vssd1 vccd1 vccd1 _17957_/B sky130_fd_sc_hd__inv_2
XFILLER_0_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25579_ _26084_/CLK _25579_/D vssd1 vssd1 vccd1 vccd1 _25579_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18120_ _18122_/A _18122_/C vssd1 vssd1 vccd1 vccd1 _18121_/A sky130_fd_sc_hd__nand2_1
X_15332_ _16799_/B vssd1 vssd1 vccd1 vccd1 _22750_/B sky130_fd_sc_hd__inv_2
X_12544_ _23193_/B _15839_/B vssd1 vssd1 vccd1 vccd1 _14267_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_26_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18051_ _18529_/C vssd1 vssd1 vccd1 vccd1 _18891_/C sky130_fd_sc_hd__buf_8
X_15263_ _15263_/A _16768_/A vssd1 vssd1 vccd1 vccd1 _15264_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17002_ _17002_/A vssd1 vssd1 vccd1 vccd1 _19082_/A sky130_fd_sc_hd__buf_6
X_14214_ _18794_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14214_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_50_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15194_ _15621_/A _16221_/B vssd1 vssd1 vccd1 vccd1 _15197_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 _24858_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14145_ _25818_/Q vssd1 vssd1 vccd1 vccd1 _18572_/B sky130_fd_sc_hd__inv_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14076_ _14118_/A hold488/X vssd1 vssd1 vccd1 vccd1 hold489/A sky130_fd_sc_hd__nand2_1
X_18953_ _18953_/A _25837_/Q _18953_/C vssd1 vssd1 vccd1 vccd1 _20094_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_123_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17904_ _18611_/A _17908_/B vssd1 vssd1 vccd1 vccd1 _17906_/A sky130_fd_sc_hd__nand2_1
X_13027_ _17580_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13027_/X sky130_fd_sc_hd__or2_1
X_18884_ _18882_/Y _18883_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25688_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17835_ _20070_/A _17835_/B vssd1 vssd1 vccd1 vccd1 _19093_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17766_ _17767_/B _17766_/B vssd1 vssd1 vccd1 vccd1 _17768_/A sky130_fd_sc_hd__nand2b_1
X_14978_ _14976_/X hold1753/X _14928_/X vssd1 vssd1 vccd1 vccd1 _14978_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19505_ _21156_/A _21913_/B _25615_/Q vssd1 vssd1 vccd1 vccd1 _21160_/C sky130_fd_sc_hd__nand3_1
X_16717_ _16980_/A _16722_/B vssd1 vssd1 vccd1 vccd1 _16719_/B sky130_fd_sc_hd__nand2_1
X_13929_ _13941_/A _13929_/B vssd1 vssd1 vccd1 vccd1 _13929_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17697_ _17764_/B vssd1 vssd1 vccd1 vccd1 _17725_/B sky130_fd_sc_hd__inv_2
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19436_ _19434_/X _19435_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19436_/Y sky130_fd_sc_hd__a21oi_1
X_16648_ _16642_/B _16639_/Y _16631_/Y _16649_/A _16641_/B vssd1 vssd1 vccd1 vccd1
+ _16658_/B sky130_fd_sc_hd__o221a_1
XFILLER_0_186_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19367_ _19452_/A _19367_/B vssd1 vssd1 vccd1 vccd1 _19367_/Y sky130_fd_sc_hd__nand2_1
X_16579_ _16596_/A _16580_/A vssd1 vssd1 vccd1 vccd1 _16581_/A sky130_fd_sc_hd__or2_1
XFILLER_0_130_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18318_ _19488_/A vssd1 vssd1 vccd1 vccd1 _21878_/B sky130_fd_sc_hd__inv_2
X_19298_ _19296_/Y _19297_/Y _19086_/X vssd1 vssd1 vccd1 vccd1 _19298_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18249_ _18535_/A hold990/X _18393_/C vssd1 vssd1 vccd1 vccd1 _18249_/X sky130_fd_sc_hd__and3_1
XFILLER_0_72_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21260_ _21260_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21260_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold501 hold501/A vssd1 vssd1 vccd1 vccd1 hold501/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold512 hold512/A vssd1 vssd1 vccd1 vccd1 hold512/X sky130_fd_sc_hd__dlygate4sd3_1
X_20211_ _19177_/A _21924_/A _25587_/Q vssd1 vssd1 vccd1 vccd1 _20214_/A sky130_fd_sc_hd__a21o_1
Xhold523 hold523/A vssd1 vssd1 vccd1 vccd1 hold523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 hold534/A vssd1 vssd1 vccd1 vccd1 hold534/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 hold545/A vssd1 vssd1 vccd1 vccd1 hold545/X sky130_fd_sc_hd__dlygate4sd3_1
X_21191_ _21191_/A _21191_/B vssd1 vssd1 vccd1 vccd1 _21643_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold556 hold556/A vssd1 vssd1 vccd1 vccd1 hold556/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold567 hold567/A vssd1 vssd1 vccd1 vccd1 hold567/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold578 hold578/A vssd1 vssd1 vccd1 vccd1 hold578/X sky130_fd_sc_hd__dlygate4sd3_1
X_20142_ _19137_/A _21855_/A _25585_/Q vssd1 vssd1 vccd1 vccd1 _20143_/B sky130_fd_sc_hd__a21o_1
Xhold589 hold589/A vssd1 vssd1 vccd1 vccd1 hold589/X sky130_fd_sc_hd__dlygate4sd3_1
X_24950_ _24950_/A _24950_/B vssd1 vssd1 vccd1 vccd1 _24950_/Y sky130_fd_sc_hd__nand2_1
X_20073_ _21692_/A _21385_/A vssd1 vssd1 vccd1 vccd1 _20075_/A sky130_fd_sc_hd__nand2_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1201 _25577_/Q vssd1 vssd1 vccd1 vccd1 _16963_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23901_ hold2048/X hold1963/X _23907_/S vssd1 vssd1 vccd1 vccd1 _23902_/A sky130_fd_sc_hd__mux2_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1212 _19696_/Y vssd1 vssd1 vccd1 vccd1 _25750_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1223 _25125_/Q vssd1 vssd1 vccd1 vccd1 _19054_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24881_ _24958_/B _24873_/Y _24875_/Y _24880_/X vssd1 vssd1 vccd1 vccd1 _24881_/X
+ sky130_fd_sc_hd__a31o_1
Xhold1234 _25738_/Q vssd1 vssd1 vccd1 vccd1 _19526_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1245 _19113_/Y vssd1 vssd1 vccd1 vccd1 _25710_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1256 _25022_/Q vssd1 vssd1 vccd1 vccd1 _17296_/B sky130_fd_sc_hd__dlygate4sd3_1
X_23832_ _23832_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23833_/A sky130_fd_sc_hd__and2_1
XFILLER_0_139_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1267 _20661_/Y vssd1 vssd1 vccd1 vccd1 _25790_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1278 _25579_/Q vssd1 vssd1 vccd1 vccd1 _16977_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1289 _13200_/X vssd1 vssd1 vccd1 vccd1 _25086_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23763_ _23763_/A vssd1 vssd1 vccd1 vccd1 _25992_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20975_ _21464_/C _21513_/C vssd1 vssd1 vccd1 vccd1 _20978_/A sky130_fd_sc_hd__nand2_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25502_ _25510_/CLK _25502_/D vssd1 vssd1 vccd1 vccd1 hold882/A sky130_fd_sc_hd__dfxtp_1
X_22714_ _22705_/Y _22713_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22714_/X sky130_fd_sc_hd__a21o_1
X_23694_ _23694_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23695_/A sky130_fd_sc_hd__and2_1
XFILLER_0_94_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25433_ _26002_/CLK _25433_/D vssd1 vssd1 vccd1 vccd1 _25433_/Q sky130_fd_sc_hd__dfxtp_1
X_22645_ _22645_/A _22645_/B vssd1 vssd1 vccd1 vccd1 _22646_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25364_ _26190_/CLK hold76/X vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__dfxtp_1
X_22576_ _22576_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _22576_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24315_ _24315_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24316_/A sky130_fd_sc_hd__and2_1
X_21527_ _21578_/A _21531_/A vssd1 vssd1 vccd1 vccd1 _21529_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25295_ _26249_/CLK hold355/X vssd1 vssd1 vccd1 vccd1 hold353/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24246_ hold2352/X hold2153/X _24279_/S vssd1 vssd1 vccd1 vccd1 _24247_/A sky130_fd_sc_hd__mux2_1
X_21458_ _21458_/A _21458_/B vssd1 vssd1 vccd1 vccd1 _21459_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20409_ _20409_/A _20409_/B _20409_/C vssd1 vssd1 vccd1 vccd1 _20410_/B sky130_fd_sc_hd__nand3_1
X_24177_ _24177_/A vssd1 vssd1 vccd1 vccd1 _26125_/D sky130_fd_sc_hd__clkbuf_1
Xoutput8 output8/A vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__buf_12
Xoutput10 _26341_/Q vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__buf_12
X_21389_ _21389_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21394_/A sky130_fd_sc_hd__nand2_1
X_23128_ _23127_/A _22849_/X _23127_/B vssd1 vssd1 vccd1 vccd1 _23129_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15950_ _15951_/B _15951_/A vssd1 vssd1 vccd1 vccd1 _15961_/B sky130_fd_sc_hd__or2_1
X_23059_ _23059_/A _23187_/B vssd1 vssd1 vccd1 vccd1 _23059_/Y sky130_fd_sc_hd__nand2_1
X_14901_ _14899_/Y _14900_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14901_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15881_ _15881_/A _15881_/B vssd1 vssd1 vccd1 vccd1 _15882_/B sky130_fd_sc_hd__nand2_1
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2480 _26072_/Q vssd1 vssd1 vccd1 vccd1 hold2480/X sky130_fd_sc_hd__dlygate4sd3_1
X_17620_ _18252_/A _17620_/B vssd1 vssd1 vccd1 vccd1 _17620_/Y sky130_fd_sc_hd__nand2_1
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14832_ _14830_/Y _14831_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14832_/Y sky130_fd_sc_hd__a21oi_1
Xhold2491 _26183_/Q vssd1 vssd1 vccd1 vccd1 hold2491/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1790 _22406_/Y vssd1 vssd1 vccd1 vccd1 _25860_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17551_ _17549_/X _17528_/X _17550_/X vssd1 vssd1 vccd1 vccd1 _17552_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_59_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14763_ _21967_/B _15778_/B vssd1 vssd1 vccd1 vccd1 _14764_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _16513_/B _16502_/B vssd1 vssd1 vccd1 vccd1 _16524_/A sky130_fd_sc_hd__nand2_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13714_ _18469_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13714_/Y sky130_fd_sc_hd__nor2_1
X_17482_ _17605_/A _17482_/B vssd1 vssd1 vccd1 vccd1 _17482_/Y sky130_fd_sc_hd__nand2_1
X_14694_ _14694_/A vssd1 vssd1 vccd1 vccd1 _22680_/A sky130_fd_sc_hd__buf_4
XFILLER_0_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19221_ _26220_/Q hold768/X vssd1 vssd1 vccd1 vccd1 _19221_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_67_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16433_ _16431_/X _16432_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 hold934/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13645_ _18243_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13645_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_160_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19152_ _19150_/Y hold606/X _19086_/X vssd1 vssd1 vccd1 vccd1 hold607/A sky130_fd_sc_hd__a21oi_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16364_ _16378_/A _16365_/A vssd1 vssd1 vccd1 vccd1 _16366_/A sky130_fd_sc_hd__or2_1
XFILLER_0_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13576_ _26230_/Q _13426_/X _13468_/X _13575_/Y vssd1 vssd1 vccd1 vccd1 _13577_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _20888_/B _21871_/A vssd1 vssd1 vccd1 vccd1 _20882_/A sky130_fd_sc_hd__nand2_2
X_15315_ _26016_/Q _25952_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15316_/A sky130_fd_sc_hd__mux2_1
X_12527_ _12527_/A vssd1 vssd1 vccd1 vccd1 _12535_/A sky130_fd_sc_hd__clkinv_4
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19083_ _19081_/X _18879_/X _19082_/X vssd1 vssd1 vccd1 vccd1 _19084_/A sky130_fd_sc_hd__a21o_1
X_16295_ _16295_/A _16295_/B vssd1 vssd1 vccd1 vccd1 _16296_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_48_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18034_ _18529_/A _18034_/B _18529_/C vssd1 vssd1 vccd1 vccd1 _18035_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_87_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15246_ _15247_/B _16761_/A vssd1 vssd1 vccd1 vccd1 _15248_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_23_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15177_ _16733_/A _15177_/B vssd1 vssd1 vccd1 vccd1 _15178_/B sky130_fd_sc_hd__and2_1
XFILLER_0_23_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14128_ _18510_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14128_/Y sky130_fd_sc_hd__nor2_1
X_19985_ _19980_/X _19984_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19985_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_185_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18936_ _18936_/A _18936_/B _18936_/C vssd1 vssd1 vccd1 vccd1 _22694_/A sky130_fd_sc_hd__nand3_2
X_14059_ _18288_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14059_/Y sky130_fd_sc_hd__nor2_1
X_18867_ _18867_/A _18867_/B vssd1 vssd1 vccd1 vccd1 _22614_/A sky130_fd_sc_hd__or2_1
XFILLER_0_118_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17818_ _19018_/A _17818_/B vssd1 vssd1 vccd1 vccd1 _17818_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_118_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18798_ _18798_/A _18798_/B vssd1 vssd1 vccd1 vccd1 _18798_/X sky130_fd_sc_hd__xor2_1
X_17749_ _17748_/Y _17708_/A _17719_/B vssd1 vssd1 vccd1 vccd1 _17750_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_134_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20760_ _20760_/A _20760_/B vssd1 vssd1 vccd1 vccd1 _21677_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_187_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19419_ _19435_/B _19509_/B vssd1 vssd1 vccd1 vccd1 _19421_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20691_ _20691_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20696_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_147_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22430_ _22586_/A vssd1 vssd1 vccd1 vccd1 _23197_/A sky130_fd_sc_hd__buf_6
XFILLER_0_57_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22361_ _22358_/X _22359_/Y _22900_/B vssd1 vssd1 vccd1 vccd1 _22361_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24100_ _24100_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24101_/A sky130_fd_sc_hd__and2_1
XFILLER_0_66_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21312_ _21636_/A _21312_/B _21311_/X vssd1 vssd1 vccd1 vccd1 _21313_/B sky130_fd_sc_hd__or3b_1
X_25080_ _26164_/CLK _25080_/D vssd1 vssd1 vccd1 vccd1 _25080_/Q sky130_fd_sc_hd__dfxtp_1
X_22292_ _22653_/A _22292_/B vssd1 vssd1 vccd1 vccd1 _22292_/X sky130_fd_sc_hd__or2_1
XFILLER_0_143_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24031_ _24031_/A vssd1 vssd1 vccd1 vccd1 _26078_/D sky130_fd_sc_hd__clkbuf_1
Xhold320 hold320/A vssd1 vssd1 vccd1 vccd1 hold320/X sky130_fd_sc_hd__dlygate4sd3_1
X_21243_ _21243_/A _21243_/B vssd1 vssd1 vccd1 vccd1 _21245_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_130_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold331 hold331/A vssd1 vssd1 vccd1 vccd1 hold331/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 hold342/A vssd1 vssd1 vccd1 vccd1 hold342/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 hold353/A vssd1 vssd1 vccd1 vccd1 hold353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 hold364/A vssd1 vssd1 vccd1 vccd1 hold364/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 hold375/A vssd1 vssd1 vccd1 vccd1 hold375/X sky130_fd_sc_hd__dlygate4sd3_1
X_21174_ _21174_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _21179_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold386 hold386/A vssd1 vssd1 vccd1 vccd1 hold386/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 hold397/A vssd1 vssd1 vccd1 vccd1 hold397/X sky130_fd_sc_hd__dlygate4sd3_1
X_20125_ _20124_/Y _21228_/A _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20125_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25982_ _26004_/CLK _25982_/D vssd1 vssd1 vccd1 vccd1 _25982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24933_ hold889/A hold999/A _24942_/S vssd1 vssd1 vccd1 vccd1 _24934_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_176_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20056_ _20058_/B _20058_/C vssd1 vssd1 vccd1 vccd1 _20057_/A sky130_fd_sc_hd__nand2_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1020 _12913_/X vssd1 vssd1 vccd1 vccd1 _25033_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 _25732_/Q vssd1 vssd1 vccd1 vccd1 _19438_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1042 _12823_/X vssd1 vssd1 vccd1 vccd1 _25016_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1053 _25004_/Q vssd1 vssd1 vccd1 vccd1 _17045_/B sky130_fd_sc_hd__dlygate4sd3_1
X_24864_ _24864_/A _24944_/S vssd1 vssd1 vccd1 vccd1 _24864_/Y sky130_fd_sc_hd__nand2_1
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1064 _12929_/X vssd1 vssd1 vccd1 vccd1 _25036_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1075 _25740_/Q vssd1 vssd1 vccd1 vccd1 _19554_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 _16873_/Y vssd1 vssd1 vccd1 vccd1 _25564_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23815_ hold1943/X _26010_/Q _23831_/S vssd1 vssd1 vccd1 vccd1 _23815_/X sky130_fd_sc_hd__mux2_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 _25042_/Q vssd1 vssd1 vccd1 vccd1 _17486_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24795_ _24795_/A vssd1 vssd1 vccd1 vccd1 _26326_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23746_ _23746_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23747_/A sky130_fd_sc_hd__and2_1
X_20958_ _20956_/Y _20192_/X _19236_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _20958_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23677_ hold2071/X hold1903/X _23677_/S vssd1 vssd1 vccd1 vccd1 _23678_/A sky130_fd_sc_hd__mux2_1
X_20889_ _20888_/B _20889_/B _20889_/C vssd1 vssd1 vccd1 vccd1 _20890_/B sky130_fd_sc_hd__nand3b_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25416_ _25425_/CLK _25416_/D vssd1 vssd1 vccd1 vccd1 _25416_/Q sky130_fd_sc_hd__dfxtp_1
X_13430_ _26206_/Q _13426_/X _13429_/X vssd1 vssd1 vccd1 vccd1 _13430_/X sky130_fd_sc_hd__a21o_1
X_22628_ _22653_/A _22628_/B vssd1 vssd1 vccd1 vccd1 _22628_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13361_ _13220_/X _14635_/A _13242_/X _19687_/A vssd1 vssd1 vccd1 vccd1 _13361_/X
+ sky130_fd_sc_hd__a22o_1
X_22559_ _22559_/A _22900_/B vssd1 vssd1 vccd1 vccd1 _22559_/Y sky130_fd_sc_hd__nand2_1
X_25347_ _26299_/CLK hold214/X vssd1 vssd1 vccd1 vccd1 hold212/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15100_ _15100_/A _15100_/B vssd1 vssd1 vccd1 vccd1 _15101_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_133_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16080_ _16081_/B _16081_/A vssd1 vssd1 vccd1 vccd1 _16097_/B sky130_fd_sc_hd__or2_2
XFILLER_0_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13292_ _26184_/Q _13239_/X _13291_/X vssd1 vssd1 vccd1 vccd1 _13292_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_107_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25278_ _26232_/CLK hold118/X vssd1 vssd1 vccd1 vccd1 hold116/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15031_ _15031_/A vssd1 vssd1 vccd1 vccd1 _15032_/A sky130_fd_sc_hd__inv_2
X_24229_ _24229_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24230_/A sky130_fd_sc_hd__and2_1
XFILLER_0_47_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19770_ _26259_/Q _19134_/X hold500/X vssd1 vssd1 vccd1 vccd1 _19770_/Y sky130_fd_sc_hd__a21oi_1
X_16982_ _16980_/Y _15816_/A _16981_/Y vssd1 vssd1 vccd1 vccd1 _16982_/Y sky130_fd_sc_hd__o21ai_1
X_18721_ _18721_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18721_/Y sky130_fd_sc_hd__nand2_1
X_15933_ _15933_/A _15933_/B vssd1 vssd1 vccd1 vccd1 _15940_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18652_ _18793_/A _18652_/B _18894_/C vssd1 vssd1 vccd1 vccd1 _18653_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_189_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ _21796_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _15866_/A sky130_fd_sc_hd__nand2_1
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17603_ _17601_/X _17528_/X _17602_/X vssd1 vssd1 vccd1 vccd1 _17604_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_99_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14815_ _15839_/A _25994_/Q vssd1 vssd1 vccd1 vccd1 _22145_/A sky130_fd_sc_hd__nand2_1
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18583_ _22267_/B _25627_/Q vssd1 vssd1 vccd1 vccd1 _18585_/A sky130_fd_sc_hd__nand2_1
X_15795_ _15795_/A _16676_/B vssd1 vssd1 vccd1 vccd1 _15798_/A sky130_fd_sc_hd__nor2_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17534_ _17534_/A _17585_/A vssd1 vssd1 vccd1 vccd1 _17535_/B sky130_fd_sc_hd__xnor2_1
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _14746_/A vssd1 vssd1 vccd1 vccd1 _14938_/A sky130_fd_sc_hd__inv_2
XFILLER_0_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17465_ _17463_/X _17241_/X _17464_/X vssd1 vssd1 vccd1 vccd1 _17466_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_74_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14677_ _14675_/Y hold231/X _14646_/X vssd1 vssd1 vccd1 vccd1 hold232/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19204_ _26219_/Q _19134_/X hold739/X vssd1 vssd1 vccd1 vccd1 _19205_/C sky130_fd_sc_hd__a21o_1
X_16416_ _16416_/A _16416_/B vssd1 vssd1 vccd1 vccd1 _16440_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13628_ _13703_/A _13628_/B vssd1 vssd1 vccd1 vccd1 _13628_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_172_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17396_ _17467_/A _17396_/B vssd1 vssd1 vccd1 vccd1 _17396_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19135_ _26215_/Q _19134_/X hold715/A vssd1 vssd1 vccd1 vccd1 _19136_/C sky130_fd_sc_hd__a21o_1
X_16347_ _16347_/A _16347_/B vssd1 vssd1 vccd1 vccd1 _16361_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_137_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13559_ _14345_/A vssd1 vssd1 vccd1 vccd1 _13559_/X sky130_fd_sc_hd__buf_6
XFILLER_0_70_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19066_ _19066_/A _19066_/B vssd1 vssd1 vccd1 vccd1 _19067_/B sky130_fd_sc_hd__xnor2_1
X_16278_ _16059_/X _16273_/A _16277_/Y vssd1 vssd1 vccd1 vccd1 _16279_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18017_ _18017_/A _18017_/B _20214_/B vssd1 vssd1 vccd1 vccd1 _18024_/A sky130_fd_sc_hd__and3_2
X_15229_ hold885/X vssd1 vssd1 vccd1 vccd1 _15231_/A sky130_fd_sc_hd__inv_2
XFILLER_0_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19968_ _26274_/Q _19134_/X hold680/X vssd1 vssd1 vccd1 vccd1 _19969_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18919_ _18919_/A _18919_/B vssd1 vssd1 vccd1 vccd1 _18919_/X sky130_fd_sc_hd__xor2_1
X_19899_ _19970_/A _19914_/B vssd1 vssd1 vccd1 vccd1 _19901_/A sky130_fd_sc_hd__xnor2_1
X_21930_ _21902_/X _21929_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _21930_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_179_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21861_ _21833_/X _21860_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _21861_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_171_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23600_ _24970_/Q _24969_/Q _24971_/Q vssd1 vssd1 vccd1 vccd1 _23600_/X sky130_fd_sc_hd__a21o_1
X_20812_ _21042_/A _20812_/B _20811_/X vssd1 vssd1 vccd1 vccd1 _20813_/B sky130_fd_sc_hd__or3b_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21792_ _21762_/X _21790_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _21792_/Y sky130_fd_sc_hd__o21ai_1
X_24580_ _24580_/A vssd1 vssd1 vccd1 vccd1 _26256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20743_ _20743_/A _25857_/Q vssd1 vssd1 vccd1 vccd1 _20748_/B sky130_fd_sc_hd__nand2_1
X_23531_ _23519_/X _23530_/X _24949_/S vssd1 vssd1 vccd1 vccd1 _23531_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_147_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23462_ _24956_/S hold272/A _23461_/X vssd1 vssd1 vccd1 vccd1 _23462_/Y sky130_fd_sc_hd__o21ai_1
X_26250_ _26281_/CLK _26250_/D vssd1 vssd1 vccd1 vccd1 _26250_/Q sky130_fd_sc_hd__dfxtp_2
X_20674_ _20677_/A _20677_/C vssd1 vssd1 vccd1 vccd1 _20675_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_169_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22413_ _22413_/A _22413_/B vssd1 vssd1 vccd1 vccd1 _22414_/B sky130_fd_sc_hd__nand2_1
X_25201_ _25743_/CLK hold738/X vssd1 vssd1 vccd1 vccd1 hold736/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23393_ _24940_/S hold278/A _23392_/X vssd1 vssd1 vccd1 vccd1 _23393_/Y sky130_fd_sc_hd__o21ai_1
X_26181_ _26181_/CLK _26181_/D vssd1 vssd1 vccd1 vccd1 _26181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22344_ _22344_/A _22387_/B vssd1 vssd1 vccd1 vccd1 _22344_/Y sky130_fd_sc_hd__nand2_1
X_25132_ _25712_/CLK hold717/X vssd1 vssd1 vccd1 vccd1 hold715/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25063_ _26148_/CLK _25063_/D vssd1 vssd1 vccd1 vccd1 _25063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22275_ _22496_/A _22742_/B vssd1 vssd1 vccd1 vccd1 _22287_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24014_ hold2480/X hold2253/X _24047_/S vssd1 vssd1 vccd1 vccd1 _24015_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_131_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21226_ _21226_/A _21226_/B vssd1 vssd1 vccd1 vccd1 _21227_/A sky130_fd_sc_hd__nand2_1
Xhold150 hold150/A vssd1 vssd1 vccd1 vccd1 hold150/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold161 hold161/A vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 hold172/A vssd1 vssd1 vccd1 vccd1 hold172/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 hold183/A vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 hold194/A vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
X_21157_ _21157_/A _21157_/B vssd1 vssd1 vccd1 vccd1 _21160_/B sky130_fd_sc_hd__nand2_1
X_20108_ _21708_/A _21402_/A vssd1 vssd1 vccd1 vccd1 _20117_/A sky130_fd_sc_hd__nand2_1
X_25965_ _26032_/CLK _25965_/D vssd1 vssd1 vccd1 vccd1 _25965_/Q sky130_fd_sc_hd__dfxtp_1
X_21088_ _21580_/B _21529_/C vssd1 vssd1 vccd1 vccd1 _21089_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_176_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24916_ hold894/A hold933/A _24944_/S vssd1 vssd1 vccd1 vccd1 _24917_/B sky130_fd_sc_hd__mux2_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12930_ _14260_/A vssd1 vssd1 vccd1 vccd1 _12930_/X sky130_fd_sc_hd__clkbuf_8
X_20039_ _20039_/A _20039_/B vssd1 vssd1 vccd1 vccd1 _20040_/A sky130_fd_sc_hd__nand2_1
X_25896_ _26080_/CLK _25896_/D vssd1 vssd1 vccd1 vccd1 _25896_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24847_ _24845_/X _24846_/X _24858_/S vssd1 vssd1 vccd1 vccd1 _24847_/X sky130_fd_sc_hd__mux2_1
X_12861_ _26235_/Q _25604_/Q vssd1 vssd1 vccd1 vccd1 _14358_/A sky130_fd_sc_hd__xor2_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _14645_/A hold368/X vssd1 vssd1 vccd1 vccd1 hold369/A sky130_fd_sc_hd__nand2_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _25567_/Q vssd1 vssd1 vccd1 vccd1 _22982_/B sky130_fd_sc_hd__inv_2
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _12746_/X hold2/X _14910_/B _12791_/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__o211a_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24778_ hold2666/X hold2655/X _24817_/S vssd1 vssd1 vccd1 vccd1 _24779_/A sky130_fd_sc_hd__mux2_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14531_ _14585_/A hold227/X vssd1 vssd1 vccd1 vccd1 hold228/A sky130_fd_sc_hd__nand2_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23729_ _23729_/A vssd1 vssd1 vccd1 vccd1 _25981_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17250_ _19373_/A _17250_/B vssd1 vssd1 vccd1 vccd1 _17535_/A sky130_fd_sc_hd__xor2_4
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _14465_/A hold29/X vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__nand2_1
X_16201_ _16212_/A hold882/X vssd1 vssd1 vccd1 vccd1 _16201_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_181_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13413_ _13413_/A vssd1 vssd1 vccd1 vccd1 _19816_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_183_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17181_ _19303_/A _17181_/B vssd1 vssd1 vccd1 vccd1 _17499_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_3_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14393_ _14391_/Y hold48/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16132_ _16161_/A vssd1 vssd1 vccd1 vccd1 _16132_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_180_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13344_ _26192_/Q _13239_/X _13343_/X vssd1 vssd1 vccd1 vccd1 _13344_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16063_ _16063_/A _16697_/B _16071_/A vssd1 vssd1 vccd1 vccd1 _16063_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_161_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13275_ _18679_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13275_/X sky130_fd_sc_hd__or2_1
X_15014_ _15014_/A _15034_/A vssd1 vssd1 vccd1 vccd1 _15029_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_122_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19822_ _19820_/X _19821_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19822_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16965_ _22145_/B _16970_/B vssd1 vssd1 vccd1 vccd1 _16967_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19753_ _19751_/Y _19752_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19753_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15916_ _21933_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _15918_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_155_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18704_ _19758_/A vssd1 vssd1 vccd1 vccd1 _22408_/B sky130_fd_sc_hd__inv_2
X_19684_ _26253_/Q hold925/X vssd1 vssd1 vccd1 vccd1 _19684_/Y sky130_fd_sc_hd__nand2_1
X_16896_ _16897_/B _16897_/A vssd1 vssd1 vccd1 vccd1 _16896_/X sky130_fd_sc_hd__or2_1
XFILLER_0_188_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18635_ _18635_/A _20321_/A vssd1 vssd1 vccd1 vccd1 _18966_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15847_ _16660_/B vssd1 vssd1 vccd1 vccd1 _16686_/B sky130_fd_sc_hd__buf_8
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18566_ _25882_/Q _22236_/A vssd1 vssd1 vccd1 vccd1 _18574_/A sky130_fd_sc_hd__or2_2
X_15778_ _16665_/A _15778_/B vssd1 vssd1 vccd1 vccd1 _16967_/A sky130_fd_sc_hd__nand2_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17517_ _17605_/A _17517_/B vssd1 vssd1 vccd1 vccd1 _17517_/Y sky130_fd_sc_hd__nand2_1
X_14729_ _25841_/Q _13466_/A _14728_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14730_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18497_ _18497_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18497_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17448_ _17448_/A _17448_/B vssd1 vssd1 vccd1 vccd1 _17448_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_28_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17379_ _21211_/B _25873_/Q _25809_/Q vssd1 vssd1 vccd1 vccd1 _17380_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_160_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19118_ _20284_/A _18117_/C _20288_/C vssd1 vssd1 vccd1 vccd1 _19220_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_172_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20390_ _20390_/A _20390_/B vssd1 vssd1 vccd1 vccd1 _20394_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19049_ _19049_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _19049_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_112_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22060_ _22653_/A _22060_/B vssd1 vssd1 vccd1 vccd1 _22060_/X sky130_fd_sc_hd__or2_1
XFILLER_0_112_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21011_ _21011_/A _21011_/B vssd1 vssd1 vccd1 vccd1 _21012_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25750_ _25750_/CLK _25750_/D vssd1 vssd1 vccd1 vccd1 _25750_/Q sky130_fd_sc_hd__dfxtp_1
X_22962_ _23188_/A _22962_/B vssd1 vssd1 vccd1 vccd1 _22962_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24701_ hold2602/X _26296_/Q _24740_/S vssd1 vssd1 vccd1 vccd1 _24701_/X sky130_fd_sc_hd__mux2_1
X_21913_ _25807_/Q _21913_/B vssd1 vssd1 vccd1 vccd1 _21913_/Y sky130_fd_sc_hd__nor2_1
X_25681_ _26313_/CLK _25681_/D vssd1 vssd1 vccd1 vccd1 _25681_/Q sky130_fd_sc_hd__dfxtp_1
X_22893_ _22893_/A _22893_/B vssd1 vssd1 vccd1 vccd1 _22893_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24632_ _24632_/A vssd1 vssd1 vccd1 vccd1 _26273_/D sky130_fd_sc_hd__clkbuf_1
X_21844_ _21844_/A _21844_/B vssd1 vssd1 vccd1 vccd1 _21844_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_167_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21775_ _21775_/A _21775_/B vssd1 vssd1 vccd1 vccd1 _21775_/Y sky130_fd_sc_hd__nand2_1
X_24563_ hold2582/X _26251_/Q _24587_/S vssd1 vssd1 vccd1 vccd1 _24563_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26302_ _26302_/CLK _26302_/D vssd1 vssd1 vccd1 vccd1 _26302_/Q sky130_fd_sc_hd__dfxtp_2
X_23514_ hold71/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23514_/X sky130_fd_sc_hd__or2b_1
X_20726_ _21384_/C _21660_/B vssd1 vssd1 vccd1 vccd1 _20728_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_148_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24494_ _24494_/A vssd1 vssd1 vccd1 vccd1 _26228_/D sky130_fd_sc_hd__clkbuf_1
X_26233_ _26235_/CLK _26233_/D vssd1 vssd1 vccd1 vccd1 _26233_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_162_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20657_ _21042_/A _20657_/B _20656_/X vssd1 vssd1 vccd1 vccd1 _20658_/B sky130_fd_sc_hd__or3b_1
X_23445_ _23439_/X _23444_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _23445_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23376_ _23376_/A _23376_/B vssd1 vssd1 vccd1 vccd1 _23380_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26164_ _26164_/CLK _26164_/D vssd1 vssd1 vccd1 vccd1 _26164_/Q sky130_fd_sc_hd__dfxtp_1
X_20588_ _20588_/A _25853_/Q vssd1 vssd1 vccd1 vccd1 _20593_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25115_ _26198_/CLK _25115_/D vssd1 vssd1 vccd1 vccd1 _25115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22327_ _25821_/Q _22327_/B vssd1 vssd1 vccd1 vccd1 _22327_/Y sky130_fd_sc_hd__nor2_1
X_26095_ _26096_/CLK _26095_/D vssd1 vssd1 vccd1 vccd1 _26095_/Q sky130_fd_sc_hd__dfxtp_1
X_13060_ _26273_/Q _25642_/Q vssd1 vssd1 vccd1 vccd1 _14479_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_131_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22258_ _22256_/X _22257_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _22258_/Y sky130_fd_sc_hd__a21oi_2
X_25046_ _26130_/CLK _25046_/D vssd1 vssd1 vccd1 vccd1 _25046_/Q sky130_fd_sc_hd__dfxtp_1
X_21209_ _21207_/Y _21208_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21209_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22189_ _22189_/A _25852_/Q vssd1 vssd1 vccd1 vccd1 _22189_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16750_ _16858_/A _16750_/B vssd1 vssd1 vccd1 vccd1 _16750_/Y sky130_fd_sc_hd__nand2_1
X_25948_ _26014_/CLK _25948_/D vssd1 vssd1 vccd1 vccd1 _25948_/Q sky130_fd_sc_hd__dfxtp_1
X_13962_ _14000_/A hold853/X vssd1 vssd1 vccd1 vccd1 _13962_/Y sky130_fd_sc_hd__nand2_1
X_15701_ _15701_/A _15718_/A vssd1 vssd1 vccd1 vccd1 _15701_/Y sky130_fd_sc_hd__nand2_1
X_12913_ _12840_/X _12911_/X _12827_/X _12912_/X vssd1 vssd1 vccd1 vccd1 _12913_/X
+ sky130_fd_sc_hd__o211a_1
X_16681_ _16681_/A _16681_/B vssd1 vssd1 vccd1 vccd1 _16683_/A sky130_fd_sc_hd__nand2_1
X_25879_ _25901_/CLK _25879_/D vssd1 vssd1 vccd1 vccd1 _25879_/Q sky130_fd_sc_hd__dfxtp_2
X_13893_ _13888_/Y _13892_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold852/A sky130_fd_sc_hd__a21oi_1
X_18420_ _19560_/A vssd1 vssd1 vccd1 vccd1 _22040_/B sky130_fd_sc_hd__inv_2
X_15632_ _16914_/B vssd1 vssd1 vccd1 vccd1 _23031_/B sky130_fd_sc_hd__inv_2
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _17269_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12844_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18351_ _18555_/A _18698_/A vssd1 vssd1 vccd1 vccd1 _18352_/B sky130_fd_sc_hd__xnor2_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _25566_/Q vssd1 vssd1 vccd1 vccd1 _22965_/B sky130_fd_sc_hd__inv_2
XFILLER_0_115_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12775_ hold992/X _12748_/X _12774_/X vssd1 vssd1 vccd1 vccd1 hold993/A sky130_fd_sc_hd__a21o_1
XFILLER_0_16_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _21022_/B _25866_/Q _21045_/B vssd1 vssd1 vccd1 vccd1 _17303_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _14512_/Y hold126/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold127/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ _18446_/A _19554_/B _21716_/A vssd1 vssd1 vccd1 vccd1 _18283_/C sky130_fd_sc_hd__nand3_1
X_15494_ _15495_/B _16855_/A vssd1 vssd1 vccd1 vccd1 _15496_/A sky130_fd_sc_hd__nor2_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17233_ _20883_/B _25861_/Q _25797_/Q vssd1 vssd1 vccd1 vccd1 _17234_/B sky130_fd_sc_hd__mux2_2
X_14445_ _14443_/Y hold18/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_181_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17164_ _17272_/A _17164_/B vssd1 vssd1 vccd1 vccd1 _17164_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14376_ _14376_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14376_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_135_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16115_ _16133_/A _16133_/B _16134_/A vssd1 vssd1 vccd1 vccd1 _16125_/A sky130_fd_sc_hd__a21o_1
Xhold908 hold908/A vssd1 vssd1 vccd1 vccd1 hold908/X sky130_fd_sc_hd__buf_1
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13327_ _18839_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13327_/X sky130_fd_sc_hd__or2_1
Xhold919 hold919/A vssd1 vssd1 vccd1 vccd1 hold919/X sky130_fd_sc_hd__dlygate4sd3_1
X_17095_ _17095_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17095_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16046_ hold800/X vssd1 vssd1 vccd1 vccd1 _16049_/B sky130_fd_sc_hd__inv_2
XFILLER_0_177_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13258_ _13207_/X _13256_/X _13192_/X _13257_/X vssd1 vssd1 vccd1 vccd1 _13258_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13189_ _26296_/Q _19303_/A vssd1 vssd1 vccd1 vccd1 _14551_/A sky130_fd_sc_hd__xor2_1
Xhold2309 _26159_/Q vssd1 vssd1 vccd1 vccd1 hold2309/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_23_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19805_ _19821_/B _19888_/B vssd1 vssd1 vccd1 vccd1 _19807_/A sky130_fd_sc_hd__xnor2_1
X_17997_ _25859_/Q _21800_/A vssd1 vssd1 vccd1 vccd1 _18005_/A sky130_fd_sc_hd__or2_2
Xhold1608 _25619_/Q vssd1 vssd1 vccd1 vccd1 _17467_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1619 _21510_/Y vssd1 vssd1 vccd1 vccd1 _25824_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16948_ _16948_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16948_/Y sky130_fd_sc_hd__nand2_1
X_19736_ _19728_/X _19735_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19736_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_189_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16879_ _16977_/A _16879_/B vssd1 vssd1 vccd1 vccd1 _16879_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19667_ _19723_/A _19667_/B vssd1 vssd1 vccd1 vccd1 _19667_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_189_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18618_ _19026_/A _18618_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18618_/X sky130_fd_sc_hd__and3_1
XFILLER_0_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19598_ _26247_/Q _19483_/X hold614/X vssd1 vssd1 vccd1 vccd1 _19598_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18549_ _18611_/A _25753_/Q vssd1 vssd1 vccd1 vccd1 _18551_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21560_ _21611_/A _21563_/A vssd1 vssd1 vccd1 vccd1 _21561_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_185_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20511_ _20511_/A _22165_/B _20511_/C vssd1 vssd1 vccd1 vccd1 _20514_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_90_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21491_ _21491_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21491_/Y sky130_fd_sc_hd__nand2_1
X_23230_ _23232_/A vssd1 vssd1 vccd1 vccd1 _24867_/S sky130_fd_sc_hd__inv_8
XFILLER_0_172_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20442_ _22988_/B vssd1 vssd1 vccd1 vccd1 _22396_/B sky130_fd_sc_hd__inv_2
XFILLER_0_27_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23161_ _23161_/A _23193_/B _23161_/C vssd1 vssd1 vccd1 vccd1 _23161_/X sky130_fd_sc_hd__and3_1
XFILLER_0_28_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20373_ _21515_/A vssd1 vssd1 vccd1 vccd1 _21514_/A sky130_fd_sc_hd__inv_4
XFILLER_0_141_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22112_ _22093_/X _22111_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _22112_/Y sky130_fd_sc_hd__o21ai_1
X_23092_ _23188_/A _23092_/B vssd1 vssd1 vccd1 vccd1 _23092_/X sky130_fd_sc_hd__or2_1
XFILLER_0_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_208_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _26112_/CLK sky130_fd_sc_hd__clkbuf_16
X_22043_ _19560_/A _22042_/A _22042_/Y vssd1 vssd1 vccd1 vccd1 _22045_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_167_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25802_ _25802_/CLK _25802_/D vssd1 vssd1 vccd1 vccd1 _25802_/Q sky130_fd_sc_hd__dfxtp_1
X_23994_ _23994_/A vssd1 vssd1 vccd1 vccd1 _26066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25733_ _26286_/CLK _25733_/D vssd1 vssd1 vccd1 vccd1 _25733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22945_ _23188_/A _22945_/B vssd1 vssd1 vccd1 vccd1 _22945_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25664_ _26297_/CLK _25664_/D vssd1 vssd1 vccd1 vccd1 _25664_/Q sky130_fd_sc_hd__dfxtp_1
X_22876_ _22876_/A _22876_/B vssd1 vssd1 vccd1 vccd1 _22877_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_168_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24615_ hold2586/X _26268_/Q _24664_/S vssd1 vssd1 vccd1 vccd1 _24615_/X sky130_fd_sc_hd__mux2_1
X_21827_ _21799_/X _21826_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _21827_/Y sky130_fd_sc_hd__o21ai_1
X_25595_ _25596_/CLK _25595_/D vssd1 vssd1 vccd1 vccd1 _25595_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12560_ _12560_/A _24836_/B _12564_/A vssd1 vssd1 vccd1 vccd1 _12561_/A sky130_fd_sc_hd__and3_1
X_24546_ _24546_/A vssd1 vssd1 vccd1 vccd1 _26245_/D sky130_fd_sc_hd__clkbuf_1
X_21758_ _21756_/Y _21757_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21758_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20709_ _20709_/A _20709_/B vssd1 vssd1 vccd1 vccd1 _21387_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_47_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12491_ _12491_/A vssd1 vssd1 vccd1 vccd1 _23193_/B sky130_fd_sc_hd__buf_8
X_24477_ hold2723/X hold2617/X _24510_/S vssd1 vssd1 vccd1 vccd1 _24478_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21689_ _21692_/B _21693_/A vssd1 vssd1 vccd1 vccd1 _21691_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_163_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14230_ _14236_/A hold383/X vssd1 vssd1 vccd1 vccd1 hold384/A sky130_fd_sc_hd__nand2_1
X_26216_ _26216_/CLK _26216_/D vssd1 vssd1 vccd1 vccd1 _26216_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_124_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23428_ _24940_/S hold218/A _23427_/X vssd1 vssd1 vccd1 vccd1 _23428_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26147_ _26148_/CLK _26147_/D vssd1 vssd1 vccd1 vccd1 _26147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14161_ _14180_/A _14161_/B vssd1 vssd1 vccd1 vccd1 _14161_/Y sky130_fd_sc_hd__nand2_1
X_23359_ _23360_/B _23360_/A vssd1 vssd1 vccd1 vccd1 _23359_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13112_ _26154_/Q _13065_/X _13111_/X vssd1 vssd1 vccd1 vccd1 _13112_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_132_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26078_ _26079_/CLK _26078_/D vssd1 vssd1 vccd1 vccd1 _26078_/Q sky130_fd_sc_hd__dfxtp_1
X_14092_ _14180_/A _14092_/B vssd1 vssd1 vccd1 vccd1 _14092_/Y sky130_fd_sc_hd__nand2_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25029_ _26112_/CLK _25029_/D vssd1 vssd1 vccd1 vccd1 _25029_/Q sky130_fd_sc_hd__dfxtp_1
X_13043_ _13018_/X _13041_/X _13005_/X _13042_/X vssd1 vssd1 vccd1 vccd1 _13043_/X
+ sky130_fd_sc_hd__o211a_1
X_17920_ _25649_/Q vssd1 vssd1 vccd1 vccd1 _21855_/A sky130_fd_sc_hd__inv_2
XFILLER_0_79_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17851_ _25657_/Q vssd1 vssd1 vccd1 vccd1 _22106_/A sky130_fd_sc_hd__inv_2
X_16802_ _16803_/B _16803_/A vssd1 vssd1 vccd1 vccd1 _16802_/X sky130_fd_sc_hd__or2_1
X_17782_ _17738_/A _17740_/B _17771_/C vssd1 vssd1 vccd1 vccd1 _17783_/B sky130_fd_sc_hd__o21ai_1
X_14994_ _14992_/X hold2247/X _14928_/X vssd1 vssd1 vccd1 vccd1 _14994_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16733_ _16733_/A _16733_/B vssd1 vssd1 vccd1 vccd1 _16733_/Y sky130_fd_sc_hd__nand2_1
X_19521_ _19537_/B _19607_/B vssd1 vssd1 vccd1 vccd1 _19523_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13945_ _25786_/Q vssd1 vssd1 vccd1 vccd1 _17896_/B sky130_fd_sc_hd__inv_2
XFILLER_0_152_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19452_ _19452_/A _19452_/B vssd1 vssd1 vccd1 vccd1 _19452_/Y sky130_fd_sc_hd__nand2_1
X_16664_ hold689/X vssd1 vssd1 vccd1 vccd1 _16667_/B sky130_fd_sc_hd__inv_2
XFILLER_0_159_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13876_ _17834_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13876_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_69_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15615_ _15560_/A _15694_/A _15695_/A vssd1 vssd1 vccd1 vccd1 _15615_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_158_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18403_ _18445_/A _18408_/B vssd1 vssd1 vccd1 vccd1 _18405_/A sky130_fd_sc_hd__nand2_1
X_19383_ _19380_/Y _19381_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19383_/Y sky130_fd_sc_hd__a21oi_1
X_12827_ _23377_/B vssd1 vssd1 vccd1 vccd1 _12827_/X sky130_fd_sc_hd__buf_4
XFILLER_0_57_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16595_ _16592_/Y _16593_/Y _16594_/X vssd1 vssd1 vccd1 vccd1 hold963/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_189_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18334_ _18332_/X _18269_/X _18333_/X vssd1 vssd1 vccd1 vccd1 _18335_/A sky130_fd_sc_hd__a21o_1
X_15546_ _15546_/A _15546_/B vssd1 vssd1 vccd1 vccd1 _15547_/A sky130_fd_sc_hd__nand2_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12758_ _26215_/Q _25584_/Q vssd1 vssd1 vccd1 vccd1 _14295_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_189_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18265_ _21053_/B _21775_/A vssd1 vssd1 vccd1 vccd1 _21047_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_189_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15477_ hold916/X _15479_/A vssd1 vssd1 vccd1 vccd1 _15481_/A sky130_fd_sc_hd__nor2_1
X_12689_ _12689_/A vssd1 vssd1 vccd1 vccd1 _12713_/B sky130_fd_sc_hd__inv_2
XFILLER_0_154_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17216_ _17216_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17216_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_142_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14428_ _14428_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14428_/Y sky130_fd_sc_hd__nand2_1
X_18196_ _18196_/A _18196_/B vssd1 vssd1 vccd1 vccd1 _21971_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_170_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17147_ _17423_/A _17147_/B vssd1 vssd1 vccd1 vccd1 _17147_/X sky130_fd_sc_hd__xor2_1
Xhold705 hold705/A vssd1 vssd1 vccd1 vccd1 hold705/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14359_ _14404_/A hold362/X vssd1 vssd1 vccd1 vccd1 hold363/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold716 hold716/A vssd1 vssd1 vccd1 vccd1 hold716/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold727 hold727/A vssd1 vssd1 vccd1 vccd1 hold727/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold738 hold738/A vssd1 vssd1 vccd1 vccd1 hold738/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17078_ _17076_/X _23187_/B _17077_/X vssd1 vssd1 vccd1 vccd1 _17079_/A sky130_fd_sc_hd__a21o_1
Xhold749 hold749/A vssd1 vssd1 vccd1 vccd1 hold749/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16029_ _16006_/A _16053_/A _16028_/Y vssd1 vssd1 vccd1 vccd1 _16031_/A sky130_fd_sc_hd__a21o_1
Xhold2106 _24990_/Q vssd1 vssd1 vccd1 vccd1 _12689_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2117 _15081_/Y vssd1 vssd1 vccd1 vccd1 _25433_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2128 _25973_/Q vssd1 vssd1 vccd1 vccd1 hold2128/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2139 _23279_/X vssd1 vssd1 vccd1 vccd1 _23280_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1405 _25111_/Q vssd1 vssd1 vccd1 vccd1 _18941_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 _19269_/Y vssd1 vssd1 vccd1 vccd1 _25720_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1427 _25553_/Q vssd1 vssd1 vccd1 vccd1 _16799_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1438 _16835_/Y vssd1 vssd1 vccd1 vccd1 _25558_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1449 _25402_/Q vssd1 vssd1 vccd1 vccd1 _14822_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19719_ _19720_/B _19720_/A vssd1 vssd1 vccd1 vccd1 _19719_/X sky130_fd_sc_hd__or2_1
X_20991_ _21235_/A _20991_/B vssd1 vssd1 vccd1 vccd1 _20991_/Y sky130_fd_sc_hd__nand2_1
X_22730_ _22730_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22730_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22661_ _22652_/Y _22660_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22661_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_48_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24400_ hold2363/X hold2310/X _24433_/S vssd1 vssd1 vccd1 vccd1 _24401_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21612_ _21612_/A _21661_/B vssd1 vssd1 vccd1 vccd1 _21613_/C sky130_fd_sc_hd__nand2_1
X_25380_ _25418_/CLK hold40/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dfxtp_1
X_22592_ _22592_/A _22592_/B vssd1 vssd1 vccd1 vccd1 _22592_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_168_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24331_ _24331_/A vssd1 vssd1 vccd1 vccd1 _26175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21543_ _21546_/A _21596_/A vssd1 vssd1 vccd1 vccd1 _21545_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_145_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24262_ _24262_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24263_/A sky130_fd_sc_hd__and2_1
XFILLER_0_90_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21474_ _21474_/A _21474_/B vssd1 vssd1 vccd1 vccd1 _21475_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26001_ _26001_/CLK _26001_/D vssd1 vssd1 vccd1 vccd1 _26001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23213_ _23213_/A vssd1 vssd1 vccd1 vccd1 _25906_/D sky130_fd_sc_hd__inv_2
XFILLER_0_16_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20425_ _20425_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _20425_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_114_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24193_ _24193_/A vssd1 vssd1 vccd1 vccd1 _26130_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23144_ _23143_/A _22849_/X _23143_/B vssd1 vssd1 vccd1 vccd1 _23145_/C sky130_fd_sc_hd__o21ai_1
X_20356_ _20356_/A _20357_/A vssd1 vssd1 vccd1 vccd1 _20359_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_144_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23075_ _23075_/A _23187_/B vssd1 vssd1 vccd1 vccd1 _23075_/Y sky130_fd_sc_hd__nand2_1
X_20287_ _20287_/A _25845_/Q vssd1 vssd1 vccd1 vccd1 _20291_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_105_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22026_ _22026_/A _22026_/B vssd1 vssd1 vccd1 vccd1 _22028_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_179_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2640 _24566_/X vssd1 vssd1 vccd1 vccd1 _24567_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2651 _15219_/Y vssd1 vssd1 vccd1 vccd1 _25441_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2662 _24645_/X vssd1 vssd1 vccd1 vccd1 _24646_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2673 _15501_/Y vssd1 vssd1 vccd1 vccd1 _25457_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2684 _26332_/Q vssd1 vssd1 vccd1 vccd1 hold2684/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2695 _26333_/Q vssd1 vssd1 vccd1 vccd1 hold2695/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1950 _24293_/X vssd1 vssd1 vccd1 vccd1 _24294_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1961 _26139_/Q vssd1 vssd1 vccd1 vccd1 hold1961/X sky130_fd_sc_hd__dlygate4sd3_1
X_23977_ _26060_/Q hold2422/X _24001_/S vssd1 vssd1 vccd1 vccd1 _23977_/X sky130_fd_sc_hd__mux2_1
Xhold1972 _26112_/Q vssd1 vssd1 vccd1 vccd1 hold1972/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1983 _24963_/X vssd1 vssd1 vccd1 vccd1 _26341_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1994 _23665_/X vssd1 vssd1 vccd1 vccd1 _23666_/A sky130_fd_sc_hd__dlygate4sd3_1
X_25716_ _25716_/CLK _25716_/D vssd1 vssd1 vccd1 vccd1 _25716_/Q sky130_fd_sc_hd__dfxtp_1
X_13730_ _13760_/A hold380/X vssd1 vssd1 vccd1 vccd1 hold381/A sky130_fd_sc_hd__nand2_1
XFILLER_0_98_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22928_ _23188_/A _22928_/B vssd1 vssd1 vccd1 vccd1 _22928_/X sky130_fd_sc_hd__or2_1
XFILLER_0_58_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13661_ hold630/X _13660_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold631/A sky130_fd_sc_hd__a21oi_1
X_25647_ _25712_/CLK _25647_/D vssd1 vssd1 vccd1 vccd1 _25647_/Q sky130_fd_sc_hd__dfxtp_2
X_22859_ _22859_/A _23168_/B vssd1 vssd1 vccd1 vccd1 _22860_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_116_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15400_ _15400_/A vssd1 vssd1 vccd1 vccd1 _16387_/A sky130_fd_sc_hd__inv_2
XFILLER_0_13_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _12613_/B _12613_/A vssd1 vssd1 vccd1 vccd1 _12614_/A sky130_fd_sc_hd__or2_1
X_16380_ _16380_/A _16380_/B vssd1 vssd1 vccd1 vccd1 _16489_/A sky130_fd_sc_hd__nand2_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25578_ _26084_/CLK _25578_/D vssd1 vssd1 vccd1 vccd1 _25578_/Q sky130_fd_sc_hd__dfxtp_1
X_13592_ _13642_/A hold455/X vssd1 vssd1 vccd1 vccd1 hold456/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15331_ _15827_/A _15407_/B _15408_/A vssd1 vssd1 vccd1 vccd1 _15331_/X sky130_fd_sc_hd__a21o_1
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12543_ _17685_/A vssd1 vssd1 vccd1 vccd1 _17707_/B sky130_fd_sc_hd__inv_2
X_24529_ hold2557/X _26240_/Q _24587_/S vssd1 vssd1 vccd1 vccd1 _24529_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_109_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18050_ _18100_/A vssd1 vssd1 vccd1 vccd1 _18793_/A sky130_fd_sc_hd__buf_8
X_15262_ _15262_/A vssd1 vssd1 vccd1 vccd1 _16768_/A sky130_fd_sc_hd__inv_2
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17001_ _24871_/B _21203_/A _20957_/A vssd1 vssd1 vccd1 vccd1 _17002_/A sky130_fd_sc_hd__or3_1
XFILLER_0_35_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14213_ _25829_/Q vssd1 vssd1 vccd1 vccd1 _18794_/B sky130_fd_sc_hd__inv_2
X_15193_ _22552_/B _15812_/B vssd1 vssd1 vccd1 vccd1 _16221_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 _24946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14144_ _14236_/A hold434/X vssd1 vssd1 vccd1 vccd1 hold435/A sky130_fd_sc_hd__nand2_1
XFILLER_0_158_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14075_ hold696/X _14074_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold697/A sky130_fd_sc_hd__a21oi_1
X_18952_ _18952_/A _25773_/Q _18952_/C vssd1 vssd1 vccd1 vccd1 _18953_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_120_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17903_ _25857_/Q _21728_/A vssd1 vssd1 vccd1 vccd1 _17911_/A sky130_fd_sc_hd__or2_2
X_13026_ _26138_/Q _12907_/X _13025_/X vssd1 vssd1 vccd1 vccd1 _13026_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18883_ _18986_/A _19630_/A vssd1 vssd1 vccd1 vccd1 _18883_/Y sky130_fd_sc_hd__nand2_1
X_17834_ _17834_/A _17834_/B vssd1 vssd1 vccd1 vccd1 _17835_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14977_ _14977_/A _14982_/A vssd1 vssd1 vccd1 vccd1 _14977_/Y sky130_fd_sc_hd__nand2_1
X_17765_ _17722_/A _17763_/Y _17764_/X vssd1 vssd1 vccd1 vccd1 _17767_/B sky130_fd_sc_hd__a21boi_1
X_19504_ _19504_/A _21157_/B vssd1 vssd1 vccd1 vccd1 _19504_/Y sky130_fd_sc_hd__nor2_1
X_16716_ _16714_/Y _16715_/Y _16594_/X vssd1 vssd1 vccd1 vccd1 _16716_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13928_ _26286_/Q _13801_/X _13793_/X _13927_/Y vssd1 vssd1 vccd1 vccd1 _13929_/B
+ sky130_fd_sc_hd__a22o_1
X_17696_ _17696_/A _17794_/A vssd1 vssd1 vccd1 vccd1 _17764_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_107_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16647_ _16647_/A _16647_/B vssd1 vssd1 vccd1 vccd1 _16649_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_159_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19435_ _19435_/A _19435_/B vssd1 vssd1 vccd1 vccd1 _19435_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_187_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13859_ _26275_/Q _13801_/X _13793_/X _13858_/Y vssd1 vssd1 vccd1 vccd1 _13860_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16578_ _16555_/A _16597_/A _16577_/Y vssd1 vssd1 vccd1 vccd1 _16580_/A sky130_fd_sc_hd__a21o_1
X_19366_ _19358_/X _19365_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19366_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_186_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15529_ _15529_/A vssd1 vssd1 vccd1 vccd1 _16869_/A sky130_fd_sc_hd__inv_2
X_18317_ _18315_/Y _18316_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25660_/D sky130_fd_sc_hd__a21oi_1
X_19297_ _19452_/A _19297_/B vssd1 vssd1 vccd1 vccd1 _19297_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_5_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18248_ _19045_/B _18248_/B vssd1 vssd1 vccd1 vccd1 _18248_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18179_ _18177_/X _17528_/X _18178_/X vssd1 vssd1 vccd1 vccd1 _18180_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_114_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold502 hold502/A vssd1 vssd1 vccd1 vccd1 hold502/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold513 hold513/A vssd1 vssd1 vccd1 vccd1 hold513/X sky130_fd_sc_hd__dlygate4sd3_1
X_20210_ _21450_/A vssd1 vssd1 vccd1 vccd1 _21449_/A sky130_fd_sc_hd__inv_2
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold524 hold524/A vssd1 vssd1 vccd1 vccd1 hold524/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_29_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21190_ _21189_/B _21190_/B _21190_/C vssd1 vssd1 vccd1 vccd1 _21191_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_123_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold535 hold535/A vssd1 vssd1 vccd1 vccd1 hold535/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 hold546/A vssd1 vssd1 vccd1 vccd1 hold546/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 hold557/A vssd1 vssd1 vccd1 vccd1 hold557/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 hold568/A vssd1 vssd1 vccd1 vccd1 hold568/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20141_ _20141_/A vssd1 vssd1 vccd1 vccd1 _20145_/A sky130_fd_sc_hd__inv_2
Xhold579 hold579/A vssd1 vssd1 vccd1 vccd1 hold579/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20072_ _20072_/A _20072_/B _20981_/B vssd1 vssd1 vccd1 vccd1 _20076_/A sky130_fd_sc_hd__nand3_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1202 _16964_/Y vssd1 vssd1 vccd1 vccd1 _25577_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23900_ _23900_/A vssd1 vssd1 vccd1 vccd1 _26037_/D sky130_fd_sc_hd__clkbuf_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24880_ _24877_/X _24879_/Y _24867_/S _24949_/S vssd1 vssd1 vccd1 vccd1 _24880_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1213 _25813_/Q vssd1 vssd1 vccd1 vccd1 _21331_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1224 _13442_/X vssd1 vssd1 vccd1 vccd1 _25125_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1235 _19527_/Y vssd1 vssd1 vccd1 vccd1 _25738_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1246 _25745_/Q vssd1 vssd1 vccd1 vccd1 _19624_/B sky130_fd_sc_hd__dlygate4sd3_1
X_23831_ hold1900/X _26015_/Q _23831_/S vssd1 vssd1 vccd1 vccd1 _23831_/X sky130_fd_sc_hd__mux2_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1257 _12855_/X vssd1 vssd1 vccd1 vccd1 _25022_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1268 _25049_/Q vssd1 vssd1 vccd1 vccd1 _17536_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 _16978_/Y vssd1 vssd1 vccd1 vccd1 _25579_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23762_ _23762_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23763_/A sky130_fd_sc_hd__and2_1
XFILLER_0_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20974_ _20974_/A _20974_/B vssd1 vssd1 vccd1 vccd1 _21513_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_178_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25501_ _25501_/CLK _25501_/D vssd1 vssd1 vccd1 vccd1 hold860/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22713_ _22713_/A _22900_/B vssd1 vssd1 vccd1 vccd1 _22713_/Y sky130_fd_sc_hd__nand2_1
X_23693_ hold2163/X hold2111/X _23754_/S vssd1 vssd1 vccd1 vccd1 _23694_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_48_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25432_ _25913_/CLK _25432_/D vssd1 vssd1 vccd1 vccd1 _25432_/Q sky130_fd_sc_hd__dfxtp_1
X_22644_ _22645_/B _22645_/A vssd1 vssd1 vccd1 vccd1 _22646_/A sky130_fd_sc_hd__or2_1
XFILLER_0_165_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25363_ _26190_/CLK hold358/X vssd1 vssd1 vccd1 vccd1 hold356/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22575_ _22575_/A _22575_/B vssd1 vssd1 vccd1 vccd1 _22576_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24314_ hold2209/X _26170_/Q _24356_/S vssd1 vssd1 vccd1 vccd1 _24314_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_173_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21526_ _21524_/Y _21525_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21526_/Y sky130_fd_sc_hd__a21oi_1
X_25294_ _26284_/CLK hold49/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24245_ _24245_/A vssd1 vssd1 vccd1 vccd1 _26147_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21457_ _21636_/A _21457_/B _21456_/X vssd1 vssd1 vccd1 vccd1 _21458_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20408_ _20408_/A _20408_/B vssd1 vssd1 vccd1 vccd1 _20410_/A sky130_fd_sc_hd__nand2_1
X_24176_ _24176_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24177_/A sky130_fd_sc_hd__and2_1
XFILLER_0_82_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21388_ _21388_/A _21388_/B vssd1 vssd1 vccd1 vccd1 _21389_/A sky130_fd_sc_hd__nand2_1
Xoutput9 output9/A vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_12
XFILLER_0_43_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23127_ _23127_/A _23127_/B _23191_/C vssd1 vssd1 vccd1 vccd1 _23129_/A sky130_fd_sc_hd__or3_1
X_20339_ _20339_/A _20339_/B vssd1 vssd1 vccd1 vccd1 _20340_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23058_ _23058_/A _23058_/B vssd1 vssd1 vccd1 vccd1 _23059_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_101_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14900_ _14900_/A _14900_/B vssd1 vssd1 vccd1 vccd1 _14900_/Y sky130_fd_sc_hd__nand2_1
X_22009_ _19416_/A _22008_/A _22008_/Y vssd1 vssd1 vccd1 vccd1 _22011_/A sky130_fd_sc_hd__o21ai_1
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15880_ _15881_/B _15881_/A vssd1 vssd1 vccd1 vccd1 _15882_/A sky130_fd_sc_hd__or2_1
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2470 _25681_/Q vssd1 vssd1 vccd1 vccd1 _13289_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14831_ _14900_/A _14831_/B vssd1 vssd1 vccd1 vccd1 _14831_/Y sky130_fd_sc_hd__nand2_1
Xhold2481 _25695_/Q vssd1 vssd1 vccd1 vccd1 _13377_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2492 _25693_/Q vssd1 vssd1 vccd1 vccd1 _13365_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1780 _25887_/Q vssd1 vssd1 vccd1 vccd1 _22971_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17550_ _17624_/A _17550_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17550_/X sky130_fd_sc_hd__and3_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14762_ _14768_/B _21968_/A vssd1 vssd1 vccd1 vccd1 _21967_/B sky130_fd_sc_hd__xnor2_2
Xhold1791 _25871_/Q vssd1 vssd1 vccd1 vccd1 _22689_/B sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16501_ _16501_/A _16501_/B vssd1 vssd1 vccd1 vccd1 _16502_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ _25749_/Q vssd1 vssd1 vccd1 vccd1 _18469_/B sky130_fd_sc_hd__inv_2
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17481_ _17481_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17481_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_98_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14693_ _14693_/A vssd1 vssd1 vccd1 vccd1 _14903_/A sky130_fd_sc_hd__inv_2
XFILLER_0_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16432_ _16473_/A hold933/X vssd1 vssd1 vccd1 vccd1 _16432_/Y sky130_fd_sc_hd__nand2_1
X_19220_ _19220_/A _19220_/B vssd1 vssd1 vccd1 vccd1 _19220_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_168_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13644_ _14120_/A vssd1 vssd1 vccd1 vccd1 _13756_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_184_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19151_ _19186_/A hold605/X vssd1 vssd1 vccd1 vccd1 hold606/A sky130_fd_sc_hd__nand2_1
XFILLER_0_82_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16363_ _16340_/A _16379_/B _16362_/X vssd1 vssd1 vccd1 vccd1 _16365_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_183_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _17813_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13575_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_82_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18102_ _18102_/A _18102_/B _18102_/C vssd1 vssd1 vccd1 vccd1 _21871_/A sky130_fd_sc_hd__nand3_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _16790_/B vssd1 vssd1 vccd1 vccd1 _22734_/B sky130_fd_sc_hd__inv_2
XFILLER_0_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ _15774_/B _15773_/S vssd1 vssd1 vccd1 vccd1 _12527_/A sky130_fd_sc_hd__nand2_8
X_19082_ _19082_/A _19082_/B _22786_/A vssd1 vssd1 vccd1 vccd1 _19082_/X sky130_fd_sc_hd__and3_1
XFILLER_0_42_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16294_ _16294_/A hold863/X _16691_/B vssd1 vssd1 vccd1 vccd1 _16295_/B sky130_fd_sc_hd__and3_1
XFILLER_0_109_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18033_ _18528_/A _25725_/Q vssd1 vssd1 vccd1 vccd1 _18035_/A sky130_fd_sc_hd__nand2_1
X_15245_ _16260_/A _15778_/B vssd1 vssd1 vccd1 vccd1 _16761_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_124_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15176_ _15177_/B _16733_/A vssd1 vssd1 vccd1 vccd1 _15178_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_151_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14127_ _25815_/Q vssd1 vssd1 vccd1 vccd1 _18510_/B sky130_fd_sc_hd__inv_2
XFILLER_0_120_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19984_ _19982_/X _19983_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19984_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14058_ _25804_/Q vssd1 vssd1 vccd1 vccd1 _18288_/B sky130_fd_sc_hd__inv_2
X_18935_ _18955_/A _18935_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18936_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_182_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13009_ _12891_/X _14446_/A _12909_/X _25632_/Q vssd1 vssd1 vccd1 vccd1 _13009_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18866_ _25641_/Q _22615_/B vssd1 vssd1 vccd1 vccd1 _18867_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_98_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17817_ _19038_/A _18372_/A vssd1 vssd1 vccd1 vccd1 _17818_/B sky130_fd_sc_hd__xnor2_4
X_18797_ _18974_/A _19024_/A vssd1 vssd1 vccd1 vccd1 _18798_/B sky130_fd_sc_hd__xnor2_1
X_17748_ _17748_/A _17748_/B vssd1 vssd1 vccd1 vccd1 _17748_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_134_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17679_ _17679_/A _17679_/B vssd1 vssd1 vccd1 vccd1 _17691_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19418_ _20993_/A _19416_/Y _20998_/C vssd1 vssd1 vccd1 vccd1 _19509_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_134_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20690_ _20690_/A _20690_/B vssd1 vssd1 vccd1 vccd1 _20691_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19349_ _19350_/B _19350_/A vssd1 vssd1 vccd1 vccd1 _19349_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22360_ _22786_/A vssd1 vssd1 vccd1 vccd1 _22900_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21311_ _21310_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21311_/X
+ sky130_fd_sc_hd__a211o_1
X_22291_ _22289_/Y _22290_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _22291_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24030_ _24030_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24031_/A sky130_fd_sc_hd__and2_1
X_21242_ _21244_/B _21244_/C vssd1 vssd1 vccd1 vccd1 _21243_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_131_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold310 hold310/A vssd1 vssd1 vccd1 vccd1 hold310/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 hold321/A vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 hold332/A vssd1 vssd1 vccd1 vccd1 hold332/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold343 hold343/A vssd1 vssd1 vccd1 vccd1 hold343/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 hold354/A vssd1 vssd1 vccd1 vccd1 hold354/X sky130_fd_sc_hd__dlygate4sd3_1
X_21173_ _21173_/A _21173_/B vssd1 vssd1 vccd1 vccd1 _21174_/A sky130_fd_sc_hd__nand2_1
Xhold365 hold365/A vssd1 vssd1 vccd1 vccd1 hold365/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 hold376/A vssd1 vssd1 vccd1 vccd1 hold376/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold387 hold387/A vssd1 vssd1 vccd1 vccd1 hold387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 hold398/A vssd1 vssd1 vccd1 vccd1 hold398/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_20124_ _26279_/Q hold707/X vssd1 vssd1 vccd1 vccd1 _20124_/Y sky130_fd_sc_hd__nand2_1
X_25981_ _26004_/CLK _25981_/D vssd1 vssd1 vccd1 vccd1 _25981_/Q sky130_fd_sc_hd__dfxtp_1
X_24932_ _24957_/S _24932_/B vssd1 vssd1 vccd1 vccd1 _24932_/Y sky130_fd_sc_hd__nor2_1
X_20055_ _20055_/A _20055_/B vssd1 vssd1 vccd1 vccd1 _20058_/B sky130_fd_sc_hd__nand2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1010 _13181_/X vssd1 vssd1 vccd1 vccd1 _25083_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1021 _25102_/Q vssd1 vssd1 vccd1 vccd1 _18759_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 _19439_/Y vssd1 vssd1 vccd1 vccd1 _25732_/D sky130_fd_sc_hd__dlygate4sd3_1
X_24863_ _15589_/A _15604_/A _24863_/S vssd1 vssd1 vccd1 vccd1 _24863_/X sky130_fd_sc_hd__mux2_1
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1043 _25024_/Q vssd1 vssd1 vccd1 vccd1 _17322_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1054 _12762_/X vssd1 vssd1 vccd1 vccd1 _25004_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1065 _25127_/Q vssd1 vssd1 vccd1 vccd1 _19068_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1076 _19555_/Y vssd1 vssd1 vccd1 vccd1 _25740_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23814_ _23814_/A vssd1 vssd1 vccd1 vccd1 _26009_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 _25113_/Q vssd1 vssd1 vccd1 vccd1 _18968_/B sky130_fd_sc_hd__dlygate4sd3_1
X_24794_ _24794_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24795_/A sky130_fd_sc_hd__and2_1
Xhold1098 _12960_/X vssd1 vssd1 vccd1 vccd1 _25042_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23745_ _14743_/B _25987_/Q _23754_/S vssd1 vssd1 vccd1 vccd1 _23745_/X sky130_fd_sc_hd__mux2_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20957_ _20957_/A vssd1 vssd1 vccd1 vccd1 _20957_/X sky130_fd_sc_hd__buf_8
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23676_ _23676_/A vssd1 vssd1 vccd1 vccd1 _25964_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20888_ _20888_/A _20888_/B vssd1 vssd1 vccd1 vccd1 _20890_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25415_ _25859_/CLK _25415_/D vssd1 vssd1 vccd1 vccd1 _25415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22627_ _22627_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _22627_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_113_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25346_ _26299_/CLK hold73/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dfxtp_1
X_13360_ _26323_/Q _19687_/A vssd1 vssd1 vccd1 vccd1 _14635_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_180_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22558_ _16743_/B _22421_/X _22552_/X _22553_/Y _22557_/X vssd1 vssd1 vccd1 vccd1
+ _22559_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21509_ _21573_/A _21509_/B vssd1 vssd1 vccd1 vccd1 _21509_/Y sky130_fd_sc_hd__nand2_1
X_25277_ _26232_/CLK hold325/X vssd1 vssd1 vccd1 vccd1 hold323/A sky130_fd_sc_hd__dfxtp_1
X_13291_ _13220_/X _14602_/A _13242_/X _19532_/A vssd1 vssd1 vccd1 vccd1 _13291_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22489_ _18776_/A _25828_/Q _22487_/Y _22488_/Y vssd1 vssd1 vccd1 vccd1 _22490_/B
+ sky130_fd_sc_hd__a31o_1
X_15030_ _15030_/A _15030_/B vssd1 vssd1 vccd1 vccd1 _15031_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_122_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24228_ hold2263/X _26142_/Q _24279_/S vssd1 vssd1 vccd1 vccd1 _24228_/X sky130_fd_sc_hd__mux2_1
X_24159_ _24159_/A vssd1 vssd1 vccd1 vccd1 _26119_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16981_ _15813_/A _16980_/Y _15621_/A vssd1 vssd1 vccd1 vccd1 _16981_/Y sky130_fd_sc_hd__a21oi_1
X_18720_ _18718_/X _18269_/X _18719_/X vssd1 vssd1 vccd1 vccd1 _18721_/A sky130_fd_sc_hd__a21o_1
X_15932_ _15932_/A _15932_/B vssd1 vssd1 vccd1 vccd1 _15933_/B sky130_fd_sc_hd__nand2_1
X_15863_ hold774/X vssd1 vssd1 vccd1 vccd1 _15866_/B sky130_fd_sc_hd__inv_2
X_18651_ _18792_/A _25758_/Q vssd1 vssd1 vccd1 vccd1 _18653_/A sky130_fd_sc_hd__nand2_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14814_ _14812_/Y _14813_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14814_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17602_ _17624_/A _17602_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _17602_/X sky130_fd_sc_hd__and3_1
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15794_ _23172_/B _15812_/B vssd1 vssd1 vccd1 vccd1 _16676_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_118_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18582_ _19673_/A vssd1 vssd1 vccd1 vccd1 _22267_/B sky130_fd_sc_hd__inv_2
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14745_ _21899_/B _15543_/B vssd1 vssd1 vccd1 vccd1 _14746_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_114_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17533_ _17531_/Y _17532_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _17533_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17464_ _17624_/A _17464_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17464_/X sky130_fd_sc_hd__and3_1
X_14676_ _14688_/A hold230/X vssd1 vssd1 vccd1 vccd1 hold231/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16415_ _16439_/B vssd1 vssd1 vccd1 vccd1 _16420_/B sky130_fd_sc_hd__inv_2
XFILLER_0_117_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19203_ _19202_/Y _19130_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19205_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13627_ _26238_/Q _13612_/X _13605_/X _13626_/Y vssd1 vssd1 vccd1 vccd1 _13628_/B
+ sky130_fd_sc_hd__a22o_1
X_17395_ _17395_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17395_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_8__f_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_8__f_clk/X
+ sky130_fd_sc_hd__clkbuf_16
X_16346_ _16346_/A hold968/X _16691_/B vssd1 vssd1 vccd1 vccd1 _16347_/B sky130_fd_sc_hd__and3_1
XFILLER_0_27_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19134_ _21228_/A vssd1 vssd1 vccd1 vccd1 _19134_/X sky130_fd_sc_hd__buf_8
X_13558_ _13583_/A _13558_/B vssd1 vssd1 vccd1 vccd1 _13558_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12509_ _24979_/Q _24978_/Q _24976_/Q _24977_/Q vssd1 vssd1 vccd1 vccd1 _12515_/B
+ sky130_fd_sc_hd__or4_1
X_19065_ _19063_/Y _19064_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25706_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16277_ _16171_/B _16272_/B _16275_/X _16276_/Y vssd1 vssd1 vccd1 vccd1 _16277_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_140_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13489_ _26216_/Q _13426_/X _13468_/X _13488_/Y vssd1 vssd1 vccd1 vccd1 _13490_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15228_ hold885/X _15230_/A vssd1 vssd1 vccd1 vccd1 _15232_/A sky130_fd_sc_hd__nor2_1
X_18016_ _25843_/Q vssd1 vssd1 vccd1 vccd1 _20214_/B sky130_fd_sc_hd__inv_2
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15159_ _15159_/A vssd1 vssd1 vccd1 vccd1 _16726_/A sky130_fd_sc_hd__inv_2
XFILLER_0_140_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19967_ _19966_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19969_/A
+ sky130_fd_sc_hd__a211o_1
X_18918_ _19017_/B _19066_/B vssd1 vssd1 vccd1 vccd1 _18919_/B sky130_fd_sc_hd__xnor2_1
X_19898_ _19999_/A _18908_/A _20004_/C vssd1 vssd1 vccd1 vccd1 _19970_/A sky130_fd_sc_hd__o21a_2
X_18849_ _18951_/A _18853_/B vssd1 vssd1 vccd1 vccd1 _18851_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_179_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21860_ _21858_/X _21859_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _21860_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20811_ _20810_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20811_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21791_ _21791_/A vssd1 vssd1 vccd1 vccd1 _21791_/X sky130_fd_sc_hd__buf_4
XFILLER_0_49_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23530_ _23524_/X _23529_/X _24867_/S vssd1 vssd1 vccd1 vccd1 _23530_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20742_ _20745_/A _20745_/C vssd1 vssd1 vccd1 vccd1 _20743_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23461_ hold56/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23461_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_163_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20673_ _20673_/A _20673_/B vssd1 vssd1 vccd1 vccd1 _20677_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_107_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25200_ _26281_/CLK hold685/X vssd1 vssd1 vccd1 vccd1 hold683/A sky130_fd_sc_hd__dfxtp_1
X_22412_ _22413_/B _22413_/A vssd1 vssd1 vccd1 vccd1 _22414_/A sky130_fd_sc_hd__or2_1
XFILLER_0_61_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26180_ _26181_/CLK _26180_/D vssd1 vssd1 vccd1 vccd1 _26180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23392_ hold140/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23392_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25131_ _25711_/CLK hold499/X vssd1 vssd1 vccd1 vccd1 hold497/A sky130_fd_sc_hd__dfxtp_1
X_22343_ _22653_/A _22343_/B vssd1 vssd1 vccd1 vccd1 _22343_/X sky130_fd_sc_hd__or2_1
XFILLER_0_115_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25062_ _26148_/CLK _25062_/D vssd1 vssd1 vccd1 vccd1 _25062_/Q sky130_fd_sc_hd__dfxtp_1
X_22274_ _22890_/B vssd1 vssd1 vccd1 vccd1 _22496_/A sky130_fd_sc_hd__inv_2
XFILLER_0_20_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24013_ _24013_/A vssd1 vssd1 vccd1 vccd1 _26072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold140 hold140/A vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__dlygate4sd3_1
X_21225_ _21225_/A _21225_/B _21225_/C vssd1 vssd1 vccd1 vccd1 _21226_/B sky130_fd_sc_hd__nand3_1
Xhold151 hold151/A vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold162 hold162/A vssd1 vssd1 vccd1 vccd1 hold162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 hold173/A vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold184 hold184/A vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
X_21156_ _21156_/A _21913_/B vssd1 vssd1 vccd1 vccd1 _21157_/A sky130_fd_sc_hd__nand2_1
Xhold195 hold195/A vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
X_20107_ _20107_/A _20107_/B vssd1 vssd1 vccd1 vccd1 _21402_/A sky130_fd_sc_hd__nand2_4
X_25964_ _26042_/CLK _25964_/D vssd1 vssd1 vccd1 vccd1 _25964_/Q sky130_fd_sc_hd__dfxtp_1
X_21087_ _21577_/C _21532_/B vssd1 vssd1 vccd1 vccd1 _21089_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_176_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24915_ _16390_/B _16399_/Y _24944_/S vssd1 vssd1 vccd1 vccd1 _24915_/X sky130_fd_sc_hd__mux2_1
X_20038_ _21042_/A _20038_/B _20037_/X vssd1 vssd1 vccd1 vccd1 _20039_/B sky130_fd_sc_hd__or3b_1
X_25895_ _25895_/CLK _25895_/D vssd1 vssd1 vccd1 vccd1 _25895_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24846_ _15305_/B _15320_/B _24860_/S vssd1 vssd1 vccd1 vccd1 _24846_/X sky130_fd_sc_hd__mux2_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ _12840_/X _12858_/X _12827_/X _12859_/X vssd1 vssd1 vccd1 vccd1 _12860_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12791_ _25010_/Q _14264_/A vssd1 vssd1 vccd1 vccd1 _12791_/X sky130_fd_sc_hd__or2_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24777_ _24777_/A vssd1 vssd1 vccd1 vccd1 _26320_/D sky130_fd_sc_hd__clkbuf_1
X_21989_ _22729_/A vssd1 vssd1 vccd1 vccd1 _22245_/A sky130_fd_sc_hd__inv_2
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14590_/A vssd1 vssd1 vccd1 vccd1 _14585_/A sky130_fd_sc_hd__clkbuf_8
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23728_ _23728_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23729_/A sky130_fd_sc_hd__and2_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _14461_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14461_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_95_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23659_ hold2109/X hold1936/X _23677_/S vssd1 vssd1 vccd1 vccd1 _23660_/A sky130_fd_sc_hd__mux2_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16200_ _16188_/Y _16190_/Y _16214_/A _16199_/Y vssd1 vssd1 vccd1 vccd1 _16200_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13412_ _13315_/X _13410_/X _23629_/B _13411_/X vssd1 vssd1 vccd1 vccd1 hold974/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17180_ _20741_/B _25857_/Q _25793_/Q vssd1 vssd1 vccd1 vccd1 _17181_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_187_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14392_ _14404_/A hold47/X vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__nand2_1
XFILLER_0_52_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16131_ _16125_/B _16134_/B _16124_/A vssd1 vssd1 vccd1 vccd1 _16161_/A sky130_fd_sc_hd__o21ai_1
X_25329_ _25650_/CLK hold67/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dfxtp_1
X_13343_ _13220_/X _14626_/A _13242_/X _19644_/A vssd1 vssd1 vccd1 vccd1 _13343_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16062_ _16160_/A _16062_/B vssd1 vssd1 vccd1 vccd1 _16071_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_106_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13274_ _26181_/Q _13239_/X _13273_/X vssd1 vssd1 vccd1 vccd1 _13274_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_59_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15013_ _15013_/A _15013_/B vssd1 vssd1 vccd1 vccd1 _15034_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_121_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19821_ _19821_/A _19821_/B vssd1 vssd1 vccd1 vccd1 _19821_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_166_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19752_ _19975_/A _19752_/B vssd1 vssd1 vccd1 vccd1 _19752_/Y sky130_fd_sc_hd__nand2_1
X_16964_ _16962_/Y _16963_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _16964_/Y sky130_fd_sc_hd__a21oi_1
X_18703_ _18701_/Y _18702_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25679_/D sky130_fd_sc_hd__a21oi_1
X_15915_ hold551/X vssd1 vssd1 vccd1 vccd1 _15918_/B sky130_fd_sc_hd__inv_2
XFILLER_0_21_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19683_ _26253_/Q _19483_/X hold925/X vssd1 vssd1 vccd1 vccd1 _19683_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16895_ _16935_/A _16900_/B vssd1 vssd1 vccd1 vccd1 _16897_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_155_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18634_ _20330_/B _22329_/A vssd1 vssd1 vccd1 vccd1 _20321_/A sky130_fd_sc_hd__nand2_2
X_15846_ _15869_/B _15846_/B vssd1 vssd1 vccd1 vccd1 _15857_/A sky130_fd_sc_hd__or2_1
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18565_ _18565_/A _18565_/B vssd1 vssd1 vccd1 vccd1 _22236_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_188_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15777_ _15777_/A vssd1 vssd1 vccd1 vccd1 _16665_/A sky130_fd_sc_hd__inv_2
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ _26131_/Q _12907_/X _12988_/X vssd1 vssd1 vccd1 vccd1 _12989_/X sky130_fd_sc_hd__a21o_1
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17516_ _17516_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17516_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_185_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14728_ _25841_/Q _12527_/A _14923_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14728_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_185_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18496_ _18494_/X _18269_/X _18495_/X vssd1 vssd1 vccd1 vccd1 _18497_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_115_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14659_ _14657_/Y hold42/X _14646_/X vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__a21oi_1
X_17447_ _17498_/A _17615_/B vssd1 vssd1 vccd1 vccd1 _17448_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_180_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _25784_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17378_ _25617_/Q vssd1 vssd1 vccd1 vccd1 _21211_/B sky130_fd_sc_hd__inv_2
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19117_ _20284_/A _21992_/A _25589_/Q vssd1 vssd1 vccd1 vccd1 _20288_/C sky130_fd_sc_hd__nand3_2
X_16329_ _16676_/A _16329_/B vssd1 vssd1 vccd1 vccd1 _16331_/A sky130_fd_sc_hd__or2_1
XFILLER_0_160_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19048_ _19046_/X _18879_/X _19047_/X vssd1 vssd1 vccd1 vccd1 _19049_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_70_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21010_ _21010_/A _21010_/B _21010_/C vssd1 vssd1 vccd1 vccd1 _21011_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22961_ _22961_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22961_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24700_ _24700_/A vssd1 vssd1 vccd1 vccd1 _26295_/D sky130_fd_sc_hd__clkbuf_1
X_21912_ _21912_/A _25871_/Q vssd1 vssd1 vccd1 vccd1 _21912_/Y sky130_fd_sc_hd__nand2_1
X_25680_ _26313_/CLK _25680_/D vssd1 vssd1 vccd1 vccd1 _25680_/Q sky130_fd_sc_hd__dfxtp_1
X_22892_ _22892_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _22901_/A sky130_fd_sc_hd__nand2_1
X_24631_ _24631_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24632_/A sky130_fd_sc_hd__and2_1
X_21843_ _21843_/A _25869_/Q vssd1 vssd1 vccd1 vccd1 _21843_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_139_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24562_ _24562_/A vssd1 vssd1 vccd1 vccd1 _26250_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21774_ _18266_/A _25803_/Q _21772_/Y _21773_/Y vssd1 vssd1 vccd1 vccd1 _21775_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26301_ _26301_/CLK _26301_/D vssd1 vssd1 vccd1 vccd1 _26301_/Q sky130_fd_sc_hd__dfxtp_2
X_23513_ _23510_/Y _23512_/Y _24858_/S vssd1 vssd1 vccd1 vccd1 _23513_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_65_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20725_ _20725_/A _20725_/B _21335_/C vssd1 vssd1 vccd1 vccd1 _20729_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_93_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_171_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _25791_/CLK sky130_fd_sc_hd__clkbuf_16
X_24493_ _24493_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24494_/A sky130_fd_sc_hd__and2_1
X_26232_ _26232_/CLK _26232_/D vssd1 vssd1 vccd1 vccd1 _26232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23444_ _23441_/Y _23443_/Y _24957_/S vssd1 vssd1 vccd1 vccd1 _23444_/X sky130_fd_sc_hd__mux2_1
X_20656_ _20655_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20656_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26163_ _26164_/CLK _26163_/D vssd1 vssd1 vccd1 vccd1 _26163_/Q sky130_fd_sc_hd__dfxtp_1
X_23375_ _23376_/B _23376_/A vssd1 vssd1 vccd1 vccd1 _23375_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20587_ _20590_/A _20590_/C vssd1 vssd1 vccd1 vccd1 _20588_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25114_ _26198_/CLK _25114_/D vssd1 vssd1 vccd1 vccd1 _25114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22326_ _22326_/A _25885_/Q vssd1 vssd1 vccd1 vccd1 _22326_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_131_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26094_ _26096_/CLK _26094_/D vssd1 vssd1 vccd1 vccd1 hold721/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25045_ _26130_/CLK _25045_/D vssd1 vssd1 vccd1 vccd1 _25045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22257_ _22257_/A _23154_/A _22257_/C vssd1 vssd1 vccd1 vccd1 _22257_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_108_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21208_ _21235_/A _21208_/B vssd1 vssd1 vccd1 vccd1 _21208_/Y sky130_fd_sc_hd__nand2_1
X_22188_ _22676_/A _22840_/B vssd1 vssd1 vccd1 vccd1 _22198_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_100_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21139_ _21610_/C vssd1 vssd1 vccd1 vccd1 _21613_/B sky130_fd_sc_hd__inv_2
XFILLER_0_79_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13961_ hold778/X _13960_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold779/A sky130_fd_sc_hd__a21oi_1
X_25947_ _26012_/CLK _25947_/D vssd1 vssd1 vccd1 vccd1 _25947_/Q sky130_fd_sc_hd__dfxtp_1
X_15700_ _15718_/A _15701_/A vssd1 vssd1 vccd1 vccd1 _15700_/X sky130_fd_sc_hd__or2_1
X_12912_ _17414_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12912_/X sky130_fd_sc_hd__or2_1
X_16680_ _16680_/A _16680_/B vssd1 vssd1 vccd1 vccd1 _16681_/B sky130_fd_sc_hd__nor2_1
X_25878_ _25878_/CLK _25878_/D vssd1 vssd1 vccd1 vccd1 _25878_/Q sky130_fd_sc_hd__dfxtp_2
X_13892_ _13941_/A _13892_/B vssd1 vssd1 vccd1 vccd1 _13892_/Y sky130_fd_sc_hd__nand2_1
X_15631_ _15631_/A vssd1 vssd1 vccd1 vccd1 _15640_/B sky130_fd_sc_hd__inv_2
X_24829_ hold2618/X _26338_/Q _24835_/S vssd1 vssd1 vccd1 vccd1 _24829_/X sky130_fd_sc_hd__mux2_1
X_12843_ _26103_/Q _12748_/X _12842_/X vssd1 vssd1 vccd1 vccd1 _12843_/X sky130_fd_sc_hd__a21o_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15562_ _15562_/A vssd1 vssd1 vccd1 vccd1 _24864_/A sky130_fd_sc_hd__inv_2
XFILLER_0_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18350_ _18350_/A _21156_/A vssd1 vssd1 vccd1 vccd1 _18698_/A sky130_fd_sc_hd__xor2_4
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _12726_/B _14304_/A _12752_/X _25587_/Q vssd1 vssd1 vccd1 vccd1 _12774_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _14525_/A hold125/X vssd1 vssd1 vccd1 vccd1 hold126/A sky130_fd_sc_hd__nand2_1
X_17301_ _25610_/Q vssd1 vssd1 vccd1 vccd1 _21022_/B sky130_fd_sc_hd__inv_2
XFILLER_0_90_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ _16451_/A _16711_/A vssd1 vssd1 vccd1 vccd1 _16855_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18281_ _18445_/A _18287_/B vssd1 vssd1 vccd1 vccd1 _18283_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_162_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _26171_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17232_ _25605_/Q vssd1 vssd1 vccd1 vccd1 _20883_/B sky130_fd_sc_hd__inv_2
X_14444_ _14465_/A hold17/X vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__nand2_1
XFILLER_0_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17163_ _17163_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17163_/Y sky130_fd_sc_hd__nand2_1
X_14375_ _14373_/Y hold87/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16114_ _16125_/B _16114_/B vssd1 vssd1 vccd1 vccd1 _16134_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13326_ _14064_/A vssd1 vssd1 vccd1 vccd1 _13944_/A sky130_fd_sc_hd__clkbuf_16
Xhold909 hold909/A vssd1 vssd1 vccd1 vccd1 hold909/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17094_ _17092_/X _23187_/B _17093_/X vssd1 vssd1 vccd1 vccd1 _17095_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_80_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16045_ _16043_/X hold705/X _15805_/X vssd1 vssd1 vccd1 vccd1 hold706/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13257_ _18618_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13257_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13188_ _13188_/A vssd1 vssd1 vccd1 vccd1 _19303_/A sky130_fd_sc_hd__buf_4
XFILLER_0_23_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19804_ _20596_/A _19802_/Y _20601_/C vssd1 vssd1 vccd1 vccd1 _19888_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_23_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17996_ _17996_/A _17996_/B vssd1 vssd1 vccd1 vccd1 _21800_/A sky130_fd_sc_hd__nand2_1
Xhold1609 _17468_/Y vssd1 vssd1 vccd1 vccd1 _25619_/D sky130_fd_sc_hd__dlygate4sd3_1
X_19735_ _19733_/X _19734_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19735_/Y sky130_fd_sc_hd__a21oi_1
X_16947_ _16945_/X _16711_/X _16946_/Y _25896_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16948_/A sky130_fd_sc_hd__a32o_1
X_19666_ _19658_/X _19665_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19666_/Y sky130_fd_sc_hd__o21ai_1
X_16878_ _16878_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16878_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_95_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18617_ _18617_/A _18617_/B vssd1 vssd1 vccd1 vccd1 _18617_/X sky130_fd_sc_hd__xor2_1
X_15829_ _15829_/A _15829_/B vssd1 vssd1 vccd1 vccd1 _15834_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_189_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19597_ _19595_/Y _19596_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19597_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18548_ _18548_/A _25817_/Q _18548_/C vssd1 vssd1 vccd1 vccd1 _20171_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18479_ _18477_/Y _18478_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25668_/D sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_153_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _26302_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_63_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20510_ _25851_/Q vssd1 vssd1 vccd1 vccd1 _22165_/B sky130_fd_sc_hd__inv_2
XFILLER_0_7_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21490_ _21490_/A _21490_/B vssd1 vssd1 vccd1 vccd1 _21491_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20441_ _20441_/A _25888_/Q vssd1 vssd1 vccd1 vccd1 _20447_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_172_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23160_ _23159_/A _22849_/X _23159_/B vssd1 vssd1 vccd1 vccd1 _23161_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20372_ _21198_/B _21515_/A vssd1 vssd1 vccd1 vccd1 _20375_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22111_ _22109_/X _22110_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _22111_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23091_ _23091_/A _23187_/B vssd1 vssd1 vccd1 vccd1 _23091_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_101_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22042_ _22042_/A _22042_/B vssd1 vssd1 vccd1 vccd1 _22042_/Y sky130_fd_sc_hd__nand2_1
X_25801_ _25802_/CLK _25801_/D vssd1 vssd1 vccd1 vccd1 _25801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23993_ _23993_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23994_/A sky130_fd_sc_hd__and2_1
X_25732_ _25738_/CLK _25732_/D vssd1 vssd1 vccd1 vccd1 _25732_/Q sky130_fd_sc_hd__dfxtp_1
X_22944_ _22944_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22944_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_168_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25663_ _26297_/CLK _25663_/D vssd1 vssd1 vccd1 vccd1 _25663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22875_ _22875_/A _23184_/B vssd1 vssd1 vccd1 vccd1 _22876_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24614_ _24614_/A vssd1 vssd1 vccd1 vccd1 _26267_/D sky130_fd_sc_hd__clkbuf_1
X_21826_ _21824_/X _21825_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _21826_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25594_ _25594_/CLK _25594_/D vssd1 vssd1 vccd1 vccd1 _25594_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_149_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24545_ _24545_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24546_/A sky130_fd_sc_hd__and2_1
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21757_ _22058_/A _21757_/B vssd1 vssd1 vccd1 vccd1 _21757_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_144_clk clkbuf_4_11__f_clk/X vssd1 vssd1 vccd1 vccd1 _25687_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_176_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20708_ _20707_/B _20708_/B _20708_/C vssd1 vssd1 vccd1 vccd1 _20709_/B sky130_fd_sc_hd__nand3b_1
X_12490_ _24745_/A vssd1 vssd1 vccd1 vccd1 _24836_/B sky130_fd_sc_hd__buf_8
XFILLER_0_149_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24476_ _24476_/A vssd1 vssd1 vccd1 vccd1 _26222_/D sky130_fd_sc_hd__clkbuf_1
X_21688_ _21686_/Y _21687_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21688_/Y sky130_fd_sc_hd__a21oi_1
X_26215_ _26216_/CLK _26215_/D vssd1 vssd1 vccd1 vccd1 _26215_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_136_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23427_ hold86/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23427_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20639_ _20639_/A _22518_/B _20639_/C vssd1 vssd1 vccd1 vccd1 _20643_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26146_ _26146_/CLK _26146_/D vssd1 vssd1 vccd1 vccd1 _26146_/Q sky130_fd_sc_hd__dfxtp_1
X_14160_ _26323_/Q _13988_/X _13981_/X _14159_/Y vssd1 vssd1 vccd1 vccd1 _14161_/B
+ sky130_fd_sc_hd__a22o_1
X_23358_ _23358_/A vssd1 vssd1 vccd1 vccd1 _25934_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13111_ _13049_/X _14506_/A _13067_/X _25651_/Q vssd1 vssd1 vccd1 vccd1 _13111_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22309_ _17849_/A _25792_/Q _22307_/Y _22308_/Y vssd1 vssd1 vccd1 vccd1 _22310_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26077_ _26079_/CLK _26077_/D vssd1 vssd1 vccd1 vccd1 _26077_/Q sky130_fd_sc_hd__dfxtp_1
X_14091_ _26312_/Q _13988_/X _13981_/X _14090_/Y vssd1 vssd1 vccd1 vccd1 _14092_/B
+ sky130_fd_sc_hd__a22o_1
X_23289_ hold855/X _23290_/A vssd1 vssd1 vccd1 vccd1 _23289_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25028_ _26116_/CLK _25028_/D vssd1 vssd1 vccd1 vccd1 _25028_/Q sky130_fd_sc_hd__dfxtp_1
X_13042_ _17602_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13042_/X sky130_fd_sc_hd__or2_1
X_17850_ _25657_/Q _20429_/B vssd1 vssd1 vccd1 vccd1 _17853_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_100_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16801_ _16935_/A _16806_/B vssd1 vssd1 vccd1 vccd1 _16803_/B sky130_fd_sc_hd__nand2_1
X_17781_ _17781_/A _17781_/B _17781_/C vssd1 vssd1 vccd1 vccd1 _17784_/A sky130_fd_sc_hd__nand3_1
X_14993_ _14993_/A _14998_/B vssd1 vssd1 vccd1 vccd1 _14993_/Y sky130_fd_sc_hd__nand2_1
X_19520_ _21183_/A _19518_/Y _21187_/C vssd1 vssd1 vccd1 vccd1 _19607_/B sky130_fd_sc_hd__o21a_2
X_16732_ _16733_/B _16733_/A vssd1 vssd1 vccd1 vccd1 _16732_/X sky130_fd_sc_hd__or2_1
X_13944_ _13944_/A vssd1 vssd1 vccd1 vccd1 _14061_/A sky130_fd_sc_hd__clkbuf_8
X_19451_ _19443_/X _19450_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19451_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16663_ _16661_/X _16662_/Y _16594_/X vssd1 vssd1 vccd1 vccd1 hold943/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13875_ _20085_/B vssd1 vssd1 vccd1 vccd1 _17834_/B sky130_fd_sc_hd__inv_2
X_18402_ _25874_/Q _22014_/A vssd1 vssd1 vccd1 vccd1 _18411_/A sky130_fd_sc_hd__or2_2
X_15614_ _15612_/Y _15578_/X _15613_/Y vssd1 vssd1 vccd1 vccd1 _15695_/A sky130_fd_sc_hd__o21ai_1
X_12826_ _26100_/Q _12748_/X _12825_/X vssd1 vssd1 vccd1 vccd1 _12826_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_186_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19382_ _21099_/A vssd1 vssd1 vccd1 vccd1 _19382_/X sky130_fd_sc_hd__buf_8
X_16594_ _17568_/A vssd1 vssd1 vccd1 vccd1 _16594_/X sky130_fd_sc_hd__buf_6
XFILLER_0_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18333_ _18535_/A _18333_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _18333_/X sky130_fd_sc_hd__and3_1
X_15545_ _15546_/B _15546_/A vssd1 vssd1 vccd1 vccd1 _15548_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_127_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12757_ _12746_/X _12754_/X _14910_/B _12756_/X vssd1 vssd1 vccd1 vccd1 _12757_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_135_clk clkbuf_leaf_82_clk/A vssd1 vssd1 vccd1 vccd1 _25822_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15476_ _15621_/A _16435_/B vssd1 vssd1 vccd1 vccd1 _15479_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18264_ _18264_/A _18264_/B _18264_/C vssd1 vssd1 vccd1 vccd1 _21775_/A sky130_fd_sc_hd__nand3_2
X_12688_ _12688_/A vssd1 vssd1 vccd1 vccd1 _24989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17215_ _17213_/X _23187_/B _17214_/X vssd1 vssd1 vccd1 vccd1 _17216_/A sky130_fd_sc_hd__a21o_1
X_14427_ _14425_/Y hold216/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold217/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_181_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18195_ _20965_/B _19402_/A vssd1 vssd1 vccd1 vccd1 _18196_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_142_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17146_ _17478_/A _17555_/A vssd1 vssd1 vccd1 vccd1 _17147_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14358_ _14358_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14358_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold706 hold706/A vssd1 vssd1 vccd1 vccd1 hold706/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold717 hold717/A vssd1 vssd1 vccd1 vccd1 hold717/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 hold728/A vssd1 vssd1 vccd1 vccd1 hold728/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13309_ _13309_/A vssd1 vssd1 vccd1 vccd1 _19574_/A sky130_fd_sc_hd__clkbuf_8
X_17077_ _17393_/A hold960/X _19994_/B vssd1 vssd1 vccd1 vccd1 _17077_/X sky130_fd_sc_hd__and3_1
X_14289_ _14688_/A vssd1 vssd1 vccd1 vccd1 _14344_/A sky130_fd_sc_hd__buf_6
Xhold739 hold739/A vssd1 vssd1 vccd1 vccd1 hold739/X sky130_fd_sc_hd__buf_1
X_16028_ _16028_/A _16028_/B vssd1 vssd1 vccd1 vccd1 _16028_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_27_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2107 _12690_/Y vssd1 vssd1 vccd1 vccd1 _12692_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2118 _25953_/Q vssd1 vssd1 vccd1 vccd1 hold2118/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2129 _23702_/X vssd1 vssd1 vccd1 vccd1 _23703_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1406 _13358_/X vssd1 vssd1 vccd1 vccd1 _25111_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1417 _25408_/Q vssd1 vssd1 vccd1 vccd1 _14873_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1428 _16800_/Y vssd1 vssd1 vccd1 vccd1 _25553_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17979_ _19046_/A vssd1 vssd1 vccd1 vccd1 _18997_/A sky130_fd_sc_hd__inv_2
Xhold1439 _25055_/Q vssd1 vssd1 vccd1 vccd1 _17580_/B sky130_fd_sc_hd__dlygate4sd3_1
X_19718_ _19734_/B _19807_/B vssd1 vssd1 vccd1 vccd1 _19720_/A sky130_fd_sc_hd__xnor2_1
X_20990_ _20990_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _20990_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19649_ _19649_/A _19649_/B vssd1 vssd1 vccd1 vccd1 _19649_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22660_ _22660_/A _22900_/B vssd1 vssd1 vccd1 vccd1 _22660_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_133_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21611_ _21611_/A _21660_/B vssd1 vssd1 vccd1 vccd1 _21613_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_126_clk clkbuf_4_11__f_clk/X vssd1 vssd1 vccd1 vccd1 _25817_/CLK sky130_fd_sc_hd__clkbuf_16
X_22591_ _18856_/A _25832_/Q _22589_/Y _22590_/Y vssd1 vssd1 vccd1 vccd1 _22592_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24330_ _24330_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24331_/A sky130_fd_sc_hd__and2_1
X_21542_ _21540_/Y _21541_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21542_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24261_ _26152_/Q hold2235/X _24279_/S vssd1 vssd1 vccd1 vccd1 _24261_/X sky130_fd_sc_hd__mux2_1
X_21473_ _21636_/A _21473_/B _21472_/X vssd1 vssd1 vccd1 vccd1 _21474_/B sky130_fd_sc_hd__or3b_1
X_26000_ _26001_/CLK _26000_/D vssd1 vssd1 vccd1 vccd1 _26000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23212_ _23212_/A _23212_/B vssd1 vssd1 vccd1 vccd1 _23213_/A sky130_fd_sc_hd__nand2_1
X_20424_ _20424_/A _20424_/B vssd1 vssd1 vccd1 vccd1 _20425_/A sky130_fd_sc_hd__nand2_1
X_24192_ _24192_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24193_/A sky130_fd_sc_hd__and2_1
XFILLER_0_31_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23143_ _23143_/A _23143_/B _23191_/C vssd1 vssd1 vccd1 vccd1 _23145_/A sky130_fd_sc_hd__or3_1
XFILLER_0_141_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20355_ _20358_/A _20358_/C vssd1 vssd1 vccd1 vccd1 _20356_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_109_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23074_ _23074_/A _23074_/B vssd1 vssd1 vccd1 vccd1 _23075_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20286_ _20288_/B _20288_/C vssd1 vssd1 vccd1 vccd1 _20287_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22025_ _25846_/Q _25782_/Q vssd1 vssd1 vccd1 vccd1 _22026_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_179_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2630 _26227_/Q vssd1 vssd1 vccd1 vccd1 hold2630/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2641 _26318_/Q vssd1 vssd1 vccd1 vccd1 hold2641/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2652 _26285_/Q vssd1 vssd1 vccd1 vccd1 hold2652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2663 _26275_/Q vssd1 vssd1 vccd1 vccd1 hold2663/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2674 _26296_/Q vssd1 vssd1 vccd1 vccd1 hold2674/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1940 _25260_/Q vssd1 vssd1 vccd1 vccd1 _12733_/A sky130_fd_sc_hd__buf_1
Xhold2685 _24814_/X vssd1 vssd1 vccd1 vccd1 _24815_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1951 _25427_/Q vssd1 vssd1 vccd1 vccd1 _15021_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
X_23976_ _23976_/A vssd1 vssd1 vccd1 vccd1 _26060_/D sky130_fd_sc_hd__clkbuf_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2696 _26243_/Q vssd1 vssd1 vccd1 vccd1 hold2696/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1962 _24222_/X vssd1 vssd1 vccd1 vccd1 _24223_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1973 _24139_/X vssd1 vssd1 vccd1 vccd1 _24140_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1984 _24965_/Q vssd1 vssd1 vccd1 vccd1 _12559_/A sky130_fd_sc_hd__dlygate4sd3_1
X_22927_ _22927_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22927_/Y sky130_fd_sc_hd__nand2_1
X_25715_ _25716_/CLK _25715_/D vssd1 vssd1 vccd1 vccd1 _25715_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1995 _26151_/Q vssd1 vssd1 vccd1 vccd1 hold1995/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13660_ _13703_/A _13660_/B vssd1 vssd1 vccd1 vccd1 _13660_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22858_ _23167_/B _22858_/B vssd1 vssd1 vccd1 vccd1 _22860_/A sky130_fd_sc_hd__nand2_1
X_25646_ _25712_/CLK _25646_/D vssd1 vssd1 vccd1 vccd1 _25646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _12702_/A hold869/X _12613_/A vssd1 vssd1 vccd1 vccd1 hold870/A sky130_fd_sc_hd__nor3_1
XFILLER_0_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21809_ _21809_/A _25868_/Q vssd1 vssd1 vccd1 vccd1 _21809_/Y sky130_fd_sc_hd__nand2_1
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25577_ _26066_/CLK _25577_/D vssd1 vssd1 vccd1 vccd1 _25577_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_117_clk clkbuf_4_14__f_clk/X vssd1 vssd1 vccd1 vccd1 _25378_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13591_ hold591/X _13590_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold592/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22789_ _22937_/A _22789_/B vssd1 vssd1 vccd1 vccd1 _22789_/Y sky130_fd_sc_hd__nand2_1
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _15327_/B _15308_/X _15329_/Y vssd1 vssd1 vccd1 vccd1 _15408_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_108_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ _12542_/A vssd1 vssd1 vccd1 vccd1 _24996_/D sky130_fd_sc_hd__inv_2
X_24528_ _24528_/A vssd1 vssd1 vccd1 vccd1 _26239_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15261_ _15261_/A vssd1 vssd1 vccd1 vccd1 _15263_/A sky130_fd_sc_hd__inv_2
XFILLER_0_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24459_ _24459_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24460_/A sky130_fd_sc_hd__and2_1
XFILLER_0_136_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14212_ _14236_/A hold751/X vssd1 vssd1 vccd1 vccd1 hold752/A sky130_fd_sc_hd__nand2_1
XFILLER_0_123_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17000_ _21042_/A vssd1 vssd1 vccd1 vccd1 _23187_/B sky130_fd_sc_hd__clkbuf_16
X_15192_ _22555_/B _15192_/B vssd1 vssd1 vccd1 vccd1 _22552_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_149_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_8 _24946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26129_ _26130_/CLK _26129_/D vssd1 vssd1 vccd1 vccd1 _26129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14143_ hold749/X _14142_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold750/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14074_ _14180_/A _14074_/B vssd1 vssd1 vccd1 vccd1 _14074_/Y sky130_fd_sc_hd__nand2_1
X_18951_ _18951_/A _18955_/B vssd1 vssd1 vccd1 vccd1 _18953_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17902_ _17902_/A _17902_/B vssd1 vssd1 vccd1 vccd1 _21728_/A sky130_fd_sc_hd__nand2_1
X_13025_ _12891_/X _14455_/A _12909_/X _25635_/Q vssd1 vssd1 vccd1 vccd1 _13025_/X
+ sky130_fd_sc_hd__a22o_1
X_18882_ _18882_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18882_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17833_ _17834_/B _17834_/A vssd1 vssd1 vccd1 vccd1 _20070_/A sky130_fd_sc_hd__or2_2
XFILLER_0_174_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17764_ _17764_/A _17764_/B vssd1 vssd1 vccd1 vccd1 _17764_/X sky130_fd_sc_hd__or2_1
X_14976_ _14982_/A _14977_/A vssd1 vssd1 vccd1 vccd1 _14976_/X sky130_fd_sc_hd__or2_1
X_19503_ _19500_/Y _19503_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19503_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_107_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16715_ _16858_/A _16715_/B vssd1 vssd1 vccd1 vccd1 _16715_/Y sky130_fd_sc_hd__nand2_1
X_13927_ _18189_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13927_/Y sky130_fd_sc_hd__nor2_1
X_17695_ _17750_/B _25906_/Q vssd1 vssd1 vccd1 vccd1 _17696_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19434_ _19435_/B _19435_/A vssd1 vssd1 vccd1 vccd1 _19434_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16646_ _16644_/Y _16645_/Y _16594_/X vssd1 vssd1 vccd1 vccd1 hold921/A sky130_fd_sc_hd__a21oi_1
X_13858_ _18935_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13858_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_159_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12809_ _12726_/B _14325_/A _12752_/X _25594_/Q vssd1 vssd1 vccd1 vccd1 _12809_/X
+ sky130_fd_sc_hd__a22o_1
X_19365_ _19363_/X _19364_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19365_/Y sky130_fd_sc_hd__a21oi_1
X_16577_ _16577_/A vssd1 vssd1 vccd1 vccd1 _16577_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_108_clk clkbuf_4_14__f_clk/X vssd1 vssd1 vccd1 vccd1 _25420_/CLK sky130_fd_sc_hd__clkbuf_16
X_13789_ _26264_/Q _13612_/X _13605_/X _13788_/Y vssd1 vssd1 vccd1 vccd1 _13790_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18316_ _18641_/A _19230_/A vssd1 vssd1 vccd1 vccd1 _18316_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15528_ _15528_/A vssd1 vssd1 vccd1 vccd1 _15530_/A sky130_fd_sc_hd__inv_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19296_ _19288_/X _19295_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19296_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18247_ _18454_/A _18596_/A vssd1 vssd1 vccd1 vccd1 _18248_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15459_ _15459_/A _15459_/B vssd1 vssd1 vccd1 vccd1 _15466_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18178_ _18535_/A _18178_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _18178_/X sky130_fd_sc_hd__and3_1
XFILLER_0_142_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold503 hold503/A vssd1 vssd1 vccd1 vccd1 hold503/X sky130_fd_sc_hd__dlygate4sd3_1
X_17129_ _19244_/A _17129_/B vssd1 vssd1 vccd1 vccd1 _17470_/A sky130_fd_sc_hd__xor2_4
Xhold514 hold514/A vssd1 vssd1 vccd1 vccd1 hold514/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold525 hold525/A vssd1 vssd1 vccd1 vccd1 hold525/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 hold536/A vssd1 vssd1 vccd1 vccd1 hold536/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold547 hold547/A vssd1 vssd1 vccd1 vccd1 hold547/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold558 hold558/A vssd1 vssd1 vccd1 vccd1 hold558/X sky130_fd_sc_hd__dlygate4sd3_1
X_20140_ _20148_/A _20148_/C vssd1 vssd1 vccd1 vccd1 _21418_/A sky130_fd_sc_hd__nand2_2
Xhold569 hold569/A vssd1 vssd1 vccd1 vccd1 hold569/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20071_ _20978_/C vssd1 vssd1 vccd1 vccd1 _20981_/B sky130_fd_sc_hd__inv_2
XFILLER_0_110_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 _25406_/Q vssd1 vssd1 vccd1 vccd1 _14852_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 _21332_/Y vssd1 vssd1 vccd1 vccd1 _25813_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 hold2755/X vssd1 vssd1 vccd1 vccd1 _23197_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_139_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23830_ _23830_/A vssd1 vssd1 vccd1 vccd1 _26014_/D sky130_fd_sc_hd__clkbuf_1
Xhold1236 _25753_/Q vssd1 vssd1 vccd1 vccd1 _19738_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1247 _19625_/Y vssd1 vssd1 vccd1 vccd1 _25745_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1258 _25768_/Q vssd1 vssd1 vccd1 vccd1 _19942_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 _12996_/X vssd1 vssd1 vccd1 vccd1 _25049_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23761_ _14788_/B _14797_/B _23831_/S vssd1 vssd1 vccd1 vccd1 _23762_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20973_ _20973_/A _20973_/B _20973_/C vssd1 vssd1 vccd1 vccd1 _20974_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_71_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25500_ _26341_/CLK hold756/X vssd1 vssd1 vccd1 vccd1 hold754/A sky130_fd_sc_hd__dfxtp_1
X_22712_ _16781_/B _22421_/X _22706_/X _22707_/Y _22711_/X vssd1 vssd1 vccd1 vccd1
+ _22713_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23692_ _23692_/A vssd1 vssd1 vccd1 vccd1 _25969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25431_ _26002_/CLK _25431_/D vssd1 vssd1 vccd1 vccd1 _25431_/Q sky130_fd_sc_hd__dfxtp_1
X_22643_ _25706_/Q _22642_/A _22642_/Y vssd1 vssd1 vccd1 vccd1 _22645_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25362_ _26184_/CLK hold25/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22574_ _22574_/A _22574_/B vssd1 vssd1 vccd1 vccd1 _22575_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24313_ _24313_/A vssd1 vssd1 vccd1 vccd1 _26169_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21525_ _21573_/A _21525_/B vssd1 vssd1 vccd1 vccd1 _21525_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25293_ _26249_/CLK hold253/X vssd1 vssd1 vccd1 vccd1 hold251/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24244_ _24244_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24245_/A sky130_fd_sc_hd__and2_1
XFILLER_0_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21456_ _21455_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21456_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20407_ _20409_/B vssd1 vssd1 vccd1 vccd1 _20408_/B sky130_fd_sc_hd__inv_2
XFILLER_0_114_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24175_ hold2435/X hold2157/X _24203_/S vssd1 vssd1 vccd1 vccd1 _24176_/A sky130_fd_sc_hd__mux2_1
X_21387_ _21387_/A _21387_/B _21387_/C vssd1 vssd1 vccd1 vccd1 _21388_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23126_ _26080_/Q vssd1 vssd1 vccd1 vccd1 _23127_/A sky130_fd_sc_hd__inv_2
X_20338_ _20338_/A _21089_/B _20338_/C vssd1 vssd1 vccd1 vccd1 _20339_/B sky130_fd_sc_hd__nand3_1
X_23057_ _23057_/A _23057_/B vssd1 vssd1 vccd1 vccd1 _23058_/B sky130_fd_sc_hd__nand2_1
X_20269_ _20269_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _20269_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_179_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22008_ _22008_/A _22008_/B vssd1 vssd1 vccd1 vccd1 _22008_/Y sky130_fd_sc_hd__nand2_1
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2460 _15461_/X vssd1 vssd1 vccd1 vccd1 _15463_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2471 _26048_/Q vssd1 vssd1 vccd1 vccd1 hold2471/X sky130_fd_sc_hd__dlygate4sd3_1
X_14830_ _14830_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14830_/Y sky130_fd_sc_hd__nand2_1
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2482 _24987_/Q vssd1 vssd1 vccd1 vccd1 _12676_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2493 _25430_/Q vssd1 vssd1 vccd1 vccd1 _15049_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1770 _22741_/Y vssd1 vssd1 vccd1 vccd1 _25873_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14761_ _15839_/A _14761_/B vssd1 vssd1 vccd1 vccd1 _21968_/A sky130_fd_sc_hd__nand2_1
Xhold1781 _22972_/Y vssd1 vssd1 vccd1 vccd1 _25887_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23959_ hold2293/X hold2183/X _24001_/S vssd1 vssd1 vccd1 vccd1 _23960_/A sky130_fd_sc_hd__mux2_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1792 _22690_/Y vssd1 vssd1 vccd1 vccd1 _25871_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16500_ _16500_/A vssd1 vssd1 vccd1 vccd1 _16513_/B sky130_fd_sc_hd__inv_2
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ _13760_/A hold542/X vssd1 vssd1 vccd1 vccd1 hold543/A sky130_fd_sc_hd__nand2_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14692_ _21721_/B _15543_/B vssd1 vssd1 vccd1 vccd1 _14693_/A sky130_fd_sc_hd__nand2_1
X_17480_ _17478_/X _17241_/X _17479_/X vssd1 vssd1 vccd1 vccd1 _17481_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_168_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16431_ _16429_/X _16430_/Y _16231_/A vssd1 vssd1 vccd1 vccd1 _16431_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25629_ _25716_/CLK _25629_/D vssd1 vssd1 vccd1 vccd1 _25629_/Q sky130_fd_sc_hd__dfxtp_4
X_13643_ _25738_/Q vssd1 vssd1 vccd1 vccd1 _18243_/B sky130_fd_sc_hd__inv_2
XFILLER_0_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19150_ _19136_/X _19147_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19150_/Y sky130_fd_sc_hd__o21ai_1
X_16362_ _16361_/B _16332_/A _16347_/B vssd1 vssd1 vccd1 vccd1 _16362_/X sky130_fd_sc_hd__a21o_1
X_13574_ _25727_/Q vssd1 vssd1 vccd1 vccd1 _17813_/B sky130_fd_sc_hd__inv_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18101_ _18955_/A _18101_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18102_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15313_ _15313_/A vssd1 vssd1 vccd1 vccd1 _15320_/B sky130_fd_sc_hd__inv_2
X_12525_ _12525_/A vssd1 vssd1 vccd1 vccd1 _15774_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16293_ _16676_/A _15287_/A _16292_/Y vssd1 vssd1 vccd1 vccd1 _16295_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19081_ _19081_/A _19081_/B vssd1 vssd1 vccd1 vccd1 _19081_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_136_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18032_ _18032_/A _20622_/B _18032_/C vssd1 vssd1 vccd1 vccd1 _20592_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_87_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15244_ _15244_/A vssd1 vssd1 vccd1 vccd1 _16260_/A sky130_fd_sc_hd__inv_2
XFILLER_0_152_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15175_ _15621_/A _16203_/B vssd1 vssd1 vccd1 vccd1 _16733_/A sky130_fd_sc_hd__or2_1
XFILLER_0_2_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14126_ _14236_/A hold757/X vssd1 vssd1 vccd1 vccd1 hold758/A sky130_fd_sc_hd__nand2_1
X_19983_ _19983_/A _19983_/B vssd1 vssd1 vccd1 vccd1 _19983_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_120_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18934_ _18954_/A _25772_/Q vssd1 vssd1 vccd1 vccd1 _18936_/A sky130_fd_sc_hd__nand2_1
X_14057_ _14118_/A hold796/X vssd1 vssd1 vccd1 vccd1 _14057_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13008_ _26263_/Q _25632_/Q vssd1 vssd1 vccd1 vccd1 _14446_/A sky130_fd_sc_hd__xor2_2
X_18865_ _25705_/Q vssd1 vssd1 vccd1 vccd1 _22615_/B sky130_fd_sc_hd__inv_2
XFILLER_0_98_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17816_ _17816_/A _20662_/A vssd1 vssd1 vccd1 vccd1 _18372_/A sky130_fd_sc_hd__xor2_4
X_18796_ _18796_/A _20634_/A vssd1 vssd1 vccd1 vccd1 _19024_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17747_ _17752_/B _17764_/A vssd1 vssd1 vccd1 vccd1 _17748_/A sky130_fd_sc_hd__xor2_1
X_14959_ _14959_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14959_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17678_ _17721_/B _17685_/A vssd1 vssd1 vccd1 vccd1 _17678_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19417_ _20993_/A _22006_/B _25609_/Q vssd1 vssd1 vccd1 vccd1 _20998_/C sky130_fd_sc_hd__nand3_1
X_16629_ _16629_/A _16629_/B _16629_/C vssd1 vssd1 vccd1 vccd1 _16630_/A sky130_fd_sc_hd__and3_1
XFILLER_0_9_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19348_ _19364_/B _19435_/B vssd1 vssd1 vccd1 vccd1 _19350_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19279_ _19280_/B _19280_/A vssd1 vssd1 vccd1 vccd1 _19279_/X sky130_fd_sc_hd__or2_1
XFILLER_0_14_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21310_ _26315_/Q hold527/X vssd1 vssd1 vccd1 vccd1 _21310_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22290_ _22561_/A _22290_/B vssd1 vssd1 vccd1 vccd1 _22290_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold300 hold300/A vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
X_21241_ _25874_/Q _21241_/B _21241_/C vssd1 vssd1 vccd1 vccd1 _21244_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold311 hold311/A vssd1 vssd1 vccd1 vccd1 hold311/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold322 hold322/A vssd1 vssd1 vccd1 vccd1 hold322/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 hold333/A vssd1 vssd1 vccd1 vccd1 hold333/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold344 hold344/A vssd1 vssd1 vccd1 vccd1 hold344/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 hold355/A vssd1 vssd1 vccd1 vccd1 hold355/X sky130_fd_sc_hd__dlygate4sd3_1
X_21172_ _21172_/A _21172_/B _21172_/C vssd1 vssd1 vccd1 vccd1 _21173_/B sky130_fd_sc_hd__nand3_1
Xhold366 hold366/A vssd1 vssd1 vccd1 vccd1 hold366/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 hold377/A vssd1 vssd1 vccd1 vccd1 hold377/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 hold388/A vssd1 vssd1 vccd1 vccd1 hold388/X sky130_fd_sc_hd__dlygate4sd3_1
X_20123_ _26279_/Q _20078_/X hold707/X vssd1 vssd1 vccd1 vccd1 _20126_/B sky130_fd_sc_hd__a21oi_1
Xhold399 hold399/A vssd1 vssd1 vccd1 vccd1 hold399/X sky130_fd_sc_hd__dlygate4sd3_1
X_25980_ _26073_/CLK _25980_/D vssd1 vssd1 vccd1 vccd1 _25980_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_141_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24931_ hold957/A hold972/A _24940_/S vssd1 vssd1 vccd1 vccd1 _24932_/B sky130_fd_sc_hd__mux2_1
X_20054_ _20054_/A _22120_/B vssd1 vssd1 vccd1 vccd1 _20055_/A sky130_fd_sc_hd__nand2_1
Xhold1000 _16268_/Y vssd1 vssd1 vccd1 vccd1 _25507_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 _25071_/Q vssd1 vssd1 vccd1 vccd1 _18058_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1022 _13302_/X vssd1 vssd1 vccd1 vccd1 _25102_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 _25068_/Q vssd1 vssd1 vccd1 vccd1 _17914_/B sky130_fd_sc_hd__dlygate4sd3_1
X_24862_ _24860_/X _24861_/X _24946_/A vssd1 vssd1 vccd1 vccd1 _24862_/X sky130_fd_sc_hd__mux2_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1044 _12865_/X vssd1 vssd1 vccd1 vccd1 _25024_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1055 _25763_/Q vssd1 vssd1 vccd1 vccd1 _19878_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1066 _13452_/X vssd1 vssd1 vccd1 vccd1 _25127_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23813_ _23813_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23814_/A sky130_fd_sc_hd__and2_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1077 _25716_/Q vssd1 vssd1 vccd1 vccd1 _19214_/B sky130_fd_sc_hd__dlygate4sd3_1
X_24793_ hold2508/X _26326_/Q _24817_/S vssd1 vssd1 vccd1 vccd1 _24793_/X sky130_fd_sc_hd__mux2_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1088 _13370_/X vssd1 vssd1 vccd1 vccd1 _25113_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 _25568_/Q vssd1 vssd1 vccd1 vccd1 _16900_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23744_ _23744_/A vssd1 vssd1 vccd1 vccd1 _25986_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20956_ _26302_/Q hold437/X vssd1 vssd1 vccd1 vccd1 _20956_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23675_ _23675_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23676_/A sky130_fd_sc_hd__and2_1
XFILLER_0_36_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20887_ _20889_/B _20889_/C vssd1 vssd1 vccd1 vccd1 _20888_/A sky130_fd_sc_hd__nand2_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25414_ _25859_/CLK _25414_/D vssd1 vssd1 vccd1 vccd1 _25414_/Q sky130_fd_sc_hd__dfxtp_1
X_22626_ _22626_/A _22626_/B vssd1 vssd1 vccd1 vccd1 _22627_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_181_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25345_ _26171_/CLK hold376/X vssd1 vssd1 vccd1 vccd1 hold374/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22557_ _22557_/A _23001_/B _22557_/C vssd1 vssd1 vccd1 vccd1 _22557_/X sky130_fd_sc_hd__and3_1
XFILLER_0_106_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21508_ _21508_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21508_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_122_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25276_ _26109_/CLK hold247/X vssd1 vssd1 vccd1 vccd1 hold245/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13290_ _26312_/Q _19532_/A vssd1 vssd1 vccd1 vccd1 _14602_/A sky130_fd_sc_hd__xor2_1
X_22488_ _25828_/Q _22488_/B vssd1 vssd1 vccd1 vccd1 _22488_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_51_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24227_ _24227_/A vssd1 vssd1 vccd1 vccd1 _26141_/D sky130_fd_sc_hd__clkbuf_1
X_21439_ _26323_/Q hold647/X vssd1 vssd1 vccd1 vccd1 _21439_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_146_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24158_ _24158_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24159_/A sky130_fd_sc_hd__and2_1
X_23109_ _15724_/B _22893_/A _22829_/X vssd1 vssd1 vccd1 vccd1 _23109_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16980_ _16980_/A _25580_/Q vssd1 vssd1 vccd1 vccd1 _16980_/Y sky130_fd_sc_hd__nand2_1
X_24089_ hold1832/X _26097_/Q _24126_/S vssd1 vssd1 vccd1 vccd1 _24089_/X sky130_fd_sc_hd__mux2_1
X_15931_ _15932_/B _15932_/A vssd1 vssd1 vccd1 vccd1 _15933_/A sky130_fd_sc_hd__or2_1
XFILLER_0_120_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18650_ _18650_/A _25822_/Q _18650_/C vssd1 vssd1 vccd1 vccd1 _20370_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_189_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15862_ _15860_/X hold693/X _15805_/X vssd1 vssd1 vccd1 vccd1 hold694/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2290 _15047_/Y vssd1 vssd1 vccd1 vccd1 _25429_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17601_ _17601_/A _17601_/B vssd1 vssd1 vccd1 vccd1 _17601_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_189_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14813_ _14900_/A _14813_/B vssd1 vssd1 vccd1 vccd1 _14813_/Y sky130_fd_sc_hd__nand2_1
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18581_ _18579_/Y _18580_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25673_/D sky130_fd_sc_hd__a21oi_1
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ _23175_/B _15793_/B vssd1 vssd1 vccd1 vccd1 _23172_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_87_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17532_ _17605_/A _17532_/B vssd1 vssd1 vccd1 vccd1 _17532_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_93_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ _14750_/B _21900_/A vssd1 vssd1 vccd1 vccd1 _21899_/B sky130_fd_sc_hd__xnor2_2
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17463_ _17463_/A _17463_/B vssd1 vssd1 vccd1 vccd1 _17463_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_156_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14675_ _14675_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _14675_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_184_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19202_ _26219_/Q hold739/X vssd1 vssd1 vccd1 vccd1 _19202_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16414_ _16441_/A _16414_/B vssd1 vssd1 vccd1 vccd1 _16439_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_104_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13626_ _18172_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13626_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_67_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17394_ _17392_/X _17241_/X _17393_/X vssd1 vssd1 vccd1 vccd1 _17395_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_55_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19133_ _22786_/A vssd1 vssd1 vccd1 vccd1 _23195_/B sky130_fd_sc_hd__buf_8
XFILLER_0_109_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16345_ _16346_/A _16691_/B hold968/X vssd1 vssd1 vccd1 vccd1 _16347_/A sky130_fd_sc_hd__a21oi_1
X_13557_ _26227_/Q _13426_/X _13468_/X _13556_/Y vssd1 vssd1 vccd1 vccd1 _13558_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12508_ hold868/A _24974_/Q _24973_/Q _24972_/Q vssd1 vssd1 vccd1 vccd1 _12515_/A
+ sky130_fd_sc_hd__or4_1
X_19064_ _19186_/A _19064_/B vssd1 vssd1 vccd1 vccd1 _19064_/Y sky130_fd_sc_hd__nand2_1
X_16276_ _16276_/A _16276_/B vssd1 vssd1 vccd1 vccd1 _16276_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_125_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13488_ _17927_/B _13518_/B vssd1 vssd1 vccd1 vccd1 _13488_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18015_ _21924_/A _25587_/Q vssd1 vssd1 vccd1 vccd1 _18017_/B sky130_fd_sc_hd__nand2_1
X_15227_ _15795_/A _16248_/B vssd1 vssd1 vccd1 vccd1 _15230_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_140_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15158_ _15158_/A vssd1 vssd1 vccd1 vccd1 _15160_/A sky130_fd_sc_hd__inv_2
XFILLER_0_10_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14109_ _26315_/Q _13988_/X _13981_/X _14108_/Y vssd1 vssd1 vccd1 vccd1 _14110_/B
+ sky130_fd_sc_hd__a22o_1
X_15089_ _15089_/A _15106_/A vssd1 vssd1 vccd1 vccd1 _15089_/Y sky130_fd_sc_hd__nand2_1
X_19966_ _26274_/Q hold680/X vssd1 vssd1 vccd1 vccd1 _19966_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18917_ _18917_/A _19999_/A vssd1 vssd1 vccd1 vccd1 _19066_/B sky130_fd_sc_hd__xor2_4
X_19897_ _19999_/A _22665_/B _25643_/Q vssd1 vssd1 vccd1 vccd1 _20004_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18848_ _25896_/Q _22589_/A vssd1 vssd1 vccd1 vccd1 _18856_/A sky130_fd_sc_hd__or2_2
XFILLER_0_101_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18779_ _19026_/A _18779_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18779_/X sky130_fd_sc_hd__and3_1
XFILLER_0_179_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20810_ _26297_/Q hold623/X vssd1 vssd1 vccd1 vccd1 _20810_/Y sky130_fd_sc_hd__nand2_1
X_21790_ _21787_/X _21788_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _21790_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_166_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20741_ _20741_/A _20741_/B vssd1 vssd1 vccd1 vccd1 _20745_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_187_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23460_ _24956_/S hold113/A _23459_/X vssd1 vssd1 vccd1 vccd1 _23460_/Y sky130_fd_sc_hd__o21ai_1
X_20672_ _20672_/A _22539_/B vssd1 vssd1 vccd1 vccd1 _20673_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_175_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22411_ _19758_/A _22410_/A _22410_/Y vssd1 vssd1 vccd1 vccd1 _22413_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23391_ _23391_/A vssd1 vssd1 vccd1 vccd1 _24940_/S sky130_fd_sc_hd__buf_12
XFILLER_0_174_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_clk _25759_/CLK vssd1 vssd1 vccd1 vccd1 _25898_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25130_ _25711_/CLK hold454/X vssd1 vssd1 vccd1 vccd1 hold452/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22342_ _22340_/Y _22341_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _22342_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25061_ _26142_/CLK _25061_/D vssd1 vssd1 vccd1 vccd1 _25061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22273_ _22273_/A _22273_/B vssd1 vssd1 vccd1 vccd1 _22890_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_143_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24012_ _24012_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24013_/A sky130_fd_sc_hd__and2_1
XFILLER_0_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold130 hold130/A vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
X_21224_ _21659_/C _21610_/C vssd1 vssd1 vccd1 vccd1 _21225_/C sky130_fd_sc_hd__nand2_1
Xhold141 hold141/A vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold152 hold152/A vssd1 vssd1 vccd1 vccd1 hold152/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 hold163/A vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 hold174/A vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21155_ _21153_/Y _21154_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21155_/Y sky130_fd_sc_hd__a21oi_1
Xhold185 hold185/A vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 hold196/A vssd1 vssd1 vccd1 vccd1 hold196/X sky130_fd_sc_hd__dlygate4sd3_1
X_20106_ _20106_/A _20106_/B _20106_/C vssd1 vssd1 vccd1 vccd1 _20107_/B sky130_fd_sc_hd__nand3_1
X_25963_ _26042_/CLK _25963_/D vssd1 vssd1 vccd1 vccd1 _25963_/Q sky130_fd_sc_hd__dfxtp_1
X_21086_ _21086_/A _21086_/B _21086_/C vssd1 vssd1 vccd1 vccd1 _21090_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_42_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_97_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _25998_/CLK sky130_fd_sc_hd__clkbuf_16
X_24914_ _24946_/A _24914_/B vssd1 vssd1 vccd1 vccd1 _24914_/Y sky130_fd_sc_hd__nor2_1
X_20037_ _20036_/Y _21228_/A _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20037_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25894_ _25895_/CLK _25894_/D vssd1 vssd1 vccd1 vccd1 _25894_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24845_ _15263_/A _15290_/B _24860_/S vssd1 vssd1 vccd1 vccd1 _24845_/X sky130_fd_sc_hd__mux2_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ hold1/X _12748_/X _12789_/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__a21o_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21988_ _23167_/A _22729_/A vssd1 vssd1 vccd1 vccd1 _21996_/A sky130_fd_sc_hd__nand2_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24776_ _24776_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24777_/A sky130_fd_sc_hd__and2_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23727_ _25980_/Q hold2161/X _23754_/S vssd1 vssd1 vccd1 vccd1 _23727_/X sky130_fd_sc_hd__mux2_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20939_ _22485_/B vssd1 vssd1 vccd1 vccd1 _21943_/B sky130_fd_sc_hd__inv_2
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _14458_/Y hold225/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold226/A sky130_fd_sc_hd__a21oi_1
X_23658_ _23658_/A vssd1 vssd1 vccd1 vccd1 _25958_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13411_ hold973/X _13944_/A vssd1 vssd1 vccd1 vccd1 _13411_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22609_ _16757_/B _22421_/X _22603_/X _22604_/Y _22608_/X vssd1 vssd1 vccd1 vccd1
+ _22610_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14391_ _14391_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14391_/Y sky130_fd_sc_hd__nand2_1
X_23589_ hold832/X _25918_/Q hold829/X _25916_/Q vssd1 vssd1 vccd1 vccd1 _23590_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_153_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _25650_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_52_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16130_ _16128_/X hold645/X _16076_/X vssd1 vssd1 vccd1 vccd1 hold646/A sky130_fd_sc_hd__a21oi_1
X_13342_ _26320_/Q _19644_/A vssd1 vssd1 vccd1 vccd1 _14626_/A sky130_fd_sc_hd__xor2_1
X_25328_ _26152_/CLK hold136/X vssd1 vssd1 vccd1 vccd1 hold134/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16061_ _16062_/B _16160_/A vssd1 vssd1 vccd1 vccd1 _16063_/A sky130_fd_sc_hd__or2_1
X_13273_ _13220_/X _14593_/A _13242_/X _19488_/A vssd1 vssd1 vccd1 vccd1 _13273_/X
+ sky130_fd_sc_hd__a22o_1
X_25259_ _26046_/CLK _25259_/D vssd1 vssd1 vccd1 vccd1 _25259_/Q sky130_fd_sc_hd__dfxtp_1
X_15012_ _22173_/B _15778_/B _15013_/B vssd1 vssd1 vccd1 vccd1 _15014_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_20_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19820_ _19821_/B _19821_/A vssd1 vssd1 vccd1 vccd1 _19820_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19751_ _19743_/X _19750_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19751_/Y sky130_fd_sc_hd__o21ai_1
X_16963_ _16977_/A _16963_/B vssd1 vssd1 vccd1 vccd1 _16963_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_88_clk clkbuf_leaf_95_clk/A vssd1 vssd1 vccd1 vccd1 _26052_/CLK sky130_fd_sc_hd__clkbuf_16
X_18702_ _18986_/A _19504_/A vssd1 vssd1 vccd1 vccd1 _18702_/Y sky130_fd_sc_hd__nand2_1
X_15914_ _15912_/X _15913_/Y _15805_/X vssd1 vssd1 vccd1 vccd1 hold859/A sky130_fd_sc_hd__a21oi_1
X_19682_ _19680_/Y _19681_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19682_/Y sky130_fd_sc_hd__a21oi_1
X_16894_ _16892_/Y _16893_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16894_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18633_ _18633_/A _18633_/B _18633_/C vssd1 vssd1 vccd1 vccd1 _22329_/A sky130_fd_sc_hd__nand3_2
X_15845_ _15857_/B _15845_/B vssd1 vssd1 vccd1 vccd1 _15869_/B sky130_fd_sc_hd__nand2_1
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18564_ _20200_/B _19659_/A vssd1 vssd1 vccd1 vccd1 _18565_/B sky130_fd_sc_hd__nand2_1
X_15776_ _23156_/B _15776_/B vssd1 vssd1 vccd1 vccd1 _15777_/A sky130_fd_sc_hd__nand2_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _12891_/X _14434_/A _12909_/X _25628_/Q vssd1 vssd1 vccd1 vccd1 _12988_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_188_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17515_ _17513_/X _17241_/X _17514_/X vssd1 vssd1 vccd1 vccd1 _17516_/A sky130_fd_sc_hd__a21o_1
X_14727_ _14727_/A vssd1 vssd1 vccd1 vccd1 _14923_/A sky130_fd_sc_hd__inv_2
XFILLER_0_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18495_ _18535_/A _18495_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18495_/X sky130_fd_sc_hd__and3_1
XFILLER_0_28_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17446_ _17444_/Y _17445_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _17446_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14658_ _14688_/A hold41/X vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__nand2_1
XFILLER_0_157_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13609_ _13703_/A _13609_/B vssd1 vssd1 vccd1 vccd1 _13609_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_156_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17377_ _17375_/Y _17376_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _17377_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14589_ _14589_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14589_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_clk _25184_/CLK vssd1 vssd1 vccd1 vccd1 _26252_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_172_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19116_ _19115_/C _17873_/B _20113_/A vssd1 vssd1 vccd1 vccd1 _19961_/B sky130_fd_sc_hd__a21boi_4
X_16328_ hold906/X vssd1 vssd1 vccd1 vccd1 _16331_/B sky130_fd_sc_hd__inv_2
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19047_ _19082_/A _19047_/B _22786_/A vssd1 vssd1 vccd1 vccd1 _19047_/X sky130_fd_sc_hd__and3_1
XFILLER_0_3_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16259_ hold999/X vssd1 vssd1 vccd1 vccd1 _16262_/B sky130_fd_sc_hd__inv_2
XFILLER_0_129_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19949_ _19950_/B _19950_/A vssd1 vssd1 vccd1 vccd1 _19949_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_79_clk clkbuf_leaf_82_clk/A vssd1 vssd1 vccd1 vccd1 _25864_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22960_ _22960_/A _22960_/B vssd1 vssd1 vccd1 vccd1 _22961_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_156_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21911_ _23136_/A vssd1 vssd1 vccd1 vccd1 _23135_/A sky130_fd_sc_hd__inv_2
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22891_ _22891_/A _22891_/B vssd1 vssd1 vccd1 vccd1 _22892_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21842_ _23104_/A vssd1 vssd1 vccd1 vccd1 _23103_/A sky130_fd_sc_hd__inv_2
X_24630_ hold2735/X hold2733/X _24664_/S vssd1 vssd1 vccd1 vccd1 _24631_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_78_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24561_ _24561_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24562_/A sky130_fd_sc_hd__and2_1
X_21773_ _25803_/Q _21773_/B vssd1 vssd1 vccd1 vccd1 _21773_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_93_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26300_ _26303_/CLK _26300_/D vssd1 vssd1 vccd1 vccd1 _26300_/Q sky130_fd_sc_hd__dfxtp_2
X_23512_ _24944_/S hold344/A _23511_/X vssd1 vssd1 vccd1 vccd1 _23512_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20724_ _21660_/B _21387_/B vssd1 vssd1 vccd1 vccd1 _20725_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_110_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24492_ hold2630/X hold2600/X _24510_/S vssd1 vssd1 vccd1 vccd1 _24493_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_147_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26231_ _26231_/CLK _26231_/D vssd1 vssd1 vccd1 vccd1 _26231_/Q sky130_fd_sc_hd__dfxtp_2
X_23443_ _24922_/S hold407/A _23442_/X vssd1 vssd1 vccd1 vccd1 _23443_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_163_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20655_ _26293_/Q hold638/X vssd1 vssd1 vccd1 vccd1 _20655_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23374_ _23374_/A vssd1 vssd1 vccd1 vccd1 _25937_/D sky130_fd_sc_hd__clkbuf_1
X_26162_ _26289_/CLK _26162_/D vssd1 vssd1 vccd1 vccd1 _26162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20586_ _20586_/A _20586_/B vssd1 vssd1 vccd1 vccd1 _20590_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22325_ _22325_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _22325_/X sky130_fd_sc_hd__and2_1
X_25113_ _26325_/CLK _25113_/D vssd1 vssd1 vccd1 vccd1 _25113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26093_ _26093_/CLK _26093_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25044_ _26130_/CLK _25044_/D vssd1 vssd1 vccd1 vccd1 _25044_/Q sky130_fd_sc_hd__dfxtp_1
X_22256_ _22257_/A _22257_/C _23154_/A vssd1 vssd1 vccd1 vccd1 _22256_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_104_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21207_ _21207_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21207_/Y sky130_fd_sc_hd__nand2_1
X_22187_ _22187_/A _22841_/A vssd1 vssd1 vccd1 vccd1 _22198_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21138_ _21561_/C _21610_/C vssd1 vssd1 vccd1 vccd1 _21141_/A sky130_fd_sc_hd__nand2_1
X_25946_ _26009_/CLK _25946_/D vssd1 vssd1 vccd1 vccd1 _25946_/Q sky130_fd_sc_hd__dfxtp_1
X_13960_ _14061_/A _13960_/B vssd1 vssd1 vccd1 vccd1 _13960_/Y sky130_fd_sc_hd__nand2_1
X_21069_ _21636_/A _21069_/B _21068_/X vssd1 vssd1 vccd1 vccd1 _21070_/B sky130_fd_sc_hd__or3b_1
X_12911_ _26116_/Q _12907_/X _12910_/X vssd1 vssd1 vccd1 vccd1 _12911_/X sky130_fd_sc_hd__a21o_1
X_25877_ _25877_/CLK _25877_/D vssd1 vssd1 vccd1 vccd1 _25877_/Q sky130_fd_sc_hd__dfxtp_2
X_13891_ _26280_/Q _13801_/X _13793_/X _13890_/Y vssd1 vssd1 vccd1 vccd1 _13892_/B
+ sky130_fd_sc_hd__a22o_1
X_15630_ _15628_/Y _15629_/Y _15464_/X vssd1 vssd1 vccd1 vccd1 hold947/A sky130_fd_sc_hd__a21oi_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24828_ _24828_/A vssd1 vssd1 vccd1 vccd1 _26337_/D sky130_fd_sc_hd__clkbuf_1
X_12842_ _12726_/B _14343_/A _12752_/X _25600_/Q vssd1 vssd1 vccd1 vccd1 _12842_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _15559_/X _15560_/Y _15464_/X vssd1 vssd1 vccd1 vccd1 _15561_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12773_ _26218_/Q _25587_/Q vssd1 vssd1 vccd1 vccd1 _14304_/A sky130_fd_sc_hd__xor2_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24759_ _24759_/A vssd1 vssd1 vccd1 vccd1 _26314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _17298_/Y _17299_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _17300_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14512_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14512_/Y sky130_fd_sc_hd__nand2_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18280_ _25868_/Q _21809_/A vssd1 vssd1 vccd1 vccd1 _18290_/A sky130_fd_sc_hd__or2_2
X_15492_ _15492_/A vssd1 vssd1 vccd1 vccd1 _16451_/A sky130_fd_sc_hd__inv_2
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17231_ _17229_/Y _17230_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _17231_/Y sky130_fd_sc_hd__a21oi_1
X_14443_ _14443_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14443_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_83_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17162_ _17160_/X _23187_/B _17161_/X vssd1 vssd1 vccd1 vccd1 _17163_/A sky130_fd_sc_hd__a21o_1
X_14374_ _14404_/A hold86/X vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16113_ _16113_/A _16113_/B vssd1 vssd1 vccd1 vccd1 _16114_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_181_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13325_ _26189_/Q _13239_/X _13324_/X vssd1 vssd1 vccd1 vccd1 _13325_/X sky130_fd_sc_hd__a21o_1
X_17093_ _17393_/A _25007_/Q _19994_/B vssd1 vssd1 vccd1 vccd1 _17093_/X sky130_fd_sc_hd__and3_1
XFILLER_0_12_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16044_ _16212_/A hold704/X vssd1 vssd1 vccd1 vccd1 hold705/A sky130_fd_sc_hd__nand2_1
X_13256_ _26178_/Q _13239_/X _13255_/X vssd1 vssd1 vccd1 vccd1 _13256_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_0_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13187_ _13109_/X _13185_/X _13096_/X _13186_/X vssd1 vssd1 vccd1 vccd1 _13187_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19803_ _20596_/A _22488_/B _25636_/Q vssd1 vssd1 vccd1 vccd1 _20601_/C sky130_fd_sc_hd__nand3_1
X_17995_ _20818_/B _19331_/A vssd1 vssd1 vccd1 vccd1 _17996_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_159_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16946_ _16946_/A _16946_/B vssd1 vssd1 vccd1 vccd1 _16946_/Y sky130_fd_sc_hd__nand2_1
X_19734_ _19734_/A _19734_/B vssd1 vssd1 vccd1 vccd1 _19734_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_1_clk _26093_/CLK vssd1 vssd1 vccd1 vccd1 _26216_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19665_ _19663_/X _19664_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19665_/Y sky130_fd_sc_hd__a21oi_1
X_16877_ _16875_/X _16711_/X _16876_/Y _25886_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16878_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_56_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18616_ _18818_/A _18960_/A vssd1 vssd1 vccd1 vccd1 _18617_/B sky130_fd_sc_hd__xnor2_2
X_15828_ _15828_/A vssd1 vssd1 vccd1 vccd1 _15828_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_172_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19596_ _19723_/A _19596_/B vssd1 vssd1 vccd1 vccd1 _19596_/Y sky130_fd_sc_hd__nand2_1
X_18547_ _18793_/A _19738_/B _18894_/C vssd1 vssd1 vccd1 vccd1 _18548_/C sky130_fd_sc_hd__nand3_1
X_15759_ _15761_/B _16960_/A vssd1 vssd1 vccd1 vccd1 _15760_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_87_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18478_ _18641_/A _19345_/A vssd1 vssd1 vccd1 vccd1 _18478_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17429_ _17426_/Y _17427_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _17429_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20440_ _20443_/A _20443_/C vssd1 vssd1 vccd1 vccd1 _20441_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20371_ _20371_/A _20371_/B vssd1 vssd1 vccd1 vccd1 _21515_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_67_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22110_ _22110_/A _23074_/A _22110_/C vssd1 vssd1 vccd1 vccd1 _22110_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_67_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23090_ _23090_/A _23090_/B vssd1 vssd1 vccd1 vccd1 _23091_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22041_ _18432_/A _25811_/Q _22039_/Y _22040_/Y vssd1 vssd1 vccd1 vccd1 _22042_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25800_ _25803_/CLK _25800_/D vssd1 vssd1 vccd1 vccd1 _25800_/Q sky130_fd_sc_hd__dfxtp_1
X_23992_ hold2053/X _26066_/Q _24001_/S vssd1 vssd1 vccd1 vccd1 _23992_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_98_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25731_ _25784_/CLK _25731_/D vssd1 vssd1 vccd1 vccd1 _25731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22943_ _22943_/A _22943_/B vssd1 vssd1 vccd1 vccd1 _22944_/A sky130_fd_sc_hd__xor2_1
X_25662_ _26164_/CLK _25662_/D vssd1 vssd1 vccd1 vccd1 _25662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22874_ _23183_/B _22874_/B vssd1 vssd1 vccd1 vccd1 _22876_/A sky130_fd_sc_hd__nand2_1
X_24613_ _24613_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24614_/A sky130_fd_sc_hd__and2_1
X_21825_ _21825_/A _21825_/B _22926_/A vssd1 vssd1 vccd1 vccd1 _21825_/Y sky130_fd_sc_hd__nand3_1
X_25593_ _26112_/CLK _25593_/D vssd1 vssd1 vccd1 vccd1 _25593_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21756_ _21727_/X _21755_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _21756_/Y sky130_fd_sc_hd__o21ai_1
X_24544_ hold2732/X hold2647/X _24587_/S vssd1 vssd1 vccd1 vccd1 _24545_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_47_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20707_ _20707_/A _20707_/B vssd1 vssd1 vccd1 vccd1 _20709_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_136_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24475_ _24475_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24476_/A sky130_fd_sc_hd__and2_1
X_21687_ _22058_/A _21687_/B vssd1 vssd1 vccd1 vccd1 _21687_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26214_ _26216_/CLK _26214_/D vssd1 vssd1 vccd1 vccd1 _26214_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_62_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20638_ _23069_/B vssd1 vssd1 vccd1 vccd1 _22518_/B sky130_fd_sc_hd__inv_2
X_23426_ _24940_/S hold395/A _23425_/X vssd1 vssd1 vccd1 vccd1 _23426_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23357_ _23360_/A _23377_/B _23357_/C vssd1 vssd1 vccd1 vccd1 _23358_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_61_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26145_ _26146_/CLK _26145_/D vssd1 vssd1 vccd1 vccd1 _26145_/Q sky130_fd_sc_hd__dfxtp_1
X_20569_ _21596_/A vssd1 vssd1 vccd1 vccd1 _21595_/A sky130_fd_sc_hd__inv_2
XFILLER_0_85_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22308_ _25792_/Q _22308_/B vssd1 vssd1 vccd1 vccd1 _22308_/Y sky130_fd_sc_hd__nor2_1
X_13110_ _26282_/Q _25651_/Q vssd1 vssd1 vccd1 vccd1 _14506_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_104_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14090_ _18388_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14090_/Y sky130_fd_sc_hd__nor2_1
X_23288_ _23288_/A vssd1 vssd1 vccd1 vccd1 _25920_/D sky130_fd_sc_hd__clkbuf_1
X_26076_ _26079_/CLK _26076_/D vssd1 vssd1 vccd1 vccd1 _26076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ _26141_/Q _12907_/X _13040_/X vssd1 vssd1 vccd1 vccd1 _13041_/X sky130_fd_sc_hd__a21o_1
X_25027_ _26112_/CLK _25027_/D vssd1 vssd1 vccd1 vccd1 _25027_/Q sky130_fd_sc_hd__dfxtp_1
X_22239_ _22239_/A _22239_/B vssd1 vssd1 vccd1 vccd1 _22239_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16800_ _16798_/Y _16799_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16800_/Y sky130_fd_sc_hd__a21oi_1
X_17780_ _17780_/A _17780_/B vssd1 vssd1 vccd1 vccd1 _17781_/B sky130_fd_sc_hd__nand2_1
X_14992_ _14998_/B _14993_/A vssd1 vssd1 vccd1 vccd1 _14992_/X sky130_fd_sc_hd__or2_1
X_16731_ _16980_/A _16736_/B vssd1 vssd1 vccd1 vccd1 _16733_/B sky130_fd_sc_hd__nand2_1
X_25929_ _25939_/CLK hold954/X vssd1 vssd1 vccd1 vccd1 hold952/A sky130_fd_sc_hd__dfxtp_1
X_13943_ _14000_/A hold742/X vssd1 vssd1 vccd1 vccd1 hold743/A sky130_fd_sc_hd__nand2_1
XFILLER_0_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19450_ _19448_/X _19449_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19450_/Y sky130_fd_sc_hd__a21oi_1
X_16662_ _16698_/A hold942/X vssd1 vssd1 vccd1 vccd1 _16662_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13874_ _13880_/A hold602/X vssd1 vssd1 vccd1 vccd1 hold603/A sky130_fd_sc_hd__nand2_1
X_18401_ _18401_/A _18401_/B vssd1 vssd1 vccd1 vccd1 _22014_/A sky130_fd_sc_hd__nand2_1
X_15613_ _15612_/B _15590_/B _15605_/B vssd1 vssd1 vccd1 vccd1 _15613_/Y sky130_fd_sc_hd__a21oi_1
X_12825_ _12726_/B _14334_/A _12752_/X _25597_/Q vssd1 vssd1 vccd1 vccd1 _12825_/X
+ sky130_fd_sc_hd__a22o_1
X_19381_ _19452_/A _19381_/B vssd1 vssd1 vccd1 vccd1 _19381_/Y sky130_fd_sc_hd__nand2_1
X_16593_ _16698_/A hold962/X vssd1 vssd1 vccd1 vccd1 _16593_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18332_ _19073_/A _18332_/B vssd1 vssd1 vccd1 vccd1 _18332_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_55_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15544_ _16876_/A vssd1 vssd1 vccd1 vccd1 _15546_/A sky130_fd_sc_hd__inv_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _17029_/B _14264_/A vssd1 vssd1 vccd1 vccd1 _12756_/X sky130_fd_sc_hd__or2_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18263_ _18446_/A _18263_/B _18952_/C vssd1 vssd1 vccd1 vccd1 _18264_/C sky130_fd_sc_hd__nand3_1
X_15475_ _22879_/B _16369_/B vssd1 vssd1 vccd1 vccd1 _16435_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_127_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12687_ _12687_/A _24836_/B _12700_/B vssd1 vssd1 vccd1 vccd1 _12688_/A sky130_fd_sc_hd__and3_1
XFILLER_0_154_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17214_ _17393_/A _17214_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17214_/X sky130_fd_sc_hd__and3_1
XFILLER_0_53_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14426_ _14465_/A hold215/X vssd1 vssd1 vccd1 vccd1 hold216/A sky130_fd_sc_hd__nand2_1
XFILLER_0_86_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18194_ _21972_/B _25608_/Q vssd1 vssd1 vccd1 vccd1 _18196_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17145_ _19744_/A _17145_/B vssd1 vssd1 vccd1 vccd1 _17555_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_53_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14357_ _14355_/Y hold255/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold256/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold707 hold707/A vssd1 vssd1 vccd1 vccd1 hold707/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold718 hold718/A vssd1 vssd1 vccd1 vccd1 hold718/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13308_ _13207_/X _13306_/X _13300_/X _13307_/X vssd1 vssd1 vccd1 vccd1 _13308_/X
+ sky130_fd_sc_hd__o211a_1
Xhold729 hold729/A vssd1 vssd1 vccd1 vccd1 hold729/X sky130_fd_sc_hd__dlygate4sd3_1
X_17076_ _17638_/A _17076_/B vssd1 vssd1 vccd1 vccd1 _17076_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_126_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14288_ _14590_/A vssd1 vssd1 vccd1 vccd1 _14688_/A sky130_fd_sc_hd__buf_8
XFILLER_0_110_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16027_ _16027_/A _16027_/B vssd1 vssd1 vccd1 vccd1 _16028_/A sky130_fd_sc_hd__or2_1
X_13239_ _14262_/B vssd1 vssd1 vccd1 vccd1 _13239_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2108 _12692_/X vssd1 vssd1 vccd1 vccd1 _12693_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2119 _26017_/Q vssd1 vssd1 vccd1 vccd1 hold2119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1407 _25401_/Q vssd1 vssd1 vccd1 vccd1 _14813_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_97_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1418 _14874_/Y vssd1 vssd1 vccd1 vccd1 _25408_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17978_ _17978_/A _19159_/A vssd1 vssd1 vccd1 vccd1 _19046_/A sky130_fd_sc_hd__xor2_4
Xhold1429 _25797_/Q vssd1 vssd1 vccd1 vccd1 _20906_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16929_ _16930_/B _16930_/A vssd1 vssd1 vccd1 vccd1 _16929_/X sky130_fd_sc_hd__or2_1
X_19717_ _20361_/A _19715_/Y _20366_/C vssd1 vssd1 vccd1 vccd1 _19807_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19648_ _19649_/B _19649_/A vssd1 vssd1 vccd1 vccd1 _19648_/X sky130_fd_sc_hd__or2_1
XFILLER_0_172_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19579_ _19579_/A _19579_/B vssd1 vssd1 vccd1 vccd1 _19579_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_133_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21610_ _21610_/A _21610_/B _21610_/C vssd1 vssd1 vccd1 vccd1 _21614_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_153_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22590_ _25832_/Q _22590_/B vssd1 vssd1 vccd1 vccd1 _22590_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_75_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21541_ _21573_/A _21541_/B vssd1 vssd1 vccd1 vccd1 _21541_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24260_ _24260_/A vssd1 vssd1 vccd1 vccd1 _26152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21472_ _21471_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21472_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23211_ _23211_/A _23211_/B vssd1 vssd1 vccd1 vccd1 _23211_/X sky130_fd_sc_hd__xor2_1
X_20423_ _21042_/A _20423_/B _20422_/X vssd1 vssd1 vccd1 vccd1 _20424_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_126_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24191_ _24560_/A vssd1 vssd1 vccd1 vccd1 _24280_/B sky130_fd_sc_hd__buf_8
XFILLER_0_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23142_ _26081_/Q vssd1 vssd1 vccd1 vccd1 _23143_/A sky130_fd_sc_hd__inv_2
X_20354_ _20354_/A _20354_/B _20354_/C vssd1 vssd1 vccd1 vccd1 _20358_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_113_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23073_ _23073_/A _23073_/B vssd1 vssd1 vccd1 vccd1 _23074_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20285_ _20285_/A _20285_/B vssd1 vssd1 vccd1 vccd1 _20288_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22024_ _22743_/A _23184_/A vssd1 vssd1 vccd1 vccd1 _22030_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_80_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2620 _26280_/Q vssd1 vssd1 vccd1 vccd1 hold2620/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2631 _24970_/Q vssd1 vssd1 vccd1 vccd1 _12585_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2642 _26246_/Q vssd1 vssd1 vccd1 vccd1 hold2642/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2653 _26225_/Q vssd1 vssd1 vccd1 vccd1 hold2653/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2664 _26252_/Q vssd1 vssd1 vccd1 vccd1 hold2664/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2675 _26288_/Q vssd1 vssd1 vccd1 vccd1 hold2675/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1930 _26133_/Q vssd1 vssd1 vccd1 vccd1 hold1930/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1941 _14279_/Y vssd1 vssd1 vccd1 vccd1 hold1941/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2686 _26298_/Q vssd1 vssd1 vccd1 vccd1 hold2686/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1952 _15034_/B vssd1 vssd1 vccd1 vccd1 _15024_/B sky130_fd_sc_hd__dlygate4sd3_1
X_23975_ _23975_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23976_/A sky130_fd_sc_hd__and2_1
Xhold2697 _24541_/X vssd1 vssd1 vccd1 vccd1 _24542_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1963 _26038_/Q vssd1 vssd1 vccd1 vccd1 hold1963/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1974 _25967_/Q vssd1 vssd1 vccd1 vccd1 hold1974/X sky130_fd_sc_hd__dlygate4sd3_1
X_25714_ _25716_/CLK hold820/X vssd1 vssd1 vccd1 vccd1 hold818/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22926_ _22926_/A _22926_/B vssd1 vssd1 vccd1 vccd1 _22927_/A sky130_fd_sc_hd__xor2_1
Xhold1985 _26157_/Q vssd1 vssd1 vccd1 vccd1 hold1985/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1996 _24258_/X vssd1 vssd1 vccd1 vccd1 _24259_/A sky130_fd_sc_hd__dlygate4sd3_1
X_25645_ _25712_/CLK _25645_/D vssd1 vssd1 vccd1 vccd1 _25645_/Q sky130_fd_sc_hd__dfxtp_4
X_22857_ _22854_/X _22855_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _22857_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_168_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _12610_/A hold868/X _12643_/B vssd1 vssd1 vccd1 vccd1 _12613_/A sky130_fd_sc_hd__and3_1
XFILLER_0_183_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21808_ _23088_/A vssd1 vssd1 vccd1 vccd1 _23087_/A sky130_fd_sc_hd__inv_2
XFILLER_0_94_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25576_ _26066_/CLK _25576_/D vssd1 vssd1 vccd1 vccd1 _25576_/Q sky130_fd_sc_hd__dfxtp_1
X_13590_ _13703_/A _13590_/B vssd1 vssd1 vccd1 vccd1 _13590_/Y sky130_fd_sc_hd__nand2_1
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22788_ _22778_/Y _22787_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22788_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_151_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ _12518_/Y _12548_/C _12533_/X _24871_/B vssd1 vssd1 vccd1 vccd1 _12542_/A
+ sky130_fd_sc_hd__a22o_1
X_24527_ _24527_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24528_/A sky130_fd_sc_hd__and2_1
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21739_ _18246_/A _21045_/B _21737_/Y _21738_/Y vssd1 vssd1 vccd1 vccd1 _21740_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15260_ _15261_/A _15262_/A vssd1 vssd1 vccd1 vccd1 _15264_/A sky130_fd_sc_hd__nor2_1
X_24458_ hold2592/X _26217_/Q _24510_/S vssd1 vssd1 vccd1 vccd1 _24458_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14211_ hold474/X _14210_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold475/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23409_ _24942_/S hold323/A _23408_/X vssd1 vssd1 vccd1 vccd1 _23409_/Y sky130_fd_sc_hd__o21ai_1
X_15191_ _15191_/A _15774_/B vssd1 vssd1 vccd1 vccd1 _15192_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_149_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24389_ _24389_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24390_/A sky130_fd_sc_hd__and2_1
XANTENNA_9 _24946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26128_ _26130_/CLK _26128_/D vssd1 vssd1 vccd1 vccd1 _26128_/Q sky130_fd_sc_hd__dfxtp_1
X_14142_ _14180_/A _14142_/B vssd1 vssd1 vccd1 vccd1 _14142_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26059_ _26060_/CLK _26059_/D vssd1 vssd1 vccd1 vccd1 _26059_/Q sky130_fd_sc_hd__dfxtp_1
X_18950_ _25901_/Q _22717_/A vssd1 vssd1 vccd1 vccd1 _18958_/A sky130_fd_sc_hd__or2_2
X_14073_ _26309_/Q _13988_/X _13981_/X _14072_/Y vssd1 vssd1 vccd1 vccd1 _14074_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17901_ _20741_/B _19303_/A vssd1 vssd1 vccd1 vccd1 _17902_/B sky130_fd_sc_hd__nand2_1
X_13024_ _26266_/Q _25635_/Q vssd1 vssd1 vccd1 vccd1 _14455_/A sky130_fd_sc_hd__xor2_2
X_18881_ _18878_/X _18879_/X _18880_/X vssd1 vssd1 vccd1 vccd1 _18882_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17832_ _17832_/A _17832_/B vssd1 vssd1 vccd1 vccd1 _17834_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_156_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17763_ _17764_/B _17764_/A vssd1 vssd1 vccd1 vccd1 _17763_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_156_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14975_ _14982_/B _14974_/Y _14963_/B vssd1 vssd1 vccd1 vccd1 _14975_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16714_ _16714_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16714_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_117_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19502_ _19501_/Y _19272_/X _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19503_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13926_ _25783_/Q vssd1 vssd1 vccd1 vccd1 _18189_/B sky130_fd_sc_hd__inv_2
XFILLER_0_187_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17694_ _17699_/A _17699_/B vssd1 vssd1 vccd1 vccd1 _17698_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19433_ _19449_/B _19523_/B vssd1 vssd1 vccd1 vccd1 _19435_/A sky130_fd_sc_hd__xnor2_1
X_16645_ _16698_/A hold920/X vssd1 vssd1 vccd1 vccd1 _16645_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13857_ _25772_/Q vssd1 vssd1 vccd1 vccd1 _18935_/B sky130_fd_sc_hd__inv_2
XFILLER_0_53_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12808_ _26225_/Q _25594_/Q vssd1 vssd1 vccd1 vccd1 _14325_/A sky130_fd_sc_hd__xor2_2
X_19364_ _19364_/A _19364_/B vssd1 vssd1 vccd1 vccd1 _19364_/Y sky130_fd_sc_hd__nand2_1
X_16576_ _16563_/A _16550_/A _16562_/B vssd1 vssd1 vccd1 vccd1 _16577_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13788_ _18713_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13788_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18315_ _18315_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18315_/Y sky130_fd_sc_hd__nand2_1
X_15527_ _15528_/A _15529_/A vssd1 vssd1 vccd1 vccd1 _15531_/A sky130_fd_sc_hd__nor2_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12739_ _16702_/A vssd1 vssd1 vccd1 vccd1 _16773_/A sky130_fd_sc_hd__clkinv_4
X_19295_ _19293_/X _19294_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19295_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18246_ _18246_/A _21021_/A vssd1 vssd1 vccd1 vccd1 _18596_/A sky130_fd_sc_hd__xor2_4
X_15458_ _15458_/A _15458_/B vssd1 vssd1 vccd1 vccd1 _15459_/B sky130_fd_sc_hd__and2_1
XFILLER_0_155_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14409_ _14409_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14409_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_5_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18177_ _19074_/A _18177_/B vssd1 vssd1 vccd1 vccd1 _18177_/X sky130_fd_sc_hd__xor2_1
X_15389_ _15389_/A vssd1 vssd1 vccd1 vccd1 _15405_/A sky130_fd_sc_hd__inv_2
XFILLER_0_163_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17128_ _20586_/B _25853_/Q _25789_/Q vssd1 vssd1 vccd1 vccd1 _17129_/B sky130_fd_sc_hd__mux2_2
Xhold504 hold504/A vssd1 vssd1 vccd1 vccd1 hold504/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold515 hold515/A vssd1 vssd1 vccd1 vccd1 hold515/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold526 hold526/A vssd1 vssd1 vccd1 vccd1 hold526/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 hold537/A vssd1 vssd1 vccd1 vccd1 hold537/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold548 hold548/A vssd1 vssd1 vccd1 vccd1 hold548/X sky130_fd_sc_hd__dlygate4sd3_1
X_17059_ _17434_/A _17512_/A vssd1 vssd1 vccd1 vccd1 _17060_/B sky130_fd_sc_hd__xnor2_1
Xhold559 hold559/A vssd1 vssd1 vccd1 vccd1 hold559/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20070_ _20070_/A _20070_/B vssd1 vssd1 vccd1 vccd1 _20978_/C sky130_fd_sc_hd__xnor2_4
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 _14857_/Y vssd1 vssd1 vccd1 vccd1 _25406_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_148_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1215 _25098_/Q vssd1 vssd1 vccd1 vccd1 _18679_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1226 _16979_/Y vssd1 vssd1 vccd1 vccd1 hold1226/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1237 _19739_/Y vssd1 vssd1 vccd1 vccd1 _25753_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 _25567_/Q vssd1 vssd1 vccd1 vccd1 _16893_/B sky130_fd_sc_hd__buf_1
XFILLER_0_100_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1259 _19943_/Y vssd1 vssd1 vccd1 vccd1 _25768_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_164_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23760_ _23760_/A vssd1 vssd1 vccd1 vccd1 _25991_/D sky130_fd_sc_hd__clkbuf_1
X_20972_ _20972_/A _20972_/B vssd1 vssd1 vccd1 vccd1 _20974_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22711_ _22711_/A _23001_/B _22711_/C vssd1 vssd1 vccd1 vccd1 _22711_/X sky130_fd_sc_hd__and3_1
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23691_ _23691_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23692_/A sky130_fd_sc_hd__and2_1
XFILLER_0_67_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25430_ _25913_/CLK _25430_/D vssd1 vssd1 vccd1 vccd1 _25430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22642_ _22642_/A _22642_/B vssd1 vssd1 vccd1 vccd1 _22642_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_177_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22573_ _22940_/B _23088_/B vssd1 vssd1 vccd1 vccd1 _22574_/B sky130_fd_sc_hd__nand2_1
X_25361_ _26190_/CLK hold295/X vssd1 vssd1 vccd1 vccd1 hold293/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24312_ _24312_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24313_/A sky130_fd_sc_hd__and2_1
XFILLER_0_145_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21524_ _21524_/A _22902_/B vssd1 vssd1 vccd1 vccd1 _21524_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_161_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25292_ _26117_/CLK hold328/X vssd1 vssd1 vccd1 vccd1 hold326/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24243_ hold2004/X _26147_/Q _24279_/S vssd1 vssd1 vccd1 vccd1 _24243_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21455_ _26324_/Q hold839/X vssd1 vssd1 vccd1 vccd1 _21455_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_105_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20406_ _20409_/A _20409_/C vssd1 vssd1 vccd1 vccd1 _20408_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24174_ _24174_/A vssd1 vssd1 vccd1 vccd1 _26124_/D sky130_fd_sc_hd__clkbuf_1
X_21386_ _21386_/A _21434_/A vssd1 vssd1 vccd1 vccd1 _21387_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_32_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23125_ _15739_/B _22893_/A _22829_/X vssd1 vssd1 vccd1 vccd1 _23125_/Y sky130_fd_sc_hd__a21oi_1
X_20337_ _21169_/C _21499_/A vssd1 vssd1 vccd1 vccd1 _20338_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_31_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23056_ _23056_/A _23056_/B vssd1 vssd1 vccd1 vccd1 _23057_/B sky130_fd_sc_hd__nand2_1
X_20268_ _20268_/A _20268_/B vssd1 vssd1 vccd1 vccd1 _20269_/A sky130_fd_sc_hd__nand2_1
X_22007_ _18226_/A _25801_/Q _22005_/Y _22006_/Y vssd1 vssd1 vccd1 vccd1 _22008_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20199_ _20199_/A _22237_/B vssd1 vssd1 vccd1 vccd1 _20200_/A sky130_fd_sc_hd__nand2_1
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2450 _25687_/Q vssd1 vssd1 vccd1 vccd1 _13329_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2461 _15463_/Y vssd1 vssd1 vccd1 vccd1 hold2461/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2472 _25461_/Q vssd1 vssd1 vccd1 vccd1 _15562_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2483 _12680_/A vssd1 vssd1 vccd1 vccd1 _12684_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2494 _26078_/Q vssd1 vssd1 vccd1 vccd1 hold2494/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1760 _21542_/Y vssd1 vssd1 vccd1 vccd1 _25826_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _14758_/Y _14759_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14760_/Y sky130_fd_sc_hd__a21oi_1
Xhold1771 _25859_/Q vssd1 vssd1 vccd1 vccd1 _22384_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23958_ _23958_/A vssd1 vssd1 vccd1 vccd1 _26054_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1782 _25863_/Q vssd1 vssd1 vccd1 vccd1 _22485_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1793 _25621_/Q vssd1 vssd1 vccd1 vccd1 _17482_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13711_ hold378/X _13710_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold379/A sky130_fd_sc_hd__a21oi_1
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22909_ _22909_/A _22909_/B vssd1 vssd1 vccd1 vccd1 _22910_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_168_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ _14703_/B _21722_/A vssd1 vssd1 vccd1 vccd1 _21721_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23889_ hold2136/X hold2080/X _23907_/S vssd1 vssd1 vccd1 vccd1 _23890_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_169_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16430_ _16430_/A _16441_/B vssd1 vssd1 vccd1 vccd1 _16430_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25628_ _25716_/CLK _25628_/D vssd1 vssd1 vccd1 vccd1 _25628_/Q sky130_fd_sc_hd__dfxtp_4
X_13642_ _13642_/A hold596/X vssd1 vssd1 vccd1 vccd1 hold597/A sky130_fd_sc_hd__nand2_1
XFILLER_0_85_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16361_ _16361_/A _16361_/B vssd1 vssd1 vccd1 vccd1 _16379_/B sky130_fd_sc_hd__and2_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25559_ _25878_/CLK _25559_/D vssd1 vssd1 vccd1 vccd1 _25559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13573_ _13642_/A hold786/X vssd1 vssd1 vccd1 vccd1 hold787/A sky130_fd_sc_hd__nand2_1
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18100_ _18100_/A vssd1 vssd1 vccd1 vccd1 _18955_/A sky130_fd_sc_hd__clkbuf_16
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _15310_/X hold2407/X _15090_/X vssd1 vssd1 vccd1 vccd1 _15312_/Y sky130_fd_sc_hd__a21oi_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _25260_/Q _25259_/Q vssd1 vssd1 vccd1 vccd1 _12525_/A sky130_fd_sc_hd__nor2_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19080_ _19080_/A _19080_/B vssd1 vssd1 vccd1 vccd1 _19081_/B sky130_fd_sc_hd__xnor2_1
X_16292_ hold863/X vssd1 vssd1 vccd1 vccd1 _16292_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18031_ _18612_/A _25725_/Q _18083_/C vssd1 vssd1 vccd1 vccd1 _18032_/C sky130_fd_sc_hd__nand3_1
X_15243_ _22628_/B _15776_/B vssd1 vssd1 vccd1 vccd1 _15244_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15174_ _22526_/B _16369_/B vssd1 vssd1 vccd1 vccd1 _16203_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14125_ _14125_/A vssd1 vssd1 vccd1 vccd1 _14236_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19982_ _19983_/B _19983_/A vssd1 vssd1 vccd1 vccd1 _19982_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18933_ _18933_/A _25836_/Q _18933_/C vssd1 vssd1 vccd1 vccd1 _20050_/B sky130_fd_sc_hd__nand3_1
X_14056_ hold513/X _14055_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold514/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ _12930_/X _13004_/X _13005_/X _13006_/X vssd1 vssd1 vccd1 vccd1 _13007_/X
+ sky130_fd_sc_hd__o211a_1
X_18864_ _25705_/Q _20791_/B vssd1 vssd1 vccd1 vccd1 _18867_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17815_ _20668_/B _22280_/A vssd1 vssd1 vccd1 vccd1 _20662_/A sky130_fd_sc_hd__nand2_2
X_18795_ _20643_/B _22515_/A vssd1 vssd1 vccd1 vccd1 _20634_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17746_ _17709_/A _17738_/A _17709_/C vssd1 vssd1 vccd1 vccd1 _17759_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_168_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14958_ _14964_/B _14959_/A vssd1 vssd1 vccd1 vccd1 _14958_/X sky130_fd_sc_hd__or2_1
XFILLER_0_159_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13909_ _26283_/Q _13801_/X _13793_/X _13908_/Y vssd1 vssd1 vccd1 vccd1 _13910_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17677_ _17706_/A _17685_/C vssd1 vssd1 vccd1 vccd1 _17721_/B sky130_fd_sc_hd__nand2_1
X_14889_ _25859_/Q _13466_/A _14888_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14890_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_187_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16628_ _16642_/B _16628_/B vssd1 vssd1 vccd1 vccd1 _16647_/A sky130_fd_sc_hd__and2_1
X_19416_ _19416_/A _20994_/B vssd1 vssd1 vccd1 vccd1 _19416_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_174_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16559_ _16557_/X _16558_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 hold905/A sky130_fd_sc_hd__a21oi_1
X_19347_ _20855_/A _19345_/Y _20860_/C vssd1 vssd1 vccd1 vccd1 _19435_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_17_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19278_ _19294_/B _19364_/B vssd1 vssd1 vccd1 vccd1 _19280_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18229_ _18535_/A _18229_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _18229_/X sky130_fd_sc_hd__and3_1
XFILLER_0_26_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21240_ _21240_/A _25874_/Q vssd1 vssd1 vccd1 vccd1 _21244_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_130_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold301 hold301/A vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 hold312/A vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold323 hold323/A vssd1 vssd1 vccd1 vccd1 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 hold334/A vssd1 vssd1 vccd1 vccd1 hold334/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21171_ _21580_/B _21630_/B vssd1 vssd1 vccd1 vccd1 _21172_/C sky130_fd_sc_hd__nand2_1
Xhold345 hold345/A vssd1 vssd1 vccd1 vccd1 hold345/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold356 hold356/A vssd1 vssd1 vccd1 vccd1 hold356/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 hold367/A vssd1 vssd1 vccd1 vccd1 hold367/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20122_ _20122_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20127_/A sky130_fd_sc_hd__nand2_2
Xhold378 hold378/A vssd1 vssd1 vccd1 vccd1 hold378/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 hold389/A vssd1 vssd1 vccd1 vccd1 hold389/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24930_ _24930_/A _25912_/Q vssd1 vssd1 vccd1 vccd1 _24930_/Y sky130_fd_sc_hd__nand2_1
X_20053_ _21693_/A vssd1 vssd1 vccd1 vccd1 _21692_/A sky130_fd_sc_hd__inv_2
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 _25027_/Q vssd1 vssd1 vccd1 vccd1 _17353_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1012 _13114_/X vssd1 vssd1 vccd1 vccd1 _25071_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24861_ _15625_/A _15640_/B _24863_/S vssd1 vssd1 vccd1 vccd1 _24861_/X sky130_fd_sc_hd__mux2_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 _25034_/Q vssd1 vssd1 vccd1 vccd1 _17424_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 _13098_/X vssd1 vssd1 vccd1 vccd1 _25068_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1045 _25026_/Q vssd1 vssd1 vccd1 vccd1 _17343_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1056 _19879_/Y vssd1 vssd1 vccd1 vccd1 _25763_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23812_ hold2036/X hold1943/X _23831_/S vssd1 vssd1 vccd1 vccd1 _23813_/A sky130_fd_sc_hd__mux2_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1067 _25014_/Q vssd1 vssd1 vccd1 vccd1 _17187_/B sky130_fd_sc_hd__dlygate4sd3_1
X_24792_ _24792_/A vssd1 vssd1 vccd1 vccd1 _26325_/D sky130_fd_sc_hd__clkbuf_1
Xhold1078 _19215_/Y vssd1 vssd1 vccd1 vccd1 _25716_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1089 _25744_/Q vssd1 vssd1 vccd1 vccd1 _19610_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23743_ _23743_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23744_/A sky130_fd_sc_hd__and2_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20955_ _26302_/Q _20731_/X hold437/X vssd1 vssd1 vccd1 vccd1 _20959_/B sky130_fd_sc_hd__a21oi_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23674_ hold2243/X hold2071/X _23677_/S vssd1 vssd1 vccd1 vccd1 _23675_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_49_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ _20886_/A _21874_/B _20886_/C vssd1 vssd1 vccd1 vccd1 _20889_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25413_ _26004_/CLK _25413_/D vssd1 vssd1 vccd1 vccd1 _25413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22625_ _22625_/A _22625_/B vssd1 vssd1 vccd1 vccd1 _22626_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25344_ _26298_/CLK hold100/X vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22556_ _22555_/A _22454_/X _22555_/B vssd1 vssd1 vccd1 vccd1 _22557_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21507_ _21507_/A _21507_/B vssd1 vssd1 vccd1 vccd1 _21508_/A sky130_fd_sc_hd__nand2_1
X_25275_ _26231_/CLK hold337/X vssd1 vssd1 vccd1 vccd1 hold335/A sky130_fd_sc_hd__dfxtp_1
X_22487_ _22487_/A _25892_/Q vssd1 vssd1 vccd1 vccd1 _22487_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24226_ _24226_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24227_/A sky130_fd_sc_hd__and2_1
XFILLER_0_47_1140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21438_ _26323_/Q _21228_/X hold647/X vssd1 vssd1 vccd1 vccd1 _21441_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24157_ hold2307/X _26119_/Q _24203_/S vssd1 vssd1 vccd1 vccd1 _24157_/X sky130_fd_sc_hd__mux2_1
X_21369_ _21369_/A _21417_/A vssd1 vssd1 vccd1 vccd1 _21371_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_102_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23108_ _23188_/A _23108_/B vssd1 vssd1 vccd1 vccd1 _23108_/X sky130_fd_sc_hd__or2_1
X_24088_ _24088_/A vssd1 vssd1 vccd1 vccd1 _26096_/D sky130_fd_sc_hd__clkbuf_1
Xhold890 hold890/A vssd1 vssd1 vccd1 vccd1 hold890/X sky130_fd_sc_hd__dlygate4sd3_1
X_15930_ _21967_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _15932_/A sky130_fd_sc_hd__nand2_1
X_23039_ _23039_/A _23039_/B vssd1 vssd1 vccd1 vccd1 _23041_/A sky130_fd_sc_hd__nand2_1
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15861_ _15956_/A hold692/X vssd1 vssd1 vccd1 vccd1 hold693/A sky130_fd_sc_hd__nand2_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2280 _26135_/Q vssd1 vssd1 vccd1 vccd1 hold2280/X sky130_fd_sc_hd__dlygate4sd3_1
X_17600_ _17600_/A _17651_/A vssd1 vssd1 vccd1 vccd1 _17601_/B sky130_fd_sc_hd__xnor2_1
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812_ _14812_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14812_/Y sky130_fd_sc_hd__nand2_1
Xhold2291 _25982_/Q vssd1 vssd1 vccd1 vccd1 _14705_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18580_ _18641_/A _19416_/A vssd1 vssd1 vccd1 vccd1 _18580_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_99_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15792_ _15792_/A _15810_/B vssd1 vssd1 vccd1 vccd1 _15793_/B sky130_fd_sc_hd__nand2_2
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1590 _25883_/Q vssd1 vssd1 vccd1 vccd1 _22903_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17531_ _17531_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17531_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14743_ _15839_/A _14743_/B vssd1 vssd1 vccd1 vccd1 _21900_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17462_ _17512_/A _17629_/B vssd1 vssd1 vccd1 vccd1 _17463_/B sky130_fd_sc_hd__xnor2_1
X_14674_ _14672_/Y hold348/X _14646_/X vssd1 vssd1 vccd1 vccd1 hold349/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16413_ _16413_/A _16413_/B vssd1 vssd1 vccd1 vccd1 _16414_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_156_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19201_ _19198_/Y _19200_/Y _19086_/X vssd1 vssd1 vccd1 vccd1 _19201_/Y sky130_fd_sc_hd__a21oi_1
X_13625_ _25735_/Q vssd1 vssd1 vccd1 vccd1 _18172_/B sky130_fd_sc_hd__inv_2
X_17393_ _17393_/A _17393_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17393_/X sky130_fd_sc_hd__and3_1
XFILLER_0_184_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19132_ _19129_/Y _19130_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19136_/A
+ sky130_fd_sc_hd__a211o_1
X_16344_ _16341_/Y _16342_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 hold907/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13556_ _17989_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13556_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_55_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12507_ _23923_/A _24970_/Q _12560_/A _12507_/D vssd1 vssd1 vccd1 vccd1 _24050_/B
+ sky130_fd_sc_hd__or4_4
X_19063_ _19063_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _19063_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16275_ _16264_/B _16269_/A _16252_/B _16269_/X _16263_/A vssd1 vssd1 vccd1 vccd1
+ _16275_/X sky130_fd_sc_hd__o221a_1
X_13487_ hold815/A vssd1 vssd1 vccd1 vccd1 _17927_/B sky130_fd_sc_hd__inv_2
XFILLER_0_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18014_ _25651_/Q vssd1 vssd1 vccd1 vccd1 _21924_/A sky130_fd_sc_hd__inv_2
X_15226_ _22603_/B _15776_/B vssd1 vssd1 vccd1 vccd1 _16248_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_124_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15157_ _15158_/A _15159_/A vssd1 vssd1 vccd1 vccd1 _15161_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_121_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14108_ _18450_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14108_/Y sky130_fd_sc_hd__nor2_1
X_15088_ _15106_/A _15089_/A vssd1 vssd1 vccd1 vccd1 _15088_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19965_ _19963_/Y _19964_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _19965_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14039_ _14118_/A hold371/X vssd1 vssd1 vccd1 vccd1 hold372/A sky130_fd_sc_hd__nand2_1
X_18916_ _20006_/B _22667_/A vssd1 vssd1 vccd1 vccd1 _19999_/A sky130_fd_sc_hd__nand2_2
X_19896_ _19896_/A _19980_/B _19896_/C vssd1 vssd1 vccd1 vccd1 _19896_/X sky130_fd_sc_hd__and3_1
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18847_ _18847_/A _18847_/B vssd1 vssd1 vccd1 vccd1 _22589_/A sky130_fd_sc_hd__or2_1
XFILLER_0_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18778_ _18778_/A _18778_/B vssd1 vssd1 vccd1 vccd1 _18778_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_136_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17729_ _17766_/B _17729_/B vssd1 vssd1 vccd1 vccd1 _17734_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20740_ _20740_/A _21729_/B vssd1 vssd1 vccd1 vccd1 _20741_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_147_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20671_ _21371_/B vssd1 vssd1 vccd1 vccd1 _21368_/C sky130_fd_sc_hd__inv_2
XFILLER_0_169_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22410_ _22410_/A _22410_/B vssd1 vssd1 vccd1 vccd1 _22410_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_163_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23390_ _24942_/S hold236/A _23389_/X vssd1 vssd1 vccd1 vccd1 _23390_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22341_ _22561_/A _22341_/B vssd1 vssd1 vccd1 vccd1 _22341_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22272_ _22272_/A _22272_/B vssd1 vssd1 vccd1 vccd1 _22273_/B sky130_fd_sc_hd__nand2_1
X_25060_ _26146_/CLK _25060_/D vssd1 vssd1 vccd1 vccd1 _25060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24011_ hold2425/X _26072_/Q _24047_/S vssd1 vssd1 vccd1 vccd1 _24011_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21223_ _21662_/B _21613_/B vssd1 vssd1 vccd1 vccd1 _21225_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_131_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold120 hold120/A vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 hold131/A vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 hold142/A vssd1 vssd1 vccd1 vccd1 hold142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 hold153/A vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 hold164/A vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlygate4sd3_1
X_21154_ _21235_/A _21154_/B vssd1 vssd1 vccd1 vccd1 _21154_/Y sky130_fd_sc_hd__nand2_1
Xhold175 hold175/A vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold186 hold186/A vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 hold197/A vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
X_20105_ _20105_/A _20105_/B vssd1 vssd1 vccd1 vccd1 _20107_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25962_ _26042_/CLK _25962_/D vssd1 vssd1 vccd1 vccd1 _25962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21085_ _21532_/B _21580_/B vssd1 vssd1 vccd1 vccd1 _21086_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24913_ hold970/A _25523_/Q _24922_/S vssd1 vssd1 vccd1 vccd1 _24914_/B sky130_fd_sc_hd__mux2_1
X_20036_ _26277_/Q hold722/X vssd1 vssd1 vccd1 vccd1 _20036_/Y sky130_fd_sc_hd__nand2_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25893_ _25893_/CLK _25893_/D vssd1 vssd1 vccd1 vccd1 _25893_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24844_ _24840_/X _24843_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _24844_/X sky130_fd_sc_hd__mux2_1
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24775_ hold2636/X _26320_/Q _24817_/S vssd1 vssd1 vccd1 vccd1 _24775_/X sky130_fd_sc_hd__mux2_1
X_21987_ _21987_/A _21987_/B vssd1 vssd1 vccd1 vccd1 _22729_/A sky130_fd_sc_hd__nand2_2
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23726_ _23726_/A vssd1 vssd1 vccd1 vccd1 _25980_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ _20938_/A _25863_/Q vssd1 vssd1 vccd1 vccd1 _20944_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_139_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23657_ _23657_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23658_/A sky130_fd_sc_hd__and2_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20869_ _21676_/A _21448_/C vssd1 vssd1 vccd1 vccd1 _20871_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_187_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13410_ _26203_/Q _13239_/X _13409_/X vssd1 vssd1 vccd1 vccd1 _13410_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22608_ _22608_/A _23001_/B _22608_/C vssd1 vssd1 vccd1 vccd1 _22608_/X sky130_fd_sc_hd__and3_1
XFILLER_0_148_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14390_ _14388_/Y hold252/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold253/A sky130_fd_sc_hd__a21oi_1
X_23588_ hold985/X _25922_/Q hold855/X _25920_/Q vssd1 vssd1 vccd1 vccd1 _23590_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_0_9_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25327_ _26151_/CLK hold250/X vssd1 vssd1 vccd1 vccd1 hold248/A sky130_fd_sc_hd__dfxtp_1
X_13341_ _13341_/A vssd1 vssd1 vccd1 vccd1 _19644_/A sky130_fd_sc_hd__clkbuf_8
X_22539_ _25830_/Q _22539_/B vssd1 vssd1 vccd1 vccd1 _22539_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_51_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16060_ _16055_/Y _15846_/B _16059_/X vssd1 vssd1 vccd1 vccd1 _16160_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_161_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25258_ _26046_/CLK _25258_/D vssd1 vssd1 vccd1 vccd1 _25258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13272_ _26309_/Q _19488_/A vssd1 vssd1 vccd1 vccd1 _14593_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_161_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15011_ _15009_/X hold2197/X _14928_/X vssd1 vssd1 vccd1 vccd1 _15011_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24209_ _24209_/A vssd1 vssd1 vccd1 vccd1 _26135_/D sky130_fd_sc_hd__clkbuf_1
X_25189_ _26273_/CLK hold814/X vssd1 vssd1 vccd1 vccd1 hold812/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19750_ _19748_/X _19749_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19750_/Y sky130_fd_sc_hd__a21oi_1
X_16962_ _16962_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16962_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18701_ _18701_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18701_/Y sky130_fd_sc_hd__nand2_1
X_15913_ _15956_/A hold858/X vssd1 vssd1 vccd1 vccd1 _15913_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_21_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16893_ _16977_/A _16893_/B vssd1 vssd1 vccd1 vccd1 _16893_/Y sky130_fd_sc_hd__nand2_1
X_19681_ _19723_/A _19681_/B vssd1 vssd1 vccd1 vccd1 _19681_/Y sky130_fd_sc_hd__nand2_1
X_15844_ _15844_/A _15844_/B vssd1 vssd1 vccd1 vccd1 _15845_/B sky130_fd_sc_hd__nand2_1
X_18632_ _18955_/A _18632_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18633_/C sky130_fd_sc_hd__nand3_1
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15775_ _23159_/B _15775_/B vssd1 vssd1 vccd1 vccd1 _23156_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18563_ _22237_/B _25626_/Q vssd1 vssd1 vccd1 vccd1 _18565_/A sky130_fd_sc_hd__nand2_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _26259_/Q _25628_/Q vssd1 vssd1 vccd1 vccd1 _14434_/A sky130_fd_sc_hd__xor2_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14726_ _21830_/B _15778_/B vssd1 vssd1 vccd1 vccd1 _14727_/A sky130_fd_sc_hd__nand2_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17514_ _17624_/A _17514_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17514_/X sky130_fd_sc_hd__and3_1
XFILLER_0_185_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18494_ _18494_/A _18494_/B vssd1 vssd1 vccd1 vccd1 _18494_/X sky130_fd_sc_hd__xor2_1
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17445_ _17467_/A _17445_/B vssd1 vssd1 vccd1 vccd1 _17445_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14657_ _14657_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _14657_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_28_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13608_ _26235_/Q _13426_/X _13605_/X _13607_/Y vssd1 vssd1 vccd1 vccd1 _13609_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_184_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17376_ _17467_/A _17376_/B vssd1 vssd1 vccd1 vccd1 _17376_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_166_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14588_ _14588_/A vssd1 vssd1 vccd1 vccd1 _14644_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_171_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16327_ _16325_/X _16326_/Y _16076_/X vssd1 vssd1 vccd1 vccd1 hold874/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19115_ _25648_/Q _19115_/B _19115_/C vssd1 vssd1 vccd1 vccd1 _20113_/A sky130_fd_sc_hd__or3_1
X_13539_ _26224_/Q _13426_/X _13468_/X _13538_/Y vssd1 vssd1 vccd1 vccd1 _13540_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19046_ _19046_/A _19046_/B vssd1 vssd1 vccd1 vccd1 _19046_/X sky130_fd_sc_hd__xor2_1
X_16258_ _16256_/X _16257_/Y _16076_/X vssd1 vssd1 vccd1 vccd1 hold890/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15209_ _22577_/B _16369_/B vssd1 vssd1 vccd1 vccd1 _15210_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16189_ _16189_/A _16189_/B vssd1 vssd1 vccd1 vccd1 _16215_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_3_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19948_ _19948_/A _19959_/A vssd1 vssd1 vccd1 vccd1 _19950_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19879_ _19877_/Y _19878_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19879_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21910_ _21910_/A _21910_/B vssd1 vssd1 vccd1 vccd1 _23136_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_156_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22890_ _23042_/A _22890_/B vssd1 vssd1 vccd1 vccd1 _22891_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21841_ _21841_/A _21841_/B vssd1 vssd1 vccd1 vccd1 _23104_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_37_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24560_ _24560_/A vssd1 vssd1 vccd1 vccd1 _24649_/B sky130_fd_sc_hd__buf_6
XFILLER_0_37_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21772_ _21772_/A _25867_/Q vssd1 vssd1 vccd1 vccd1 _21772_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_148_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23511_ hold98/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23511_/X sky130_fd_sc_hd__or2b_1
X_20723_ _21661_/B vssd1 vssd1 vccd1 vccd1 _21660_/B sky130_fd_sc_hd__inv_2
X_24491_ _24491_/A vssd1 vssd1 vccd1 vccd1 _26227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26230_ _26232_/CLK _26230_/D vssd1 vssd1 vccd1 vccd1 _26230_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23442_ hold308/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23442_/X sky130_fd_sc_hd__or2b_1
X_20654_ _26293_/Q _20078_/X hold638/X vssd1 vssd1 vccd1 vccd1 _20657_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26161_ _26289_/CLK _26161_/D vssd1 vssd1 vccd1 vccd1 _26161_/Q sky130_fd_sc_hd__dfxtp_1
X_23373_ _23373_/A _23377_/B _23373_/C vssd1 vssd1 vccd1 vccd1 _23373_/X sky130_fd_sc_hd__and3_1
X_20585_ _20585_/A _22219_/B vssd1 vssd1 vccd1 vccd1 _20586_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_144_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25112_ _26330_/CLK _25112_/D vssd1 vssd1 vccd1 vccd1 _25112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22324_ _22322_/X _15839_/B _22323_/Y _14873_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _22325_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_143_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26092_ _26221_/CLK _26092_/D vssd1 vssd1 vccd1 vccd1 _26092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25043_ _26130_/CLK _25043_/D vssd1 vssd1 vccd1 vccd1 _25043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22255_ _23007_/B vssd1 vssd1 vccd1 vccd1 _23154_/A sky130_fd_sc_hd__inv_2
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21206_ _21206_/A _21206_/B vssd1 vssd1 vccd1 vccd1 _21207_/A sky130_fd_sc_hd__nand2_1
X_22186_ _22840_/B vssd1 vssd1 vccd1 vccd1 _22841_/A sky130_fd_sc_hd__inv_2
XFILLER_0_100_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21137_ _21137_/A _21137_/B vssd1 vssd1 vccd1 vccd1 _21610_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_100_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25945_ _26009_/CLK _25945_/D vssd1 vssd1 vccd1 vccd1 _25945_/Q sky130_fd_sc_hd__dfxtp_1
X_21068_ _21067_/Y _20192_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21068_/X
+ sky130_fd_sc_hd__a211o_1
X_12910_ _12891_/X _14385_/A _12909_/X _25613_/Q vssd1 vssd1 vccd1 vccd1 _12910_/X
+ sky130_fd_sc_hd__a22o_1
X_20019_ _20019_/A _20019_/B vssd1 vssd1 vccd1 vccd1 _21370_/A sky130_fd_sc_hd__nand2_2
X_25876_ _25876_/CLK _25876_/D vssd1 vssd1 vccd1 vccd1 _25876_/Q sky130_fd_sc_hd__dfxtp_2
X_13890_ _17931_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13890_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_159_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24827_ _24827_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24828_/A sky130_fd_sc_hd__and2_1
X_12841_ _26231_/Q _25600_/Q vssd1 vssd1 vccd1 vccd1 _14343_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_69_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _15560_/A _15577_/B vssd1 vssd1 vccd1 vccd1 _15560_/Y sky130_fd_sc_hd__nand2_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _12746_/X _12770_/X _14910_/B _12771_/X vssd1 vssd1 vccd1 vccd1 hold961/A
+ sky130_fd_sc_hd__o211a_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24758_ _24758_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24759_/A sky130_fd_sc_hd__and2_1
XFILLER_0_189_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14509_/Y hold90/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__a21oi_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23709_ _23709_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23710_/A sky130_fd_sc_hd__and2_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _22893_/B _16369_/B vssd1 vssd1 vccd1 vccd1 _15492_/A sky130_fd_sc_hd__nand2_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24689_ hold2596/X _26292_/Q _24740_/S vssd1 vssd1 vccd1 vccd1 _24689_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_166_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17272_/A _17230_/B vssd1 vssd1 vccd1 vccd1 _17230_/Y sky130_fd_sc_hd__nand2_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _14440_/Y hold114/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold115/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17161_ _17393_/A _17161_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17161_/X sky130_fd_sc_hd__and3_1
XFILLER_0_80_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14373_ _14373_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14373_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_52_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16112_ _16113_/B _16113_/A vssd1 vssd1 vccd1 vccd1 _16125_/B sky130_fd_sc_hd__or2_1
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13324_ _13220_/X _14617_/A _13242_/X _19602_/A vssd1 vssd1 vccd1 vccd1 _13324_/X
+ sky130_fd_sc_hd__a22o_1
X_17092_ _17645_/A _17092_/B vssd1 vssd1 vccd1 vccd1 _17092_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_134_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16043_ _16041_/X _16042_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _16043_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_150_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13255_ _13220_/X _14581_/A _13242_/X _19444_/A vssd1 vssd1 vccd1 vccd1 _13255_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13186_ _18393_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13186_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19802_ _19802_/A _20597_/B vssd1 vssd1 vccd1 vccd1 _19802_/Y sky130_fd_sc_hd__nor2_1
X_17994_ _21801_/B _25603_/Q vssd1 vssd1 vccd1 vccd1 _17996_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19733_ _19734_/B _19734_/A vssd1 vssd1 vccd1 vccd1 _19733_/X sky130_fd_sc_hd__or2_1
X_16945_ _16946_/B _16946_/A vssd1 vssd1 vccd1 vccd1 _16945_/X sky130_fd_sc_hd__or2_1
X_19664_ _19664_/A _19664_/B vssd1 vssd1 vccd1 vccd1 _19664_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_95_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16876_ _16876_/A _16876_/B vssd1 vssd1 vccd1 vccd1 _16876_/Y sky130_fd_sc_hd__nand2_1
X_18615_ _18615_/A _20272_/A vssd1 vssd1 vccd1 vccd1 _18960_/A sky130_fd_sc_hd__xor2_4
X_15827_ _15827_/A _15827_/B vssd1 vssd1 vccd1 vccd1 _15836_/A sky130_fd_sc_hd__nand2_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19595_ _19587_/X _19594_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19595_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_172_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15758_ _15795_/A _16651_/B vssd1 vssd1 vccd1 vccd1 _16960_/A sky130_fd_sc_hd__or2_2
X_18546_ _18792_/A _18550_/B vssd1 vssd1 vccd1 vccd1 _18548_/A sky130_fd_sc_hd__nand2_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14709_ _25839_/Q _12527_/A _14916_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14709_/X
+ sky130_fd_sc_hd__a22o_1
X_15689_ _15689_/A vssd1 vssd1 vccd1 vccd1 _15691_/A sky130_fd_sc_hd__inv_2
XFILLER_0_158_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18477_ _18477_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18477_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17428_ _17568_/A vssd1 vssd1 vccd1 vccd1 _17428_/X sky130_fd_sc_hd__buf_6
XFILLER_0_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17359_ _21157_/B _25871_/Q _25807_/Q vssd1 vssd1 vccd1 vccd1 _17360_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20370_ _20370_/A _20370_/B _20370_/C vssd1 vssd1 vccd1 vccd1 _20371_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19029_ _19186_/A _19816_/A vssd1 vssd1 vccd1 vccd1 _19029_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_140_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22040_ _25811_/Q _22040_/B vssd1 vssd1 vccd1 vccd1 _22040_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_100_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23991_ _23991_/A vssd1 vssd1 vccd1 vccd1 _26065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25730_ _26236_/CLK _25730_/D vssd1 vssd1 vccd1 vccd1 _25730_/Q sky130_fd_sc_hd__dfxtp_1
X_22942_ _22942_/A _22942_/B vssd1 vssd1 vccd1 vccd1 _22943_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25661_ _26292_/CLK _25661_/D vssd1 vssd1 vccd1 vccd1 _25661_/Q sky130_fd_sc_hd__dfxtp_1
X_22873_ _22871_/X _22872_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _22873_/Y sky130_fd_sc_hd__a21oi_1
X_24612_ hold2700/X hold2586/X _24664_/S vssd1 vssd1 vccd1 vccd1 _24613_/A sky130_fd_sc_hd__mux2_1
X_21824_ _21825_/A _21825_/B _22926_/A vssd1 vssd1 vccd1 vccd1 _21824_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_149_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25592_ _26096_/CLK _25592_/D vssd1 vssd1 vccd1 vccd1 _25592_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_149_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24543_ _24543_/A vssd1 vssd1 vccd1 vccd1 _26244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21755_ _21753_/X _21754_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _21755_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20706_ _20708_/B _20708_/C vssd1 vssd1 vccd1 vccd1 _20707_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24474_ hold2565/X _26222_/Q _24510_/S vssd1 vssd1 vccd1 vccd1 _24474_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21686_ _21686_/A _22902_/B vssd1 vssd1 vccd1 vccd1 _21686_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26213_ _26296_/CLK _26213_/D vssd1 vssd1 vccd1 vccd1 _26213_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23425_ hold83/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23425_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_74_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20637_ _20637_/A _25893_/Q vssd1 vssd1 vccd1 vccd1 _20643_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_110_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26144_ _26263_/CLK _26144_/D vssd1 vssd1 vccd1 vccd1 _26144_/Q sky130_fd_sc_hd__dfxtp_1
X_23356_ _23356_/A _23356_/B vssd1 vssd1 vccd1 vccd1 _23357_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20568_ _21322_/B _21596_/A vssd1 vssd1 vccd1 vccd1 _20571_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_132_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22307_ _22307_/A _25856_/Q vssd1 vssd1 vccd1 vccd1 _22307_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26075_ _26079_/CLK _26075_/D vssd1 vssd1 vccd1 vccd1 _26075_/Q sky130_fd_sc_hd__dfxtp_1
X_23287_ _23287_/A _23377_/B _23287_/C vssd1 vssd1 vccd1 vccd1 _23288_/A sky130_fd_sc_hd__and3_1
XFILLER_0_104_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20499_ _26289_/Q hold742/X vssd1 vssd1 vccd1 vccd1 _20499_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_131_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25026_ _25604_/CLK _25026_/D vssd1 vssd1 vccd1 vccd1 _25026_/Q sky130_fd_sc_hd__dfxtp_1
X_13040_ _12891_/X _14464_/A _12909_/X _25638_/Q vssd1 vssd1 vccd1 vccd1 _13040_/X
+ sky130_fd_sc_hd__a22o_1
X_22238_ _18574_/A _25818_/Q _22236_/Y _22237_/Y vssd1 vssd1 vccd1 vccd1 _22239_/B
+ sky130_fd_sc_hd__a31o_1
X_22169_ _22167_/X _22168_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _22169_/Y sky130_fd_sc_hd__a21oi_2
X_14991_ _14986_/A _14981_/A _14981_/B vssd1 vssd1 vccd1 vccd1 _14993_/A sky130_fd_sc_hd__a21bo_1
X_16730_ _16728_/Y _16729_/Y _16594_/X vssd1 vssd1 vccd1 vccd1 _16730_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13942_ hold486/X _13941_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold487/A sky130_fd_sc_hd__a21oi_1
X_25928_ _25939_/CLK _25928_/D vssd1 vssd1 vccd1 vccd1 _25928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16661_ _16658_/B _16658_/A _16680_/B _16660_/Y vssd1 vssd1 vccd1 vccd1 _16661_/X
+ sky130_fd_sc_hd__a31o_1
X_25859_ _25859_/CLK _25859_/D vssd1 vssd1 vccd1 vccd1 _25859_/Q sky130_fd_sc_hd__dfxtp_4
X_13873_ hold723/X _13872_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold724/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15612_ _15612_/A _15612_/B vssd1 vssd1 vccd1 vccd1 _15612_/Y sky130_fd_sc_hd__nand2_1
X_18400_ _21238_/B _19546_/A vssd1 vssd1 vccd1 vccd1 _18401_/B sky130_fd_sc_hd__nand2_1
X_12824_ _26228_/Q _25597_/Q vssd1 vssd1 vccd1 vccd1 _14334_/A sky130_fd_sc_hd__xor2_2
X_16592_ _16592_/A _16697_/B vssd1 vssd1 vccd1 vccd1 _16592_/Y sky130_fd_sc_hd__nand2_1
X_19380_ _19372_/X _19379_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19380_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15543_ _16498_/A _15543_/B vssd1 vssd1 vccd1 vccd1 _16876_/A sky130_fd_sc_hd__nand2_1
X_18331_ _18534_/A _18678_/A vssd1 vssd1 vccd1 vccd1 _18332_/B sky130_fd_sc_hd__xnor2_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ _14064_/A vssd1 vssd1 vccd1 vccd1 _14264_/A sky130_fd_sc_hd__clkbuf_16
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18262_ _18445_/A _25739_/Q vssd1 vssd1 vccd1 vccd1 _18264_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_154_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15474_ _22882_/B _15474_/B vssd1 vssd1 vccd1 vccd1 _22879_/B sky130_fd_sc_hd__xor2_1
X_12686_ _12686_/A _12686_/B vssd1 vssd1 vccd1 vccd1 _12700_/B sky130_fd_sc_hd__nand2_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17213_ _17463_/A _17213_/B vssd1 vssd1 vccd1 vccd1 _17213_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_53_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14425_ _14425_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14425_/Y sky130_fd_sc_hd__nand2_1
X_18193_ _19402_/A vssd1 vssd1 vccd1 vccd1 _21972_/B sky130_fd_sc_hd__inv_2
XFILLER_0_182_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17144_ _20439_/B _25888_/Q _25824_/Q vssd1 vssd1 vccd1 vccd1 _17145_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14356_ _14404_/A hold254/X vssd1 vssd1 vccd1 vccd1 hold255/A sky130_fd_sc_hd__nand2_1
XFILLER_0_181_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13307_ _18779_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13307_/X sky130_fd_sc_hd__or2_1
Xhold708 hold708/A vssd1 vssd1 vccd1 vccd1 hold708/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold719 hold719/A vssd1 vssd1 vccd1 vccd1 hold719/X sky130_fd_sc_hd__dlygate4sd3_1
X_17075_ _17441_/A _17519_/A vssd1 vssd1 vccd1 vccd1 _17076_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14287_ _14287_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14287_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16026_ _16026_/A _16027_/B vssd1 vssd1 vccd1 vccd1 _16053_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_110_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13238_ _13207_/X _13236_/X _13192_/X _13237_/X vssd1 vssd1 vccd1 vccd1 _13238_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13169_ _13109_/X _13167_/X _13096_/X _13168_/X vssd1 vssd1 vccd1 vccd1 _13169_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2109 _25958_/Q vssd1 vssd1 vccd1 vccd1 hold2109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1408 _14814_/Y vssd1 vssd1 vccd1 vccd1 _25401_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17977_ _20178_/A _17977_/B vssd1 vssd1 vccd1 vccd1 _19159_/A sky130_fd_sc_hd__nand2_2
Xhold1419 _25109_/Q vssd1 vssd1 vccd1 vccd1 _18900_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19716_ _20361_/A _22348_/B _25630_/Q vssd1 vssd1 vccd1 vccd1 _20366_/C sky130_fd_sc_hd__nand3_1
X_16928_ _16935_/A _16933_/B vssd1 vssd1 vccd1 vccd1 _16930_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19647_ _19664_/B _19734_/B vssd1 vssd1 vccd1 vccd1 _19649_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_189_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16859_ _16857_/Y _16858_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16859_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19578_ _19579_/B _19579_/A vssd1 vssd1 vccd1 vccd1 _19578_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18529_ _18529_/A _18529_/B _18529_/C vssd1 vssd1 vccd1 vccd1 _18530_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_48_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21540_ _21540_/A _22902_/B vssd1 vssd1 vccd1 vccd1 _21540_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_118_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21471_ _26325_/Q hold440/X vssd1 vssd1 vccd1 vccd1 _21471_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23210_ _23210_/A vssd1 vssd1 vccd1 vccd1 _25905_/D sky130_fd_sc_hd__inv_2
XFILLER_0_145_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20422_ _20421_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20422_/X
+ sky130_fd_sc_hd__a211o_1
X_24190_ hold2189/X hold899/X _24203_/S vssd1 vssd1 vccd1 vccd1 _24192_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_71_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23141_ _15756_/B _22893_/A _22829_/X vssd1 vssd1 vccd1 vccd1 _23141_/Y sky130_fd_sc_hd__a21oi_1
X_20353_ _25847_/Q vssd1 vssd1 vccd1 vccd1 _20354_/B sky130_fd_sc_hd__inv_2
XFILLER_0_140_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23072_ _23072_/A _23072_/B vssd1 vssd1 vccd1 vccd1 _23073_/B sky130_fd_sc_hd__nand2_1
X_20284_ _20284_/A _21992_/A vssd1 vssd1 vccd1 vccd1 _20285_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_113_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22023_ _22742_/B vssd1 vssd1 vccd1 vccd1 _22743_/A sky130_fd_sc_hd__inv_2
XFILLER_0_87_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2610 _26304_/Q vssd1 vssd1 vccd1 vccd1 hold2610/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2621 _24655_/X vssd1 vssd1 vccd1 vccd1 _24656_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2632 _26276_/Q vssd1 vssd1 vccd1 vccd1 hold2632/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2643 _24550_/X vssd1 vssd1 vccd1 vccd1 _24551_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2654 _26215_/Q vssd1 vssd1 vccd1 vccd1 hold2654/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1920 _26167_/Q vssd1 vssd1 vccd1 vccd1 hold1920/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2665 _24569_/X vssd1 vssd1 vccd1 vccd1 _24570_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1931 _24203_/X vssd1 vssd1 vccd1 vccd1 _24204_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2676 _26322_/Q vssd1 vssd1 vccd1 vccd1 hold2676/X sky130_fd_sc_hd__dlygate4sd3_1
X_23974_ hold2510/X _26060_/Q _24001_/S vssd1 vssd1 vccd1 vccd1 _23974_/X sky130_fd_sc_hd__mux2_1
Xhold1942 _14281_/Y vssd1 vssd1 vccd1 vccd1 _25260_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2687 _26237_/Q vssd1 vssd1 vccd1 vccd1 hold2687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2698 _25912_/Q vssd1 vssd1 vccd1 vccd1 _23242_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1953 _15024_/Y vssd1 vssd1 vccd1 vccd1 hold1953/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1964 _23904_/X vssd1 vssd1 vccd1 vccd1 _23905_/A sky130_fd_sc_hd__dlygate4sd3_1
X_25713_ _25716_/CLK hold817/X vssd1 vssd1 vccd1 vccd1 hold815/A sky130_fd_sc_hd__dfxtp_1
Xhold1975 _23687_/X vssd1 vssd1 vccd1 vccd1 _23688_/A sky130_fd_sc_hd__dlygate4sd3_1
X_22925_ _22925_/A _22925_/B vssd1 vssd1 vccd1 vccd1 _22926_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1986 _24276_/X vssd1 vssd1 vccd1 vccd1 _24277_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1997 _26212_/Q vssd1 vssd1 vccd1 vccd1 hold1997/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25644_ _26148_/CLK _25644_/D vssd1 vssd1 vccd1 vccd1 _25644_/Q sky130_fd_sc_hd__dfxtp_2
X_22856_ _23245_/A vssd1 vssd1 vccd1 vccd1 _22856_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21807_ _21807_/A _21807_/B vssd1 vssd1 vccd1 vccd1 _23088_/A sky130_fd_sc_hd__nand2_4
X_25575_ _26080_/CLK _25575_/D vssd1 vssd1 vccd1 vccd1 _25575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22787_ _22787_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _22787_/Y sky130_fd_sc_hd__nand2_1
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12540_ _23278_/B vssd1 vssd1 vccd1 vccd1 _24871_/B sky130_fd_sc_hd__inv_2
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24526_ hold2660/X hold2557/X _24587_/S vssd1 vssd1 vccd1 vccd1 _24527_/A sky130_fd_sc_hd__mux2_1
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21738_ _25802_/Q _21738_/B vssd1 vssd1 vccd1 vccd1 _21738_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_93_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24457_ _24457_/A vssd1 vssd1 vccd1 vccd1 _26216_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21669_ _21669_/A _21669_/B vssd1 vssd1 vccd1 vccd1 _21670_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14210_ _14264_/A _14210_/B vssd1 vssd1 vccd1 vccd1 _14210_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23408_ hold116/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23408_/X sky130_fd_sc_hd__or2b_1
X_15190_ _26009_/Q _25945_/Q _15773_/S vssd1 vssd1 vccd1 vccd1 _15191_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24388_ hold1860/X _26194_/Q _24433_/S vssd1 vssd1 vccd1 vccd1 _24388_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_123_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26127_ _26130_/CLK _26127_/D vssd1 vssd1 vccd1 vccd1 _26127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14141_ _26320_/Q _13988_/X _13981_/X _14140_/Y vssd1 vssd1 vccd1 vccd1 _14142_/B
+ sky130_fd_sc_hd__a22o_1
X_23339_ _23339_/A _23377_/B _23339_/C vssd1 vssd1 vccd1 vccd1 _23339_/X sky130_fd_sc_hd__and3_1
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26058_ _26060_/CLK _26058_/D vssd1 vssd1 vccd1 vccd1 _26058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14072_ _18328_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14072_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17900_ _21729_/B _25601_/Q vssd1 vssd1 vccd1 vccd1 _17902_/A sky130_fd_sc_hd__nand2_1
X_25009_ _26096_/CLK _25009_/D vssd1 vssd1 vccd1 vccd1 _25009_/Q sky130_fd_sc_hd__dfxtp_1
X_13023_ _13018_/X _13021_/X _13005_/X _13022_/X vssd1 vssd1 vccd1 vccd1 _13023_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18880_ _19026_/A _18880_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18880_/X sky130_fd_sc_hd__and3_1
X_17831_ _17831_/A _17831_/B vssd1 vssd1 vccd1 vccd1 _17832_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17762_ _17771_/A _17771_/C vssd1 vssd1 vccd1 vccd1 _17770_/A sky130_fd_sc_hd__nand2_1
X_14974_ _15033_/A vssd1 vssd1 vccd1 vccd1 _14974_/Y sky130_fd_sc_hd__inv_2
X_19501_ _26240_/Q hold835/X vssd1 vssd1 vccd1 vccd1 _19501_/Y sky130_fd_sc_hd__nand2_1
X_16713_ _16710_/X _16711_/X _16712_/Y _25862_/Q _14170_/X vssd1 vssd1 vccd1 vccd1
+ _16714_/A sky130_fd_sc_hd__a32o_1
X_13925_ _14000_/A hold536/X vssd1 vssd1 vccd1 vccd1 hold537/A sky130_fd_sc_hd__nand2_1
X_17693_ _17693_/A _17693_/B _17693_/C vssd1 vssd1 vccd1 vccd1 _17699_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_159_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19432_ _21021_/A _19430_/Y _21025_/C vssd1 vssd1 vccd1 vccd1 _19523_/B sky130_fd_sc_hd__o21a_1
X_16644_ _16644_/A _16697_/B vssd1 vssd1 vccd1 vccd1 _16644_/Y sky130_fd_sc_hd__nand2_1
X_13856_ _13880_/A hold806/X vssd1 vssd1 vccd1 vccd1 hold807/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12807_ _12746_/X _12805_/X _14910_/B _12806_/X vssd1 vssd1 vccd1 vccd1 hold978/A
+ sky130_fd_sc_hd__o211a_1
X_19363_ _19364_/B _19364_/A vssd1 vssd1 vccd1 vccd1 _19363_/X sky130_fd_sc_hd__or2_1
XFILLER_0_97_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16575_ _16575_/A _16575_/B vssd1 vssd1 vccd1 vccd1 _16597_/A sky130_fd_sc_hd__nor2_1
X_13787_ _25761_/Q vssd1 vssd1 vccd1 vccd1 _18713_/B sky130_fd_sc_hd__inv_2
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18314_ _18312_/X _18269_/X _18313_/X vssd1 vssd1 vccd1 vccd1 _18315_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15526_ _15621_/A _16475_/B vssd1 vssd1 vccd1 vccd1 _15529_/A sky130_fd_sc_hd__nor2_1
X_12738_ _12548_/C _14120_/A _12737_/X vssd1 vssd1 vccd1 vccd1 _16702_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19294_ _19294_/A _19294_/B vssd1 vssd1 vccd1 vccd1 _19294_/Y sky130_fd_sc_hd__nand2_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15457_ _15458_/B _15458_/A vssd1 vssd1 vccd1 vccd1 _15459_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_155_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18245_ _21027_/B _21740_/A vssd1 vssd1 vccd1 vccd1 _21021_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12669_ _12671_/B vssd1 vssd1 vccd1 vccd1 _12674_/A sky130_fd_sc_hd__inv_2
XFILLER_0_143_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14408_ _14687_/B vssd1 vssd1 vccd1 vccd1 _14464_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15388_ _15388_/A _15388_/B vssd1 vssd1 vccd1 vccd1 _15389_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_143_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18176_ _18392_/A _18534_/A vssd1 vssd1 vccd1 vccd1 _18177_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17127_ _25597_/Q vssd1 vssd1 vccd1 vccd1 _20586_/B sky130_fd_sc_hd__inv_2
X_14339_ _14337_/Y hold324/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold325/A sky130_fd_sc_hd__a21oi_1
Xhold505 hold505/A vssd1 vssd1 vccd1 vccd1 hold505/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 hold516/A vssd1 vssd1 vccd1 vccd1 hold516/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold527 hold527/A vssd1 vssd1 vccd1 vccd1 hold527/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 hold538/A vssd1 vssd1 vccd1 vccd1 hold538/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17058_ _19659_/A _17058_/B vssd1 vssd1 vccd1 vccd1 _17512_/A sky130_fd_sc_hd__xor2_4
Xhold549 hold549/A vssd1 vssd1 vccd1 vccd1 hold549/X sky130_fd_sc_hd__dlygate4sd3_1
X_16009_ _16007_/Y _16008_/Y _15805_/X vssd1 vssd1 vccd1 vccd1 hold799/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1205 _25078_/Q vssd1 vssd1 vccd1 vccd1 _18270_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 _13276_/X vssd1 vssd1 vccd1 vccd1 _25098_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 _16983_/Y vssd1 vssd1 vccd1 vccd1 _25580_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1238 _25729_/Q vssd1 vssd1 vccd1 vccd1 _19396_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 _16894_/Y vssd1 vssd1 vccd1 vccd1 _25567_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20971_ _20973_/B vssd1 vssd1 vccd1 vccd1 _20972_/B sky130_fd_sc_hd__inv_2
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22710_ _22709_/A _22454_/X _22709_/B vssd1 vssd1 vccd1 vccd1 _22711_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23690_ hold2186/X hold2163/X _23754_/S vssd1 vssd1 vccd1 vccd1 _23691_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_73_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22641_ _18897_/A _25834_/Q _22639_/Y _22640_/Y vssd1 vssd1 vccd1 vccd1 _22642_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25360_ _26190_/CLK hold46/X vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__dfxtp_1
X_22572_ _23087_/B _22941_/B vssd1 vssd1 vccd1 vccd1 _22574_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24311_ hold2175/X _26169_/Q _24356_/S vssd1 vssd1 vccd1 vccd1 _24311_/X sky130_fd_sc_hd__mux2_1
X_21523_ _21523_/A _21523_/B vssd1 vssd1 vccd1 vccd1 _21524_/A sky130_fd_sc_hd__nand2_1
X_25291_ _26244_/CLK hold166/X vssd1 vssd1 vccd1 vccd1 hold164/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24242_ _24242_/A vssd1 vssd1 vccd1 vccd1 _26146_/D sky130_fd_sc_hd__clkbuf_1
X_21454_ _26324_/Q _21228_/X hold839/X vssd1 vssd1 vccd1 vccd1 _21457_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20405_ _20405_/A _22375_/B _20405_/C vssd1 vssd1 vccd1 vccd1 _20409_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_31_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24173_ _24173_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24174_/A sky130_fd_sc_hd__and2_1
XFILLER_0_189_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21385_ _21385_/A _21433_/A vssd1 vssd1 vccd1 vccd1 _21387_/A sky130_fd_sc_hd__nand2_1
X_23124_ _23188_/A _23124_/B vssd1 vssd1 vccd1 vccd1 _23124_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20336_ _21172_/B _21498_/A vssd1 vssd1 vccd1 vccd1 _20338_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_113_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23055_ _23055_/A _23055_/B vssd1 vssd1 vccd1 vccd1 _23057_/A sky130_fd_sc_hd__nand2_1
X_20267_ _21042_/A _20267_/B _20266_/X vssd1 vssd1 vccd1 vccd1 _20268_/B sky130_fd_sc_hd__or3b_1
X_22006_ _25801_/Q _22006_/B vssd1 vssd1 vccd1 vccd1 _22006_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_179_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20198_ _20196_/Y _20197_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _20198_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2440 _24988_/Q vssd1 vssd1 vccd1 vccd1 _12679_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2451 _26106_/Q vssd1 vssd1 vccd1 vccd1 hold2451/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2462 _15465_/Y vssd1 vssd1 vccd1 vccd1 _25455_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2473 _15575_/Y vssd1 vssd1 vccd1 vccd1 hold2473/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2484 _12677_/X vssd1 vssd1 vccd1 vccd1 _12678_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1750 _25420_/Q vssd1 vssd1 vccd1 vccd1 _14962_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2495 _26289_/Q vssd1 vssd1 vccd1 vccd1 hold2495/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1761 _25838_/Q vssd1 vssd1 vccd1 vccd1 _21757_/B sky130_fd_sc_hd__dlygate4sd3_1
X_23957_ _23957_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23958_/A sky130_fd_sc_hd__and2_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1772 _22385_/Y vssd1 vssd1 vccd1 vccd1 _25859_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1783 _22486_/Y vssd1 vssd1 vccd1 vccd1 _25863_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1794 _25884_/Q vssd1 vssd1 vccd1 vccd1 _22920_/B sky130_fd_sc_hd__clkbuf_2
X_13710_ _13823_/A _13710_/B vssd1 vssd1 vccd1 vccd1 _13710_/Y sky130_fd_sc_hd__nand2_1
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22908_ _22908_/A _22908_/B vssd1 vssd1 vccd1 vccd1 _22909_/B sky130_fd_sc_hd__nand2_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14690_ _15839_/A _25981_/Q vssd1 vssd1 vccd1 vccd1 _21722_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_86_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23888_ _23888_/A vssd1 vssd1 vccd1 vccd1 _26033_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13641_ _13636_/Y _13640_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold836/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22839_ _22837_/X _22838_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22839_/Y sky130_fd_sc_hd__a21oi_1
X_25627_ _25716_/CLK _25627_/D vssd1 vssd1 vccd1 vccd1 _25627_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_116_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _16360_/A vssd1 vssd1 vccd1 vccd1 _16378_/A sky130_fd_sc_hd__inv_2
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25558_ _25878_/CLK _25558_/D vssd1 vssd1 vccd1 vccd1 _25558_/Q sky130_fd_sc_hd__dfxtp_1
X_13572_ _13567_/Y _13571_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold850/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _15311_/A _15326_/B vssd1 vssd1 vccd1 vccd1 _15311_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _15839_/B vssd1 vssd1 vccd1 vccd1 _22829_/A sky130_fd_sc_hd__clkinv_4
X_24509_ _24509_/A vssd1 vssd1 vccd1 vccd1 _26233_/D sky130_fd_sc_hd__clkbuf_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16291_ _16289_/X hold702/X _16076_/X vssd1 vssd1 vccd1 vccd1 hold703/A sky130_fd_sc_hd__a21oi_1
X_25489_ _25933_/CLK _25489_/D vssd1 vssd1 vccd1 vccd1 _25489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15242_ _22631_/B _15242_/B vssd1 vssd1 vccd1 vccd1 _22628_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_152_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18030_ _18611_/A _18034_/B vssd1 vssd1 vccd1 vccd1 _18032_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15173_ _22529_/B _15173_/B vssd1 vssd1 vccd1 vccd1 _22526_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_23_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14124_ _14118_/Y _14123_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold822/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_162_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19981_ _19981_/A _19989_/B vssd1 vssd1 vccd1 vccd1 _19983_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14055_ _14061_/A _14055_/B vssd1 vssd1 vccd1 vccd1 _14055_/Y sky130_fd_sc_hd__nand2_1
X_18932_ _18952_/A _25772_/Q _18952_/C vssd1 vssd1 vccd1 vccd1 _18933_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_24_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13006_ _17550_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13006_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18863_ _18861_/Y _18862_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25687_/D sky130_fd_sc_hd__a21oi_1
X_17814_ _17814_/A _17814_/B _17814_/C vssd1 vssd1 vccd1 vccd1 _22280_/A sky130_fd_sc_hd__nand3_2
X_18794_ _18794_/A _18794_/B _18794_/C vssd1 vssd1 vccd1 vccd1 _22515_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17745_ _17771_/A _17745_/B _17830_/A vssd1 vssd1 vccd1 vccd1 _17760_/B sky130_fd_sc_hd__nand3_1
X_14957_ _14965_/A _14946_/A _14946_/B vssd1 vssd1 vccd1 vccd1 _14959_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_159_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13908_ _18073_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13908_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_89_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17676_ _17707_/B _25903_/Q _17685_/C vssd1 vssd1 vccd1 vccd1 _17679_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_159_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14888_ _25859_/Q _12527_/A _15076_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14888_/X
+ sky130_fd_sc_hd__a22o_1
X_19415_ _19412_/Y _19415_/B _19980_/B vssd1 vssd1 vccd1 vccd1 _19415_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_186_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16627_ _16627_/A _16627_/B vssd1 vssd1 vccd1 vccd1 _16628_/B sky130_fd_sc_hd__nand2_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13839_ _25769_/Q vssd1 vssd1 vccd1 vccd1 _18873_/B sky130_fd_sc_hd__inv_2
XFILLER_0_147_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19346_ _20855_/A _21835_/B _25604_/Q vssd1 vssd1 vccd1 vccd1 _20860_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_70_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16558_ _16698_/A hold904/X vssd1 vssd1 vccd1 vccd1 _16558_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15509_ _22914_/B _15509_/B vssd1 vssd1 vccd1 vccd1 _22911_/B sky130_fd_sc_hd__xor2_1
X_19277_ _20662_/A _19275_/Y _20666_/C vssd1 vssd1 vccd1 vccd1 _19364_/B sky130_fd_sc_hd__o21a_1
X_16489_ _16489_/A _16489_/B vssd1 vssd1 vccd1 vccd1 _16490_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_116_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18228_ _19038_/A _18228_/B vssd1 vssd1 vccd1 vccd1 _18228_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18159_ _18159_/A _18159_/B _25782_/Q vssd1 vssd1 vccd1 vccd1 _20317_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_13_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold302 hold302/A vssd1 vssd1 vccd1 vccd1 hold302/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold313 hold313/A vssd1 vssd1 vccd1 vccd1 hold313/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 hold324/A vssd1 vssd1 vccd1 vccd1 hold324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 hold335/A vssd1 vssd1 vccd1 vccd1 hold335/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21170_ _21577_/C _21627_/C vssd1 vssd1 vccd1 vccd1 _21172_/A sky130_fd_sc_hd__nand2_1
Xhold346 hold346/A vssd1 vssd1 vccd1 vccd1 hold346/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold357 hold357/A vssd1 vssd1 vccd1 vccd1 hold357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 hold368/A vssd1 vssd1 vccd1 vccd1 hold368/X sky130_fd_sc_hd__dlygate4sd3_1
X_20121_ _20121_/A _20121_/B vssd1 vssd1 vccd1 vccd1 _20122_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold379 hold379/A vssd1 vssd1 vccd1 vccd1 hold379/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20052_ _20052_/A _20052_/B vssd1 vssd1 vccd1 vccd1 _21693_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_102_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 _12880_/X vssd1 vssd1 vccd1 vccd1 _25027_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24860_ _15656_/A _15673_/B _24860_/S vssd1 vssd1 vccd1 vccd1 _24860_/X sky130_fd_sc_hd__mux2_1
Xhold1013 _25122_/Q vssd1 vssd1 vccd1 vccd1 _19033_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1024 _12919_/X vssd1 vssd1 vccd1 vccd1 _25034_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 _25073_/Q vssd1 vssd1 vccd1 vccd1 _18144_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23811_ _23811_/A vssd1 vssd1 vccd1 vccd1 _26008_/D sky130_fd_sc_hd__clkbuf_1
Xhold1046 _12875_/X vssd1 vssd1 vccd1 vccd1 _25026_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1057 _25009_/Q vssd1 vssd1 vccd1 vccd1 _17122_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1068 _12812_/X vssd1 vssd1 vccd1 vccd1 _25014_/D sky130_fd_sc_hd__dlygate4sd3_1
X_24791_ _24791_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24792_/A sky130_fd_sc_hd__and2_1
Xhold1079 _25040_/Q vssd1 vssd1 vccd1 vccd1 _17471_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23742_ _14733_/B _25986_/Q _23754_/S vssd1 vssd1 vccd1 vccd1 _23742_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_68_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20954_ _20954_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _20960_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23673_ _23673_/A vssd1 vssd1 vccd1 vccd1 _25963_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20885_ _20885_/A _25861_/Q vssd1 vssd1 vccd1 vccd1 _20889_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_166_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25412_ _25860_/CLK _25412_/D vssd1 vssd1 vccd1 vccd1 _25412_/Q sky130_fd_sc_hd__dfxtp_1
X_22624_ _22974_/B _23120_/B vssd1 vssd1 vccd1 vccd1 _22625_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_119_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25343_ _26298_/CLK hold346/X vssd1 vssd1 vccd1 vccd1 hold344/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22555_ _22555_/A _22555_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22557_/A sky130_fd_sc_hd__or3_1
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21506_ _21636_/A _21506_/B _21505_/X vssd1 vssd1 vccd1 vccd1 _21507_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_107_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25274_ _26231_/CLK hold208/X vssd1 vssd1 vccd1 vccd1 hold206/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22486_ _22484_/X _22485_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22486_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24225_ hold2318/X hold2263/X _24279_/S vssd1 vssd1 vccd1 vccd1 _24226_/A sky130_fd_sc_hd__mux2_1
X_21437_ _21437_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21442_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24156_ _24156_/A vssd1 vssd1 vccd1 vccd1 _26118_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21368_ _21368_/A _21368_/B _21368_/C vssd1 vssd1 vccd1 vccd1 _21372_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_102_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23107_ _23107_/A _23187_/B vssd1 vssd1 vccd1 vccd1 _23107_/Y sky130_fd_sc_hd__nand2_1
X_20319_ _20319_/A _20319_/B vssd1 vssd1 vccd1 vccd1 _21169_/C sky130_fd_sc_hd__nand2_4
X_24087_ _24087_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24088_/A sky130_fd_sc_hd__and2_1
Xhold880 hold880/A vssd1 vssd1 vccd1 vccd1 hold880/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21299_ _21662_/B _21707_/C vssd1 vssd1 vccd1 vccd1 _21302_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_102_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold891 hold891/A vssd1 vssd1 vccd1 vccd1 hold891/X sky130_fd_sc_hd__dlygate4sd3_1
X_23038_ _23036_/X _23037_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _23038_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15860_ _15858_/X _15859_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _15860_/X sky130_fd_sc_hd__a21o_1
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2270 _26097_/Q vssd1 vssd1 vccd1 vccd1 hold2270/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14811_ _25850_/Q _13466_/A _14810_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14812_/A
+ sky130_fd_sc_hd__a22o_1
Xhold2281 _26117_/Q vssd1 vssd1 vccd1 vccd1 hold2281/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_189_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2292 _25945_/Q vssd1 vssd1 vccd1 vccd1 hold2292/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _26043_/Q _25979_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15792_/A sky130_fd_sc_hd__mux2_1
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24989_ _24990_/CLK _24989_/D vssd1 vssd1 vccd1 vccd1 _24989_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1580 _25773_/Q vssd1 vssd1 vccd1 vccd1 _19997_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _17527_/X _17528_/X _17529_/X vssd1 vssd1 vccd1 vccd1 _17531_/A sky130_fd_sc_hd__a21o_1
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14742_ _14739_/Y _14740_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14742_/Y sky130_fd_sc_hd__a21oi_1
Xhold1591 _22904_/Y vssd1 vssd1 vccd1 vccd1 _25883_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14673_ _14688_/A hold347/X vssd1 vssd1 vccd1 vccd1 hold348/A sky130_fd_sc_hd__nand2_1
X_17461_ _17459_/Y _17460_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _17461_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_192_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _26249_/CLK sky130_fd_sc_hd__clkbuf_16
X_19200_ _19452_/A _19200_/B vssd1 vssd1 vccd1 vccd1 _19200_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16412_ _16413_/B _16413_/A vssd1 vssd1 vccd1 vccd1 _16441_/A sky130_fd_sc_hd__or2_1
XFILLER_0_168_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13624_ _13642_/A hold494/X vssd1 vssd1 vccd1 vccd1 hold495/A sky130_fd_sc_hd__nand2_1
XFILLER_0_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17392_ _17652_/A _17392_/B vssd1 vssd1 vccd1 vccd1 _17392_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_27_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19131_ _20986_/A vssd1 vssd1 vccd1 vccd1 _19131_/X sky130_fd_sc_hd__buf_12
X_16343_ _17568_/A vssd1 vssd1 vccd1 vccd1 _16343_/X sky130_fd_sc_hd__buf_6
X_13555_ _25724_/Q vssd1 vssd1 vccd1 vccd1 _17989_/B sky130_fd_sc_hd__inv_2
XFILLER_0_6_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12506_ _24969_/Q _24968_/Q _24967_/Q _24966_/Q vssd1 vssd1 vccd1 vccd1 _12507_/D
+ sky130_fd_sc_hd__or4_1
X_16274_ _16274_/A _16274_/B vssd1 vssd1 vccd1 vccd1 _16279_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_164_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19062_ _19060_/X _18879_/X _19061_/X vssd1 vssd1 vccd1 vccd1 _19063_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_82_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13486_ _13522_/A hold413/X vssd1 vssd1 vccd1 vccd1 hold414/A sky130_fd_sc_hd__nand2_1
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15225_ _22606_/B _15225_/B vssd1 vssd1 vccd1 vccd1 _22603_/B sky130_fd_sc_hd__xor2_1
X_18013_ _19176_/B _25651_/Q vssd1 vssd1 vccd1 vccd1 _18017_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_112_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15156_ _15621_/A _15156_/B vssd1 vssd1 vccd1 vccd1 _15159_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14107_ _25812_/Q vssd1 vssd1 vccd1 vccd1 _18450_/B sky130_fd_sc_hd__inv_2
XFILLER_0_26_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15087_ _15073_/A _15085_/Y _15086_/X vssd1 vssd1 vccd1 vccd1 _15089_/A sky130_fd_sc_hd__a21bo_1
X_19964_ _19975_/A _19964_/B vssd1 vssd1 vccd1 vccd1 _19964_/Y sky130_fd_sc_hd__nand2_1
X_14038_ hold711/X _14036_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold712/A sky130_fd_sc_hd__a21oi_1
X_18915_ _18915_/A _18915_/B _18915_/C vssd1 vssd1 vccd1 vccd1 _22667_/A sky130_fd_sc_hd__nand3_2
X_19895_ _26268_/Q _19134_/X hold677/X vssd1 vssd1 vccd1 vccd1 _19896_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_38_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18846_ _25640_/Q _22590_/B vssd1 vssd1 vccd1 vccd1 _18847_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18777_ _18966_/A _19017_/B vssd1 vssd1 vccd1 vccd1 _18778_/B sky130_fd_sc_hd__xnor2_1
X_15989_ _15989_/A _15999_/B vssd1 vssd1 vccd1 vccd1 _15989_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_179_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17728_ _17728_/A _17728_/B _17728_/C vssd1 vssd1 vccd1 vccd1 _17729_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_136_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17659_ _21749_/A vssd1 vssd1 vccd1 vccd1 _19089_/B sky130_fd_sc_hd__inv_2
XFILLER_0_33_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_183_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _25740_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20670_ _20670_/A _20670_/B vssd1 vssd1 vccd1 vccd1 _21371_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19329_ _19328_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19330_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_162_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22340_ _22325_/X _22339_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _22340_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22271_ _22272_/B _22272_/A vssd1 vssd1 vccd1 vccd1 _22273_/A sky130_fd_sc_hd__or2_1
XFILLER_0_60_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24010_ _24010_/A vssd1 vssd1 vccd1 vccd1 _26071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold110 hold110/A vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
X_21222_ _21222_/A _21222_/B _21222_/C vssd1 vssd1 vccd1 vccd1 _21226_/A sky130_fd_sc_hd__nand3_1
Xhold121 hold121/A vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 hold132/A vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold143 hold143/A vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 hold154/A vssd1 vssd1 vccd1 vccd1 hold154/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 hold165/A vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
X_21153_ _21153_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21153_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold176 hold176/A vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 hold187/A vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 hold198/A vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__dlygate4sd3_1
X_20104_ _20106_/C vssd1 vssd1 vccd1 vccd1 _20105_/B sky130_fd_sc_hd__inv_2
X_25961_ _26042_/CLK _25961_/D vssd1 vssd1 vccd1 vccd1 _25961_/Q sky130_fd_sc_hd__dfxtp_1
X_21084_ _21577_/C _21529_/C vssd1 vssd1 vccd1 vccd1 _21086_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24912_ _24957_/S _24912_/B vssd1 vssd1 vccd1 vccd1 _24912_/Y sky130_fd_sc_hd__nor2_1
X_20035_ _26277_/Q _19134_/X hold722/X vssd1 vssd1 vccd1 vccd1 _20038_/B sky130_fd_sc_hd__a21oi_1
X_25892_ _25898_/CLK _25892_/D vssd1 vssd1 vccd1 vccd1 _25892_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24843_ _24841_/X _24842_/X _24858_/S vssd1 vssd1 vccd1 vccd1 _24843_/X sky130_fd_sc_hd__mux2_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24774_ _24774_/A vssd1 vssd1 vccd1 vccd1 _26319_/D sky130_fd_sc_hd__clkbuf_1
X_21986_ _21986_/A _22740_/B vssd1 vssd1 vccd1 vccd1 _21987_/B sky130_fd_sc_hd__nand2_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23725_ _23725_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23726_/A sky130_fd_sc_hd__and2_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20937_ _20940_/A _20940_/C vssd1 vssd1 vccd1 vccd1 _20938_/A sky130_fd_sc_hd__nand2_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_174_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _26234_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23656_ hold2092/X _25958_/Q _23677_/S vssd1 vssd1 vccd1 vccd1 _23656_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20868_ _20868_/A _20868_/B _21403_/B vssd1 vssd1 vccd1 vccd1 _20872_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22607_ _22606_/A _22454_/X _22606_/B vssd1 vssd1 vccd1 vccd1 _22608_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23587_ _23587_/A _23587_/B _23587_/C vssd1 vssd1 vccd1 vccd1 _23593_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_153_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20799_ _20799_/A _20799_/B vssd1 vssd1 vccd1 vccd1 _21693_/B sky130_fd_sc_hd__nand2_8
XFILLER_0_91_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25326_ _25711_/CLK hold112/X vssd1 vssd1 vccd1 vccd1 hold110/A sky130_fd_sc_hd__dfxtp_1
X_13340_ _13315_/X _13338_/X _13300_/X _13339_/X vssd1 vssd1 vccd1 vccd1 _13340_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22538_ _22538_/A _25894_/Q vssd1 vssd1 vccd1 vccd1 _22538_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25257_ _25257_/CLK hold427/X vssd1 vssd1 vccd1 vccd1 hold425/A sky130_fd_sc_hd__dfxtp_1
X_13271_ _13271_/A vssd1 vssd1 vccd1 vccd1 _19488_/A sky130_fd_sc_hd__buf_4
X_22469_ _22469_/A _22469_/B vssd1 vssd1 vccd1 vccd1 _23024_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_121_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15010_ _15010_/A _15010_/B vssd1 vssd1 vccd1 vccd1 _15010_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24208_ _24208_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24209_/A sky130_fd_sc_hd__and2_1
X_25188_ _25770_/CLK hold628/X vssd1 vssd1 vccd1 vccd1 hold626/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24139_ hold1972/X _26113_/Q _24203_/S vssd1 vssd1 vccd1 vccd1 _24139_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16961_ _16959_/X _16711_/A _16960_/Y _25898_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16962_/A sky130_fd_sc_hd__a32o_1
X_18700_ _18698_/X _18269_/X _18699_/X vssd1 vssd1 vccd1 vccd1 _18701_/A sky130_fd_sc_hd__a21o_1
X_15912_ _15910_/X _15911_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _15912_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_95_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19680_ _19672_/X _19679_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19680_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_159_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16892_ _16892_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16892_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_21_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18631_ _18954_/A _25757_/Q vssd1 vssd1 vccd1 vccd1 _18633_/A sky130_fd_sc_hd__nand2_1
X_15843_ _15844_/B _15844_/A vssd1 vssd1 vccd1 vccd1 _15857_/B sky130_fd_sc_hd__or2_1
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18562_ _19659_/A vssd1 vssd1 vccd1 vccd1 _22237_/B sky130_fd_sc_hd__inv_2
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ _15774_/A _15774_/B vssd1 vssd1 vccd1 vccd1 _15775_/B sky130_fd_sc_hd__nand2_2
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ _12930_/X hold900/X _12917_/X _12985_/X vssd1 vssd1 vccd1 vccd1 hold901/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17513_ _17513_/A _17513_/B vssd1 vssd1 vccd1 vccd1 _17513_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14725_ _15543_/B vssd1 vssd1 vccd1 vccd1 _15778_/B sky130_fd_sc_hd__buf_8
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_165_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _26292_/CLK sky130_fd_sc_hd__clkbuf_16
X_18493_ _18698_/A _18838_/A vssd1 vssd1 vccd1 vccd1 _18494_/B sky130_fd_sc_hd__xnor2_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _17444_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17444_/Y sky130_fd_sc_hd__nand2_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14656_ _14654_/Y hold168/X _14646_/X vssd1 vssd1 vccd1 vccd1 hold169/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13607_ _18052_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13607_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_184_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17375_ _17375_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17375_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_32_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14587_ _14584_/Y hold210/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold211/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19114_ _19114_/A vssd1 vssd1 vccd1 vccd1 _19115_/C sky130_fd_sc_hd__inv_2
X_16326_ _16473_/A hold873/X vssd1 vssd1 vccd1 vccd1 _16326_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_131_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13538_ _17858_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13538_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_125_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19045_ _19045_/A _19045_/B vssd1 vssd1 vccd1 vccd1 _19046_/B sky130_fd_sc_hd__xnor2_1
X_16257_ _16473_/A hold889/X vssd1 vssd1 vccd1 vccd1 _16257_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_153_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13469_ _25710_/Q vssd1 vssd1 vccd1 vccd1 _13470_/A sky130_fd_sc_hd__inv_2
XFILLER_0_2_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15208_ _22580_/B _15208_/B vssd1 vssd1 vccd1 vccd1 _22577_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_152_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16188_ _16181_/A _16167_/A _16180_/B vssd1 vssd1 vccd1 vccd1 _16188_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_140_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15139_ _15776_/B vssd1 vssd1 vccd1 vccd1 _16369_/B sky130_fd_sc_hd__buf_6
XFILLER_0_142_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19947_ _19947_/A _19980_/B _19947_/C vssd1 vssd1 vccd1 vccd1 _19947_/X sky130_fd_sc_hd__and3_1
XFILLER_0_10_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19878_ _19975_/A _19878_/B vssd1 vssd1 vccd1 vccd1 _19878_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_156_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18829_ _18951_/A _18833_/B vssd1 vssd1 vccd1 vccd1 _18831_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_179_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21840_ _21840_/A _21840_/B vssd1 vssd1 vccd1 vccd1 _21841_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21771_ _23072_/A vssd1 vssd1 vccd1 vccd1 _23071_/A sky130_fd_sc_hd__inv_2
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_156_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _26303_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23510_ _24940_/S hold266/A _23509_/X vssd1 vssd1 vccd1 vccd1 _23510_/Y sky130_fd_sc_hd__o21ai_1
X_20722_ _21384_/C _21661_/B vssd1 vssd1 vccd1 vccd1 _20725_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_172_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24490_ _24490_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24491_/A sky130_fd_sc_hd__and2_1
XFILLER_0_65_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23441_ _24956_/S hold200/A _23440_/X vssd1 vssd1 vccd1 vccd1 _23441_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_175_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20653_ _20653_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20658_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26160_ _26164_/CLK _26160_/D vssd1 vssd1 vccd1 vccd1 _26160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23372_ _23372_/A _23372_/B vssd1 vssd1 vccd1 vccd1 _23372_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_18_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20584_ _20582_/Y _20583_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _20584_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25111_ _26198_/CLK _25111_/D vssd1 vssd1 vccd1 vccd1 _25111_/Q sky130_fd_sc_hd__dfxtp_1
X_22323_ _22323_/A _22387_/B vssd1 vssd1 vccd1 vccd1 _22323_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_144_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26091_ _26221_/CLK _26091_/D vssd1 vssd1 vccd1 vccd1 _26091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25042_ _26216_/CLK _25042_/D vssd1 vssd1 vccd1 vccd1 _25042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22254_ _22254_/A _22254_/B vssd1 vssd1 vccd1 vccd1 _23007_/B sky130_fd_sc_hd__nand2_4
X_21205_ _21636_/A _21205_/B _21204_/X vssd1 vssd1 vccd1 vccd1 _21206_/B sky130_fd_sc_hd__or3b_1
X_22185_ _22185_/A _22185_/B vssd1 vssd1 vccd1 vccd1 _22840_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_108_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21136_ _21136_/A _21136_/B _21136_/C vssd1 vssd1 vccd1 vccd1 _21137_/B sky130_fd_sc_hd__nand3_1
X_25944_ _26009_/CLK _25944_/D vssd1 vssd1 vccd1 vccd1 _25944_/Q sky130_fd_sc_hd__dfxtp_1
X_21067_ _26306_/Q hold512/X vssd1 vssd1 vccd1 vccd1 _21067_/Y sky130_fd_sc_hd__nand2_1
X_20018_ _20018_/A _20018_/B _20018_/C vssd1 vssd1 vccd1 vccd1 _20019_/B sky130_fd_sc_hd__nand3_1
X_25875_ _25875_/CLK _25875_/D vssd1 vssd1 vccd1 vccd1 _25875_/Q sky130_fd_sc_hd__dfxtp_2
X_12840_ _14260_/A vssd1 vssd1 vccd1 vccd1 _12840_/X sky130_fd_sc_hd__clkbuf_8
X_24826_ hold2366/X _26337_/Q _24835_/S vssd1 vssd1 vccd1 vccd1 _24826_/X sky130_fd_sc_hd__mux2_1
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12771_ hold960/X _14264_/A vssd1 vssd1 vccd1 vccd1 _12771_/X sky130_fd_sc_hd__or2_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21969_ _21967_/X _14270_/A _21968_/Y _14768_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _21970_/A sky130_fd_sc_hd__a32o_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24757_ hold2730/X _26314_/Q _24817_/S vssd1 vssd1 vccd1 vccd1 _24757_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_147_clk clkbuf_4_11__f_clk/X vssd1 vssd1 vccd1 vccd1 _26190_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14510_ _14525_/A hold89/X vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__nand2_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15490_ _22896_/B _15490_/B vssd1 vssd1 vccd1 vccd1 _22893_/B sky130_fd_sc_hd__xor2_1
X_23708_ hold1957/X _25975_/Q _23754_/S vssd1 vssd1 vccd1 vccd1 _23708_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24688_ _24688_/A vssd1 vssd1 vccd1 vccd1 _26291_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23639_ _23639_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23640_/A sky130_fd_sc_hd__and2_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ _14465_/A hold113/X vssd1 vssd1 vccd1 vccd1 hold114/A sky130_fd_sc_hd__nand2_1
XFILLER_0_83_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14372_ _14370_/Y hold219/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold220/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17160_ _17434_/A _17160_/B vssd1 vssd1 vccd1 vccd1 _17160_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16111_ _22343_/B _16691_/B vssd1 vssd1 vccd1 vccd1 _16113_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13323_ _26317_/Q _19602_/A vssd1 vssd1 vccd1 vccd1 _14617_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25309_ _26139_/CLK hold115/X vssd1 vssd1 vccd1 vccd1 hold113/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26289_ _26289_/CLK _26289_/D vssd1 vssd1 vccd1 vccd1 _26289_/Q sky130_fd_sc_hd__dfxtp_2
X_17091_ _17448_/A _17526_/A vssd1 vssd1 vccd1 vccd1 _17092_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_165_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16042_ _16042_/A _16052_/B vssd1 vssd1 vccd1 vccd1 _16042_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_122_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13254_ _26306_/Q _19444_/A vssd1 vssd1 vccd1 vccd1 _14581_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_33_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13185_ _26167_/Q _13065_/X _13184_/X vssd1 vssd1 vccd1 vccd1 _13185_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19801_ _19798_/Y _19801_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19801_/X sky130_fd_sc_hd__and3b_1
X_17993_ _19331_/A vssd1 vssd1 vccd1 vccd1 _21801_/B sky130_fd_sc_hd__inv_2
X_19732_ _19749_/B _19821_/B vssd1 vssd1 vccd1 vccd1 _19734_/A sky130_fd_sc_hd__xnor2_1
X_16944_ _22145_/B _16949_/B vssd1 vssd1 vccd1 vccd1 _16946_/B sky130_fd_sc_hd__nand2_1
X_19663_ _19664_/B _19664_/A vssd1 vssd1 vccd1 vccd1 _19663_/X sky130_fd_sc_hd__or2_1
X_16875_ _16876_/B _16876_/A vssd1 vssd1 vccd1 vccd1 _16875_/X sky130_fd_sc_hd__or2_1
X_18614_ _20281_/B _22299_/A vssd1 vssd1 vccd1 vccd1 _20272_/A sky130_fd_sc_hd__nand2_2
X_15826_ _15826_/A _15828_/A vssd1 vssd1 vccd1 vccd1 _15827_/B sky130_fd_sc_hd__nor2_1
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19594_ _19592_/X _19593_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19594_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18545_ _25881_/Q _22207_/A vssd1 vssd1 vccd1 vccd1 _18553_/A sky130_fd_sc_hd__or2_2
X_15757_ _23140_/B _15812_/B vssd1 vssd1 vccd1 vccd1 _16651_/B sky130_fd_sc_hd__nand2_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_138_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _25750_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _17500_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12969_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14708_ _14907_/B vssd1 vssd1 vccd1 vccd1 _14916_/A sky130_fd_sc_hd__inv_2
X_18476_ _18474_/X _18269_/X _18475_/X vssd1 vssd1 vccd1 vccd1 _18477_/A sky130_fd_sc_hd__a21o_1
X_15688_ _15690_/B _16930_/A vssd1 vssd1 vccd1 vccd1 _15689_/A sky130_fd_sc_hd__nor2_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17427_ _17467_/A _17427_/B vssd1 vssd1 vccd1 vccd1 _17427_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14639_ _14645_/A hold32/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17358_ _25615_/Q vssd1 vssd1 vccd1 vccd1 _21157_/B sky130_fd_sc_hd__inv_2
XFILLER_0_71_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16309_ _16309_/A _16309_/B vssd1 vssd1 vccd1 vccd1 _16334_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17289_ _20994_/B _25865_/Q _21019_/B vssd1 vssd1 vccd1 vccd1 _17290_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_42_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19028_ _19028_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _19028_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23990_ _23990_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23991_/A sky130_fd_sc_hd__and2_1
X_22941_ _23090_/A _22941_/B vssd1 vssd1 vccd1 vccd1 _22942_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22872_ _22937_/A _22872_/B vssd1 vssd1 vccd1 vccd1 _22872_/Y sky130_fd_sc_hd__nand2_1
X_25660_ _26292_/CLK _25660_/D vssd1 vssd1 vccd1 vccd1 _25660_/Q sky130_fd_sc_hd__dfxtp_1
X_21823_ _21823_/A _21823_/B vssd1 vssd1 vccd1 vccd1 _22926_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24611_ _24611_/A vssd1 vssd1 vccd1 vccd1 _26266_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_129_clk clkbuf_4_14__f_clk/X vssd1 vssd1 vccd1 vccd1 _26336_/CLK sky130_fd_sc_hd__clkbuf_16
X_25591_ _26112_/CLK _25591_/D vssd1 vssd1 vccd1 vccd1 _25591_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_92_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24542_ _24542_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24543_/A sky130_fd_sc_hd__and2_1
X_21754_ _21754_/A _21754_/B _22745_/A vssd1 vssd1 vccd1 vccd1 _21754_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20705_ _25856_/Q _20705_/B _20705_/C vssd1 vssd1 vccd1 vccd1 _20708_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_175_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24473_ _24473_/A vssd1 vssd1 vccd1 vccd1 _26221_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21685_ _21685_/A _21685_/B vssd1 vssd1 vccd1 vccd1 _21686_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26212_ _26339_/CLK _26212_/D vssd1 vssd1 vccd1 vccd1 _26212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23424_ _23421_/Y _23423_/Y _24946_/A vssd1 vssd1 vccd1 vccd1 _23424_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20636_ _20639_/A _20639_/C vssd1 vssd1 vccd1 vccd1 _20637_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_110_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26143_ _26263_/CLK _26143_/D vssd1 vssd1 vccd1 vccd1 _26143_/Q sky130_fd_sc_hd__dfxtp_1
X_23355_ _23356_/B _23356_/A vssd1 vssd1 vccd1 vccd1 _23360_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_145_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20567_ _20567_/A _20567_/B vssd1 vssd1 vccd1 vccd1 _21596_/A sky130_fd_sc_hd__nand2_4
X_22306_ _22759_/A _22907_/B vssd1 vssd1 vccd1 vccd1 _22317_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26074_ _26079_/CLK _26074_/D vssd1 vssd1 vccd1 vccd1 _26074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23286_ _23307_/A _23293_/B vssd1 vssd1 vccd1 vccd1 _23290_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_132_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20498_ _26289_/Q _20078_/X hold742/X vssd1 vssd1 vccd1 vccd1 _20501_/B sky130_fd_sc_hd__a21oi_1
X_25025_ _25604_/CLK hold984/X vssd1 vssd1 vccd1 vccd1 hold983/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22237_ _25818_/Q _22237_/B vssd1 vssd1 vccd1 vccd1 _22237_/Y sky130_fd_sc_hd__nor2_1
X_22168_ _22168_/A _23106_/A _22168_/C vssd1 vssd1 vccd1 vccd1 _22168_/Y sky130_fd_sc_hd__nand3_1
X_21119_ _21119_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _21124_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14990_ _14990_/A _14990_/B vssd1 vssd1 vccd1 vccd1 _14998_/B sky130_fd_sc_hd__nand2_1
X_22099_ _25877_/Q _22100_/A vssd1 vssd1 vccd1 vccd1 _22101_/A sky130_fd_sc_hd__or2_1
XFILLER_0_22_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25927_ _25939_/CLK _25927_/D vssd1 vssd1 vccd1 vccd1 _25927_/Q sky130_fd_sc_hd__dfxtp_1
X_13941_ _13941_/A _13941_/B vssd1 vssd1 vccd1 vccd1 _13941_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16660_ _16670_/A _16660_/B vssd1 vssd1 vccd1 vccd1 _16660_/Y sky130_fd_sc_hd__nand2_1
X_25858_ _25859_/CLK _25858_/D vssd1 vssd1 vccd1 vccd1 _25858_/Q sky130_fd_sc_hd__dfxtp_4
X_13872_ _13941_/A _13872_/B vssd1 vssd1 vccd1 vccd1 _13872_/Y sky130_fd_sc_hd__nand2_1
X_15611_ _15611_/A _15612_/A _15612_/B vssd1 vssd1 vccd1 vccd1 _15694_/A sky130_fd_sc_hd__and3_1
XFILLER_0_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24809_ _24809_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24810_/A sky130_fd_sc_hd__and2_1
X_12823_ _12746_/X _12820_/X _14910_/B _12822_/X vssd1 vssd1 vccd1 vccd1 _12823_/X
+ sky130_fd_sc_hd__o211a_1
X_16591_ _16596_/B _16591_/B vssd1 vssd1 vccd1 vccd1 _16592_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_158_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25789_ _25793_/CLK _25789_/D vssd1 vssd1 vccd1 vccd1 _25789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18330_ _18330_/A _21128_/A vssd1 vssd1 vccd1 vccd1 _18678_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_97_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15542_ _15542_/A vssd1 vssd1 vccd1 vccd1 _16498_/A sky130_fd_sc_hd__inv_2
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _26086_/Q _12748_/X _12753_/X vssd1 vssd1 vccd1 vccd1 _12754_/X sky130_fd_sc_hd__a21o_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18261_ _18261_/A _21072_/B _18261_/C vssd1 vssd1 vccd1 vccd1 _21053_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_182_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12685_ _12686_/B _12686_/A vssd1 vssd1 vccd1 vccd1 _12687_/A sky130_fd_sc_hd__or2_1
XFILLER_0_155_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15473_ _15473_/A _15812_/B vssd1 vssd1 vccd1 vccd1 _15474_/B sky130_fd_sc_hd__nand2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17212_ _17513_/A _17593_/A vssd1 vssd1 vccd1 vccd1 _17213_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14424_ _14422_/Y hold300/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold301/A sky130_fd_sc_hd__a21oi_1
X_18192_ _18192_/A _20349_/A vssd1 vssd1 vccd1 vccd1 _19081_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_37_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17143_ _25632_/Q vssd1 vssd1 vccd1 vccd1 _20439_/B sky130_fd_sc_hd__inv_2
XFILLER_0_141_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14355_ _14355_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14355_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_52_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13306_ _26186_/Q _13239_/X _13305_/X vssd1 vssd1 vccd1 vccd1 _13306_/X sky130_fd_sc_hd__a21o_1
X_14286_ _14687_/B vssd1 vssd1 vccd1 vccd1 _14343_/B sky130_fd_sc_hd__buf_6
XFILLER_0_52_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold709 hold709/A vssd1 vssd1 vccd1 vccd1 hold709/X sky130_fd_sc_hd__dlygate4sd3_1
X_17074_ _19673_/A _17074_/B vssd1 vssd1 vccd1 vccd1 _17519_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16025_ _16052_/A vssd1 vssd1 vccd1 vccd1 _16031_/B sky130_fd_sc_hd__inv_2
XFILLER_0_150_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13237_ _18557_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13237_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13168_ _18333_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13168_/X sky130_fd_sc_hd__or2_1
X_13099_ _26280_/Q _25649_/Q vssd1 vssd1 vccd1 vccd1 _14500_/A sky130_fd_sc_hd__xor2_1
X_17976_ _17976_/A _17976_/B vssd1 vssd1 vccd1 vccd1 _17977_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_100_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1409 _25551_/Q vssd1 vssd1 vccd1 vccd1 _16781_/B sky130_fd_sc_hd__buf_1
X_19715_ _19715_/A _20362_/B vssd1 vssd1 vccd1 vccd1 _19715_/Y sky130_fd_sc_hd__nor2_1
X_16927_ _16925_/Y _16926_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16927_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19646_ _20162_/A _19644_/Y _20167_/C vssd1 vssd1 vccd1 vccd1 _19734_/B sky130_fd_sc_hd__o21a_1
X_16858_ _16858_/A _16858_/B vssd1 vssd1 vccd1 vccd1 _16858_/Y sky130_fd_sc_hd__nand2_1
X_15809_ _26044_/Q _25980_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15810_/A sky130_fd_sc_hd__mux2_1
X_19577_ _19593_/B _19664_/B vssd1 vssd1 vccd1 vccd1 _19579_/A sky130_fd_sc_hd__xnor2_1
X_16789_ _16789_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16789_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_34_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18528_ _18528_/A _25752_/Q vssd1 vssd1 vccd1 vccd1 _18530_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18459_ _18457_/Y _18458_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25667_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_185_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21470_ _26325_/Q _21228_/X hold440/X vssd1 vssd1 vccd1 vccd1 _21473_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20421_ _26287_/Q hold686/X vssd1 vssd1 vccd1 vccd1 _20421_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_114_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23140_ _23188_/A _23140_/B vssd1 vssd1 vccd1 vccd1 _23140_/X sky130_fd_sc_hd__or2_1
XFILLER_0_113_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20352_ _20352_/A _25847_/Q vssd1 vssd1 vccd1 vccd1 _20358_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23071_ _23071_/A _23071_/B vssd1 vssd1 vccd1 vccd1 _23073_/A sky130_fd_sc_hd__nand2_1
X_20283_ _21482_/A vssd1 vssd1 vccd1 vccd1 _21481_/A sky130_fd_sc_hd__inv_2
XFILLER_0_178_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22022_ _23183_/A _22742_/B vssd1 vssd1 vccd1 vccd1 _22030_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2600 _26228_/Q vssd1 vssd1 vccd1 vccd1 hold2600/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2611 _26229_/Q vssd1 vssd1 vccd1 vccd1 hold2611/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2622 _25459_/Q vssd1 vssd1 vccd1 vccd1 _15528_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2633 _24642_/X vssd1 vssd1 vccd1 vccd1 _24643_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2644 _26315_/Q vssd1 vssd1 vccd1 vccd1 hold2644/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1910 _24287_/X vssd1 vssd1 vccd1 vccd1 _24288_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2655 _26321_/Q vssd1 vssd1 vccd1 vccd1 hold2655/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1921 _24308_/X vssd1 vssd1 vccd1 vccd1 _24309_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2666 _26320_/Q vssd1 vssd1 vccd1 vccd1 hold2666/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2677 _25911_/Q vssd1 vssd1 vccd1 vccd1 _23236_/A sky130_fd_sc_hd__buf_1
X_23973_ _23973_/A vssd1 vssd1 vccd1 vccd1 _26059_/D sky130_fd_sc_hd__clkbuf_1
Xhold1932 _26032_/Q vssd1 vssd1 vccd1 vccd1 hold1932/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1943 _26009_/Q vssd1 vssd1 vccd1 vccd1 hold1943/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2688 _26248_/Q vssd1 vssd1 vccd1 vccd1 hold2688/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2699 _23241_/Y vssd1 vssd1 vccd1 vccd1 _23245_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1954 _15025_/Y vssd1 vssd1 vccd1 vccd1 _25427_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1965 _25992_/Q vssd1 vssd1 vccd1 vccd1 _14797_/B sky130_fd_sc_hd__dlygate4sd3_1
X_25712_ _25712_/CLK hold607/X vssd1 vssd1 vccd1 vccd1 hold605/A sky130_fd_sc_hd__dfxtp_1
X_22924_ _22924_/A _23074_/A vssd1 vssd1 vccd1 vccd1 _22925_/B sky130_fd_sc_hd__nand2_1
Xhold1976 _26044_/Q vssd1 vssd1 vccd1 vccd1 hold1976/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1987 _26209_/Q vssd1 vssd1 vccd1 vccd1 hold1987/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1998 _24443_/X vssd1 vssd1 vccd1 vccd1 _24444_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25643_ _26148_/CLK _25643_/D vssd1 vssd1 vccd1 vccd1 _25643_/Q sky130_fd_sc_hd__dfxtp_2
X_22855_ _22937_/A _22855_/B vssd1 vssd1 vccd1 vccd1 _22855_/Y sky130_fd_sc_hd__nand2_1
X_21806_ _21806_/A _21806_/B vssd1 vssd1 vccd1 vccd1 _21807_/B sky130_fd_sc_hd__nand2_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25574_ _25893_/CLK _25574_/D vssd1 vssd1 vccd1 vccd1 _25574_/Q sky130_fd_sc_hd__dfxtp_1
X_22786_ _22786_/A vssd1 vssd1 vccd1 vccd1 _23099_/B sky130_fd_sc_hd__clkbuf_8
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24525_ _24525_/A vssd1 vssd1 vccd1 vccd1 _26238_/D sky130_fd_sc_hd__clkbuf_1
X_21737_ _21737_/A _25866_/Q vssd1 vssd1 vccd1 vccd1 _21737_/Y sky130_fd_sc_hd__nand2_1
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21668_ _21716_/A _21668_/B _21667_/X vssd1 vssd1 vccd1 vccd1 _21669_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24456_ _24456_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24457_/A sky130_fd_sc_hd__and2_1
XFILLER_0_47_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20619_ _21042_/A _20619_/B _20618_/X vssd1 vssd1 vccd1 vccd1 _20620_/B sky130_fd_sc_hd__or3b_1
X_23407_ _23395_/X _23406_/X _24949_/S vssd1 vssd1 vccd1 vccd1 _23407_/X sky130_fd_sc_hd__mux2_1
X_24387_ _24387_/A vssd1 vssd1 vccd1 vccd1 _26193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21599_ _21599_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21604_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_105_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14140_ _18551_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14140_/Y sky130_fd_sc_hd__nor2_1
X_23338_ _23336_/A hold952/X _23336_/B vssd1 vssd1 vccd1 vccd1 _23338_/X sky130_fd_sc_hd__a21o_1
X_26126_ _26130_/CLK _26126_/D vssd1 vssd1 vccd1 vccd1 _26126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14071_ _25806_/Q vssd1 vssd1 vccd1 vccd1 _18328_/B sky130_fd_sc_hd__inv_2
X_23269_ _23269_/A _23269_/B vssd1 vssd1 vccd1 vccd1 _23273_/A sky130_fd_sc_hd__nand2_1
X_26057_ _26057_/CLK _26057_/D vssd1 vssd1 vccd1 vccd1 _26057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13022_ _17572_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13022_/X sky130_fd_sc_hd__or2_1
X_25008_ _26221_/CLK _25008_/D vssd1 vssd1 vccd1 vccd1 _25008_/Q sky130_fd_sc_hd__dfxtp_1
X_17830_ _17830_/A _23203_/B vssd1 vssd1 vccd1 vccd1 _17831_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17761_ _18019_/B _17761_/B vssd1 vssd1 vccd1 vccd1 _17775_/A sky130_fd_sc_hd__nand2_2
X_14973_ _14973_/A _14973_/B vssd1 vssd1 vccd1 vccd1 _14982_/A sky130_fd_sc_hd__nand2_1
X_19500_ _26240_/Q _19483_/X hold835/X vssd1 vssd1 vccd1 vccd1 _19500_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16712_ _16712_/A _16712_/B vssd1 vssd1 vccd1 vccd1 _16712_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13924_ hold390/X _13923_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold391/A sky130_fd_sc_hd__a21oi_1
X_17692_ _17692_/A _17692_/B _17692_/C vssd1 vssd1 vccd1 vccd1 _17693_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_18_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19431_ _21021_/A _21738_/B _25610_/Q vssd1 vssd1 vccd1 vccd1 _21025_/C sky130_fd_sc_hd__nand3_1
X_16643_ _16647_/B _16643_/B vssd1 vssd1 vccd1 vccd1 _16644_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13855_ hold681/X _13854_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold682/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ hold977/X _14264_/A vssd1 vssd1 vccd1 vccd1 _12806_/X sky130_fd_sc_hd__or2_1
X_19362_ _19378_/B _19449_/B vssd1 vssd1 vccd1 vccd1 _19364_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16574_ _16574_/A _16574_/B vssd1 vssd1 vccd1 vccd1 _16596_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_130_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13786_ _13880_/A hold521/X vssd1 vssd1 vccd1 vccd1 hold522/A sky130_fd_sc_hd__nand2_1
XFILLER_0_128_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18313_ _18535_/A _18313_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _18313_/X sky130_fd_sc_hd__and3_1
XFILLER_0_85_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15525_ _22928_/B _16369_/B vssd1 vssd1 vccd1 vccd1 _16475_/B sky130_fd_sc_hd__nand2_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _14266_/A _17008_/B _14267_/B _17008_/A vssd1 vssd1 vccd1 vccd1 _12737_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19293_ _19294_/B _19294_/A vssd1 vssd1 vccd1 vccd1 _19293_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18244_ _18244_/A _18244_/B _18244_/C vssd1 vssd1 vccd1 vccd1 _21740_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_72_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15456_ _15621_/A _16424_/B vssd1 vssd1 vccd1 vccd1 _15458_/A sky130_fd_sc_hd__or2_1
X_12668_ _12668_/A vssd1 vssd1 vccd1 vccd1 _24985_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14407_ _14403_/Y hold330/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold331/A sky130_fd_sc_hd__a21oi_1
X_18175_ _18175_/A _20935_/A vssd1 vssd1 vccd1 vccd1 _18534_/A sky130_fd_sc_hd__xor2_4
X_15387_ _16817_/A _15387_/B vssd1 vssd1 vccd1 vccd1 _15388_/B sky130_fd_sc_hd__and2_1
XFILLER_0_163_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12599_ _12599_/A vssd1 vssd1 vccd1 vccd1 _12644_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_26_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17126_ _17124_/Y _17125_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _25589_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14338_ _14344_/A hold323/X vssd1 vssd1 vccd1 vccd1 hold324/A sky130_fd_sc_hd__nand2_1
Xhold506 hold506/A vssd1 vssd1 vccd1 vccd1 hold506/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold517 hold517/A vssd1 vssd1 vccd1 vccd1 hold517/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 hold528/A vssd1 vssd1 vccd1 vccd1 hold528/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold539 hold539/A vssd1 vssd1 vccd1 vccd1 hold539/X sky130_fd_sc_hd__dlygate4sd3_1
X_17057_ _20200_/B _25882_/Q _25818_/Q vssd1 vssd1 vccd1 vccd1 _17058_/B sky130_fd_sc_hd__mux2_2
X_14269_ _15839_/B vssd1 vssd1 vccd1 vccd1 _14270_/A sky130_fd_sc_hd__buf_8
X_16008_ _16212_/A hold798/X vssd1 vssd1 vccd1 vccd1 _16008_/Y sky130_fd_sc_hd__nand2_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 _13151_/X vssd1 vssd1 vccd1 vccd1 _25078_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 _25074_/Q vssd1 vssd1 vccd1 vccd1 _18178_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17959_ _20786_/B _21766_/A vssd1 vssd1 vccd1 vccd1 _20779_/A sky130_fd_sc_hd__nand2_4
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 _25062_/Q vssd1 vssd1 vccd1 vccd1 _17632_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 _19397_/Y vssd1 vssd1 vccd1 vccd1 _25729_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20970_ _20973_/A _20973_/C vssd1 vssd1 vccd1 vccd1 _20972_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_174_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19629_ _19626_/Y _19629_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19629_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_73_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22640_ _25834_/Q _22640_/B vssd1 vssd1 vccd1 vccd1 _22640_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22571_ _23088_/B vssd1 vssd1 vccd1 vccd1 _23087_/B sky130_fd_sc_hd__inv_2
XFILLER_0_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_60_clk _25472_/CLK vssd1 vssd1 vccd1 vccd1 _25539_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24310_ _24310_/A vssd1 vssd1 vccd1 vccd1 _26168_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21522_ _21636_/A _21522_/B _21521_/X vssd1 vssd1 vccd1 vccd1 _21523_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_180_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25290_ _26240_/CLK hold109/X vssd1 vssd1 vccd1 vccd1 hold107/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24241_ _24241_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24242_/A sky130_fd_sc_hd__and2_1
XFILLER_0_1_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21453_ _21453_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21458_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20404_ _25887_/Q vssd1 vssd1 vccd1 vccd1 _22375_/B sky130_fd_sc_hd__inv_2
XFILLER_0_32_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24172_ hold2340/X _26124_/Q _24203_/S vssd1 vssd1 vccd1 vccd1 _24172_/X sky130_fd_sc_hd__mux2_1
X_21384_ _21384_/A _21384_/B _21384_/C vssd1 vssd1 vccd1 vccd1 _21388_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_98_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23123_ _23123_/A _23187_/B vssd1 vssd1 vccd1 vccd1 _23123_/Y sky130_fd_sc_hd__nand2_1
X_20335_ _20335_/A _20335_/B _21086_/C vssd1 vssd1 vccd1 vccd1 _20339_/A sky130_fd_sc_hd__nand3_1
X_23054_ _23052_/X _23053_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _25892_/D sky130_fd_sc_hd__a21oi_1
X_20266_ _20265_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20266_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_179_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22005_ _22005_/A _25865_/Q vssd1 vssd1 vccd1 vccd1 _22005_/Y sky130_fd_sc_hd__nand2_1
X_20197_ _20660_/A _20197_/B vssd1 vssd1 vccd1 vccd1 _20197_/Y sky130_fd_sc_hd__nand2_1
Xhold2430 _26070_/Q vssd1 vssd1 vccd1 vccd1 hold2430/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2441 _12680_/Y vssd1 vssd1 vccd1 vccd1 _12682_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2452 _25431_/Q vssd1 vssd1 vccd1 vccd1 _15058_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2463 _25677_/Q vssd1 vssd1 vccd1 vccd1 _13265_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2474 _15576_/Y vssd1 vssd1 vccd1 vccd1 _25461_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1740 _25865_/Q vssd1 vssd1 vccd1 vccd1 _22536_/B sky130_fd_sc_hd__clkbuf_2
Xhold2485 _26287_/Q vssd1 vssd1 vccd1 vccd1 hold2485/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1751 _14962_/Y vssd1 vssd1 vccd1 vccd1 _14963_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2496 _24683_/X vssd1 vssd1 vccd1 vccd1 _24684_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23956_ hold1799/X _26054_/Q _24001_/S vssd1 vssd1 vccd1 vccd1 _23956_/X sky130_fd_sc_hd__mux2_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1762 _21758_/Y vssd1 vssd1 vccd1 vccd1 _25838_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1773 _25882_/Q vssd1 vssd1 vccd1 vccd1 _22888_/B sky130_fd_sc_hd__buf_1
XFILLER_0_99_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1784 _25620_/Q vssd1 vssd1 vccd1 vccd1 _17475_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1795 _22921_/Y vssd1 vssd1 vccd1 vccd1 _25884_/D sky130_fd_sc_hd__dlygate4sd3_1
X_22907_ _23058_/A _22907_/B vssd1 vssd1 vccd1 vccd1 _22908_/B sky130_fd_sc_hd__nand2_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23887_ _23887_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23888_/A sky130_fd_sc_hd__and2_1
X_25626_ _26135_/CLK _25626_/D vssd1 vssd1 vccd1 vccd1 _25626_/Q sky130_fd_sc_hd__dfxtp_4
X_13640_ _13703_/A _13640_/B vssd1 vssd1 vccd1 vccd1 _13640_/Y sky130_fd_sc_hd__nand2_1
X_22838_ _22937_/A _22838_/B vssd1 vssd1 vccd1 vccd1 _22838_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_184_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25557_ _25878_/CLK _25557_/D vssd1 vssd1 vccd1 vccd1 _25557_/Q sky130_fd_sc_hd__dfxtp_1
X_13571_ _13583_/A _13571_/B vssd1 vssd1 vccd1 vccd1 _13571_/Y sky130_fd_sc_hd__nand2_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22769_ _16806_/B _22421_/X _22763_/X _22764_/Y _22768_/X vssd1 vssd1 vccd1 vccd1
+ _22770_/A sky130_fd_sc_hd__a221o_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _25533_/CLK sky130_fd_sc_hd__clkbuf_16
X_15310_ _15326_/B _15311_/A vssd1 vssd1 vccd1 vccd1 _15310_/X sky130_fd_sc_hd__or2_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _12522_/A vssd1 vssd1 vccd1 vccd1 _15839_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24508_ _24508_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24509_/A sky130_fd_sc_hd__and2_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _16473_/A hold701/X vssd1 vssd1 vccd1 vccd1 hold702/A sky130_fd_sc_hd__nand2_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25488_ _25933_/CLK hold799/X vssd1 vssd1 vccd1 vccd1 hold798/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15241_ _15241_/A _15774_/B vssd1 vssd1 vccd1 vccd1 _15242_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_81_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24439_ _24439_/A vssd1 vssd1 vccd1 vccd1 _26210_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15172_ _15172_/A _15812_/B vssd1 vssd1 vccd1 vccd1 _15173_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_111_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26109_ _26109_/CLK _26109_/D vssd1 vssd1 vccd1 vccd1 _26109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14123_ _14180_/A _14123_/B vssd1 vssd1 vccd1 vccd1 _14123_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_162_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19980_ _19980_/A _19980_/B _19980_/C vssd1 vssd1 vccd1 vccd1 _19980_/X sky130_fd_sc_hd__and3_1
XFILLER_0_10_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18931_ _18951_/A _18935_/B vssd1 vssd1 vccd1 vccd1 _18933_/A sky130_fd_sc_hd__nand2_1
X_14054_ _26306_/Q _13988_/X _13981_/X _14053_/Y vssd1 vssd1 vccd1 vccd1 _14055_/B
+ sky130_fd_sc_hd__a22o_1
X_13005_ _23377_/B vssd1 vssd1 vccd1 vccd1 _13005_/X sky130_fd_sc_hd__clkbuf_8
X_18862_ _18986_/A _19616_/A vssd1 vssd1 vccd1 vccd1 _18862_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17813_ _18529_/A _17813_/B _18529_/C vssd1 vssd1 vccd1 vccd1 _17814_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_59_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18793_ _18793_/A _18793_/B _18894_/C vssd1 vssd1 vccd1 vccd1 _18794_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_59_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17744_ _17773_/B vssd1 vssd1 vccd1 vccd1 _17830_/A sky130_fd_sc_hd__inv_2
X_14956_ _14956_/A _14956_/B vssd1 vssd1 vccd1 vccd1 _14964_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_178_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13907_ _25780_/Q vssd1 vssd1 vccd1 vccd1 _18073_/B sky130_fd_sc_hd__inv_2
X_17675_ _17719_/B _23208_/B vssd1 vssd1 vccd1 vccd1 _17692_/A sky130_fd_sc_hd__nand2_1
X_14887_ _14887_/A vssd1 vssd1 vccd1 vccd1 _15076_/A sky130_fd_sc_hd__inv_2
XFILLER_0_58_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19414_ _19413_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19415_/B
+ sky130_fd_sc_hd__a211o_1
X_16626_ _16627_/B _16627_/A vssd1 vssd1 vccd1 vccd1 _16642_/B sky130_fd_sc_hd__or2_1
XFILLER_0_175_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13838_ _13880_/A hold812/X vssd1 vssd1 vccd1 vccd1 hold813/A sky130_fd_sc_hd__nand2_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19345_ _19345_/A _20856_/B vssd1 vssd1 vccd1 vccd1 _19345_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_69_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16557_ _16554_/A _16554_/B _16575_/B _16556_/Y vssd1 vssd1 vccd1 vccd1 _16557_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_174_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13769_ _25758_/Q vssd1 vssd1 vccd1 vccd1 _18652_/B sky130_fd_sc_hd__inv_2
XFILLER_0_186_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_42_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _26040_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_130_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15508_ _15508_/A _15812_/B vssd1 vssd1 vccd1 vccd1 _15509_/B sky130_fd_sc_hd__nand2_1
X_19276_ _20662_/A _22278_/B _25599_/Q vssd1 vssd1 vccd1 vccd1 _20666_/C sky130_fd_sc_hd__nand3_1
X_16488_ _16491_/A _16440_/X vssd1 vssd1 vccd1 vccd1 _16489_/B sky130_fd_sc_hd__or2b_1
XFILLER_0_169_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18227_ _18434_/A _18576_/A vssd1 vssd1 vccd1 vccd1 _18228_/B sky130_fd_sc_hd__xnor2_1
X_15439_ _15439_/A vssd1 vssd1 vccd1 vccd1 _15441_/A sky130_fd_sc_hd__inv_2
XFILLER_0_182_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18158_ _18158_/A _18158_/B vssd1 vssd1 vccd1 vccd1 _18160_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold303 hold303/A vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17109_ _17393_/A _17109_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17109_/X sky130_fd_sc_hd__and3_1
XFILLER_0_40_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold314 hold314/A vssd1 vssd1 vccd1 vccd1 hold314/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 hold325/A vssd1 vssd1 vccd1 vccd1 hold325/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18089_ _18089_/A _20624_/A vssd1 vssd1 vccd1 vccd1 _19080_/A sky130_fd_sc_hd__xor2_4
Xhold336 hold336/A vssd1 vssd1 vccd1 vccd1 hold336/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold347 hold347/A vssd1 vssd1 vccd1 vccd1 hold347/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold358 hold358/A vssd1 vssd1 vccd1 vccd1 hold358/X sky130_fd_sc_hd__dlygate4sd3_1
X_20120_ _20120_/A _21007_/C _20120_/C vssd1 vssd1 vccd1 vccd1 _20121_/B sky130_fd_sc_hd__nand3_1
Xclkbuf_4_3__f_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_3__f_clk/X
+ sky130_fd_sc_hd__clkbuf_16
Xhold369 hold369/A vssd1 vssd1 vccd1 vccd1 hold369/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20051_ _20050_/B _20051_/B _20051_/C vssd1 vssd1 vccd1 vccd1 _20052_/B sky130_fd_sc_hd__nand3b_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1003 _25069_/Q vssd1 vssd1 vccd1 vccd1 _17963_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1014 _13425_/X vssd1 vssd1 vccd1 vccd1 _25122_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1025 _25037_/Q vssd1 vssd1 vccd1 vccd1 _17449_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 _13124_/X vssd1 vssd1 vccd1 vccd1 _25073_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23810_ _23810_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23811_/A sky130_fd_sc_hd__and2_1
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1047 _25748_/Q vssd1 vssd1 vccd1 vccd1 _19667_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 _12787_/X vssd1 vssd1 vccd1 vccd1 _25009_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24790_ hold1918/X _26325_/Q _24817_/S vssd1 vssd1 vccd1 vccd1 _24790_/X sky130_fd_sc_hd__mux2_1
Xhold1069 _25044_/Q vssd1 vssd1 vccd1 vccd1 _17500_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23741_ _23741_/A vssd1 vssd1 vccd1 vccd1 _25985_/D sky130_fd_sc_hd__clkbuf_1
X_20953_ _20953_/A _20953_/B vssd1 vssd1 vccd1 vccd1 _20954_/A sky130_fd_sc_hd__nand2_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23672_ _23672_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23673_/A sky130_fd_sc_hd__and2_1
X_20884_ _20886_/A _20886_/C vssd1 vssd1 vccd1 vccd1 _20885_/A sky130_fd_sc_hd__nand2_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25411_ _26004_/CLK _25411_/D vssd1 vssd1 vccd1 vccd1 _25411_/Q sky130_fd_sc_hd__dfxtp_1
X_22623_ _23119_/B _22975_/B vssd1 vssd1 vccd1 vccd1 _22625_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_33_clk _25184_/CLK vssd1 vssd1 vccd1 vccd1 _25895_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22554_ _26049_/Q vssd1 vssd1 vccd1 vccd1 _22555_/A sky130_fd_sc_hd__inv_2
X_25342_ _26298_/CLK hold130/X vssd1 vssd1 vccd1 vccd1 hold128/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21505_ _21504_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21505_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22485_ _22561_/A _22485_/B vssd1 vssd1 vccd1 vccd1 _22485_/Y sky130_fd_sc_hd__nand2_1
X_25273_ _26231_/CLK hold334/X vssd1 vssd1 vccd1 vccd1 hold332/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24224_ _24224_/A vssd1 vssd1 vccd1 vccd1 _26140_/D sky130_fd_sc_hd__clkbuf_1
X_21436_ _21436_/A _21436_/B vssd1 vssd1 vccd1 vccd1 _21437_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_133_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24155_ _24155_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24156_/A sky130_fd_sc_hd__and2_1
X_21367_ _21417_/A _21370_/A vssd1 vssd1 vccd1 vccd1 _21368_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23106_ _23106_/A _23106_/B vssd1 vssd1 vccd1 vccd1 _23107_/A sky130_fd_sc_hd__xor2_1
X_20318_ _20318_/A _20318_/B _20318_/C vssd1 vssd1 vccd1 vccd1 _20319_/B sky130_fd_sc_hd__nand3_1
X_24086_ hold2185/X hold1832/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24087_/A sky130_fd_sc_hd__mux2_1
Xhold870 hold870/A vssd1 vssd1 vccd1 vccd1 hold870/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21298_ _21298_/A _21298_/B vssd1 vssd1 vccd1 vccd1 _21707_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_130_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold881 hold881/A vssd1 vssd1 vccd1 vccd1 hold881/X sky130_fd_sc_hd__dlygate4sd3_1
X_23037_ _23197_/A _23037_/B vssd1 vssd1 vccd1 vccd1 _23037_/Y sky130_fd_sc_hd__nand2_1
Xhold892 hold892/A vssd1 vssd1 vccd1 vccd1 hold892/X sky130_fd_sc_hd__dlygate4sd3_1
X_20249_ _20251_/A _20251_/C vssd1 vssd1 vccd1 vccd1 _20250_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2260 _24979_/Q vssd1 vssd1 vccd1 vccd1 _12629_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ _25850_/Q _12527_/A _14996_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14810_/X
+ sky130_fd_sc_hd__a22o_1
Xhold2271 _24972_/Q vssd1 vssd1 vccd1 vccd1 _12594_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2282 _24154_/X vssd1 vssd1 vccd1 vccd1 _24155_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2293 _26054_/Q vssd1 vssd1 vccd1 vccd1 hold2293/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _16977_/B vssd1 vssd1 vccd1 vccd1 _23175_/B sky130_fd_sc_hd__inv_2
X_24988_ _24990_/CLK _24988_/D vssd1 vssd1 vccd1 vccd1 _24988_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1570 _25812_/Q vssd1 vssd1 vccd1 vccd1 _21315_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14741_ _15464_/A vssd1 vssd1 vccd1 vccd1 _14741_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_93_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1581 _19998_/Y vssd1 vssd1 vccd1 vccd1 _25773_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23939_ _23939_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23940_/A sky130_fd_sc_hd__and2_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1592 _25781_/Q vssd1 vssd1 vccd1 vccd1 _20307_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17460_ _17467_/A _17460_/B vssd1 vssd1 vccd1 vccd1 _17460_/Y sky130_fd_sc_hd__nand2_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _14672_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _14672_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16411_ _16676_/A _16411_/B vssd1 vssd1 vccd1 vccd1 _16413_/A sky130_fd_sc_hd__or2_1
XFILLER_0_157_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_3_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_25609_ _26116_/CLK _25609_/D vssd1 vssd1 vccd1 vccd1 _25609_/Q sky130_fd_sc_hd__dfxtp_2
X_13623_ hold492/X _13622_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold493/A sky130_fd_sc_hd__a21oi_1
X_17391_ _17571_/A _17622_/B vssd1 vssd1 vccd1 vccd1 _17392_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_clk _25759_/CLK vssd1 vssd1 vccd1 vccd1 _25174_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_172_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19130_ _21228_/A vssd1 vssd1 vccd1 vccd1 _19130_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16342_ _16473_/A hold906/X vssd1 vssd1 vccd1 vccd1 _16342_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_39_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13554_ _13642_/A hold446/X vssd1 vssd1 vccd1 vccd1 hold447/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12505_ _23597_/A vssd1 vssd1 vccd1 vccd1 _12560_/A sky130_fd_sc_hd__inv_2
XFILLER_0_124_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19061_ _19082_/A _19061_/B _22786_/A vssd1 vssd1 vccd1 vccd1 _19061_/X sky130_fd_sc_hd__and3_1
X_16273_ _16273_/A _16273_/B _16273_/C vssd1 vssd1 vccd1 vccd1 _16274_/B sky130_fd_sc_hd__and3_1
X_13485_ hold716/X _13484_/Y _12558_/B vssd1 vssd1 vccd1 vccd1 hold717/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_164_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18012_ _18010_/Y _18011_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _25650_/D sky130_fd_sc_hd__a21oi_1
X_15224_ _15224_/A _15774_/B vssd1 vssd1 vccd1 vccd1 _15225_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_22_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15155_ _22501_/B _16369_/B vssd1 vssd1 vccd1 vccd1 _15156_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_23_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14106_ _14118_/A hold527/X vssd1 vssd1 vccd1 vccd1 hold528/A sky130_fd_sc_hd__nand2_1
X_15086_ _15066_/B _15085_/B _15077_/B vssd1 vssd1 vccd1 vccd1 _15086_/X sky130_fd_sc_hd__o21a_1
X_19963_ _19958_/X _19962_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19963_/Y sky130_fd_sc_hd__o21ai_1
X_14037_ _14345_/A vssd1 vssd1 vccd1 vccd1 _14037_/X sky130_fd_sc_hd__clkbuf_8
X_18914_ _18955_/A _18914_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18915_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_129_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19894_ _19893_/Y _19130_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19896_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18845_ _25704_/Q vssd1 vssd1 vccd1 vccd1 _22590_/B sky130_fd_sc_hd__inv_2
XFILLER_0_101_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18776_ _18776_/A _20596_/A vssd1 vssd1 vccd1 vccd1 _19017_/B sky130_fd_sc_hd__xor2_4
X_15988_ _15999_/B _15989_/A vssd1 vssd1 vccd1 vccd1 _15988_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17727_ _17727_/A vssd1 vssd1 vccd1 vccd1 _17728_/C sky130_fd_sc_hd__inv_2
X_14939_ _14939_/A _14939_/B vssd1 vssd1 vccd1 vccd1 _14947_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_4_11__f_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_11__f_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17658_ _20023_/B _21749_/A vssd1 vssd1 vccd1 vccd1 _17662_/A sky130_fd_sc_hd__nand2_1
X_16609_ _16629_/B _16629_/C vssd1 vssd1 vccd1 vccd1 _16610_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_169_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17589_ _21791_/A vssd1 vssd1 vccd1 vccd1 _18180_/B sky130_fd_sc_hd__buf_6
XFILLER_0_58_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_clk _25184_/CLK vssd1 vssd1 vccd1 vccd1 _26279_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19328_ _26228_/Q hold560/X vssd1 vssd1 vccd1 vccd1 _19328_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_46_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19259_ _20624_/A _19257_/Y _20628_/C vssd1 vssd1 vccd1 vccd1 _19350_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22270_ _19673_/A _22269_/A _22269_/Y vssd1 vssd1 vccd1 vccd1 _22272_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_170_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold100 hold100/A vssd1 vssd1 vccd1 vccd1 hold100/X sky130_fd_sc_hd__dlygate4sd3_1
X_21221_ _21613_/B _21659_/C vssd1 vssd1 vccd1 vccd1 _21222_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold111 hold111/A vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 hold122/A vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 hold133/A vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 hold144/A vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__dlygate4sd3_1
X_21152_ _23199_/A vssd1 vssd1 vccd1 vccd1 _21508_/B sky130_fd_sc_hd__buf_6
XFILLER_0_112_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold155 hold155/A vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 hold166/A vssd1 vssd1 vccd1 vccd1 hold166/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold177 hold177/A vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 hold188/A vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
X_20103_ _20106_/A _20106_/B vssd1 vssd1 vccd1 vccd1 _20105_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_186_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold199 hold199/A vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
X_25960_ _26073_/CLK _25960_/D vssd1 vssd1 vccd1 vccd1 _25960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21083_ _21580_/B vssd1 vssd1 vccd1 vccd1 _21577_/C sky130_fd_sc_hd__inv_2
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24911_ hold866/A hold935/A _24942_/S vssd1 vssd1 vccd1 vccd1 _24912_/B sky130_fd_sc_hd__mux2_1
X_20034_ _20034_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20039_/A sky130_fd_sc_hd__nand2_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25891_ _25893_/CLK _25891_/D vssd1 vssd1 vccd1 vccd1 _25891_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24842_ _15231_/A _15247_/B _24860_/S vssd1 vssd1 vccd1 vccd1 _24842_/X sky130_fd_sc_hd__mux2_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24773_ _24773_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24774_/A sky130_fd_sc_hd__and2_1
X_21985_ _22740_/B _21986_/A vssd1 vssd1 vccd1 vccd1 _21987_/A sky130_fd_sc_hd__or2_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23724_ _24560_/A vssd1 vssd1 vccd1 vccd1 _23813_/B sky130_fd_sc_hd__buf_8
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ _20936_/A _20936_/B vssd1 vssd1 vccd1 vccd1 _20940_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23655_ _23655_/A vssd1 vssd1 vccd1 vccd1 _25957_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20867_ _21676_/A _21451_/B vssd1 vssd1 vccd1 vccd1 _20868_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_187_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22606_ _22606_/A _22606_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22608_/A sky130_fd_sc_hd__or3_1
XFILLER_0_113_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23586_ _23586_/A _23586_/B vssd1 vssd1 vccd1 vccd1 _23587_/C sky130_fd_sc_hd__or2_1
X_20798_ _20797_/B _20798_/B _20798_/C vssd1 vssd1 vccd1 vccd1 _20799_/B sky130_fd_sc_hd__nand3b_2
XFILLER_0_165_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25325_ _25712_/CLK hold298/X vssd1 vssd1 vccd1 vccd1 hold296/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22537_ _22535_/X _22536_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22537_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25256_ _25257_/CLK hold433/X vssd1 vssd1 vccd1 vccd1 hold431/A sky130_fd_sc_hd__dfxtp_1
X_13270_ _13207_/X _13268_/X _13192_/X _13269_/X vssd1 vssd1 vccd1 vccd1 _13270_/X
+ sky130_fd_sc_hd__o211a_1
X_22468_ _22468_/A _22468_/B vssd1 vssd1 vccd1 vccd1 _22469_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24207_ hold2391/X hold2280/X _24279_/S vssd1 vssd1 vccd1 vccd1 _24208_/A sky130_fd_sc_hd__mux2_1
X_21419_ _21419_/A _21419_/B _21419_/C vssd1 vssd1 vccd1 vccd1 _21420_/B sky130_fd_sc_hd__nand3_1
X_22399_ _22824_/A _22974_/B vssd1 vssd1 vccd1 vccd1 _22402_/A sky130_fd_sc_hd__nand2_1
X_25187_ _25770_/CLK hold661/X vssd1 vssd1 vccd1 vccd1 hold659/A sky130_fd_sc_hd__dfxtp_1
X_24138_ _24138_/A vssd1 vssd1 vccd1 vccd1 _26112_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16960_ _16960_/A _16960_/B vssd1 vssd1 vccd1 vccd1 _16960_/Y sky130_fd_sc_hd__nand2_1
X_24069_ _24069_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24070_/A sky130_fd_sc_hd__and2_1
XFILLER_0_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15911_ _15911_/A _15921_/A vssd1 vssd1 vccd1 vccd1 _15911_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_159_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16891_ _16889_/X _16711_/X _16890_/Y _25888_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16892_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_95_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18630_ _18630_/A _25821_/Q _18630_/C vssd1 vssd1 vccd1 vccd1 _20330_/B sky130_fd_sc_hd__nand3_2
X_15842_ _21721_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _15844_/A sky130_fd_sc_hd__nand2_1
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2090 _26190_/Q vssd1 vssd1 vccd1 vccd1 hold2090/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18561_ _18559_/Y _18560_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25672_/D sky130_fd_sc_hd__a21oi_1
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _26042_/Q _25978_/Q _15773_/S vssd1 vssd1 vccd1 vccd1 _15774_/A sky130_fd_sc_hd__mux2_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12985_ _25047_/Q _13133_/B vssd1 vssd1 vccd1 vccd1 _12985_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17512_ _17512_/A _17562_/A vssd1 vssd1 vccd1 vccd1 _17513_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14724_ _14731_/B _21831_/A vssd1 vssd1 vccd1 vccd1 _21830_/B sky130_fd_sc_hd__xnor2_2
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18492_ _18492_/A _20054_/A vssd1 vssd1 vccd1 vccd1 _18838_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_157_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17443_ _17441_/X _17241_/X _17442_/X vssd1 vssd1 vccd1 vccd1 _17444_/A sky130_fd_sc_hd__a21o_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14655_ _14688_/A hold167/X vssd1 vssd1 vccd1 vccd1 hold168/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ _25732_/Q vssd1 vssd1 vccd1 vccd1 _18052_/B sky130_fd_sc_hd__inv_2
XFILLER_0_185_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17374_ _17372_/X _17241_/X _17373_/X vssd1 vssd1 vccd1 vccd1 _17375_/A sky130_fd_sc_hd__a21o_1
X_14586_ _15464_/A vssd1 vssd1 vccd1 vccd1 _14586_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19113_ _19111_/Y _19112_/Y _19086_/X vssd1 vssd1 vccd1 vccd1 _19113_/Y sky130_fd_sc_hd__a21oi_1
X_16325_ _16323_/X _16324_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _16325_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_184_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13537_ _25721_/Q vssd1 vssd1 vccd1 vccd1 _17858_/B sky130_fd_sc_hd__inv_2
XFILLER_0_171_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19044_ _19042_/Y _19043_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25703_/D sky130_fd_sc_hd__a21oi_1
X_16256_ _16252_/B _16252_/A _16269_/B _16255_/Y vssd1 vssd1 vccd1 vccd1 _16256_/X
+ sky130_fd_sc_hd__a31o_1
X_13468_ _14170_/A vssd1 vssd1 vccd1 vccd1 _13468_/X sky130_fd_sc_hd__buf_12
XFILLER_0_113_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15207_ _15207_/A _15776_/B vssd1 vssd1 vccd1 vccd1 _15208_/B sky130_fd_sc_hd__nand2_2
X_16187_ _16185_/X _16186_/Y _16076_/X vssd1 vssd1 vccd1 vccd1 _25501_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13399_ _19005_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13399_/X sky130_fd_sc_hd__or2_1
XFILLER_0_51_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15138_ _22479_/B _15138_/B vssd1 vssd1 vccd1 vccd1 _22476_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_26_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15069_ _15069_/A vssd1 vssd1 vccd1 vccd1 _15108_/A sky130_fd_sc_hd__inv_2
X_19946_ _26272_/Q _19134_/X hold812/X vssd1 vssd1 vccd1 vccd1 _19947_/C sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_4_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _25716_/CLK sky130_fd_sc_hd__clkbuf_16
X_19877_ _19870_/X _19876_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19877_/Y sky130_fd_sc_hd__o21ai_1
X_18828_ _25895_/Q _22563_/A vssd1 vssd1 vccd1 vccd1 _18836_/A sky130_fd_sc_hd__or2_2
XFILLER_0_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18759_ _19026_/A _18759_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18759_/X sky130_fd_sc_hd__and3_1
X_21770_ _21770_/A _21770_/B vssd1 vssd1 vccd1 vccd1 _23072_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_72_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20721_ _20721_/A _20721_/B vssd1 vssd1 vccd1 vccd1 _21661_/B sky130_fd_sc_hd__nand2_8
XFILLER_0_187_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23440_ hold329/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23440_/X sky130_fd_sc_hd__or2b_1
X_20652_ _20652_/A _20652_/B vssd1 vssd1 vccd1 vccd1 _20653_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23371_ _23376_/A vssd1 vssd1 vccd1 vccd1 _23373_/A sky130_fd_sc_hd__inv_2
XFILLER_0_116_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20583_ _20660_/A _20583_/B vssd1 vssd1 vccd1 vccd1 _20583_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25110_ _26193_/CLK _25110_/D vssd1 vssd1 vccd1 vccd1 _25110_/Q sky130_fd_sc_hd__dfxtp_1
X_22322_ _22653_/A _22322_/B vssd1 vssd1 vccd1 vccd1 _22322_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26090_ _26221_/CLK _26090_/D vssd1 vssd1 vccd1 vccd1 hold992/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22253_ _22253_/A _25854_/Q vssd1 vssd1 vccd1 vccd1 _22254_/B sky130_fd_sc_hd__nand2_1
X_25041_ _26216_/CLK _25041_/D vssd1 vssd1 vccd1 vccd1 _25041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21204_ _21202_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21204_/X
+ sky130_fd_sc_hd__a211o_1
X_22184_ _22184_/A _22855_/B vssd1 vssd1 vccd1 vccd1 _22185_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21135_ _21135_/A _21135_/B vssd1 vssd1 vccd1 vccd1 _21137_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25943_ _26073_/CLK _25943_/D vssd1 vssd1 vccd1 vccd1 _25943_/Q sky130_fd_sc_hd__dfxtp_1
X_21066_ _26306_/Q _20731_/X hold512/X vssd1 vssd1 vccd1 vccd1 _21069_/B sky130_fd_sc_hd__a21oi_1
X_20017_ _20017_/A _20017_/B vssd1 vssd1 vccd1 vccd1 _20019_/A sky130_fd_sc_hd__nand2_1
X_25874_ _25877_/CLK _25874_/D vssd1 vssd1 vccd1 vccd1 _25874_/Q sky130_fd_sc_hd__dfxtp_2
X_24825_ _24825_/A vssd1 vssd1 vccd1 vccd1 _26336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _26089_/Q _12748_/X _12769_/X vssd1 vssd1 vccd1 vccd1 _12770_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_16_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24756_ _24756_/A vssd1 vssd1 vccd1 vccd1 _26313_/D sky130_fd_sc_hd__clkbuf_1
X_21968_ _21968_/A _22145_/B vssd1 vssd1 vccd1 vccd1 _21968_/Y sky130_fd_sc_hd__nand2_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23707_ _23707_/A vssd1 vssd1 vccd1 vccd1 _25974_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20919_ _21480_/C _21709_/A vssd1 vssd1 vccd1 vccd1 _20921_/A sky130_fd_sc_hd__nand2_1
X_24687_ _24687_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24688_/A sky130_fd_sc_hd__and2_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21899_ _22653_/A _21899_/B vssd1 vssd1 vccd1 vccd1 _21899_/X sky130_fd_sc_hd__or2_1
XFILLER_0_83_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _14440_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14440_/Y sky130_fd_sc_hd__nand2_1
X_23638_ hold2094/X _25952_/Q _23677_/S vssd1 vssd1 vccd1 vccd1 _23638_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_37_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14371_ _14404_/A hold218/X vssd1 vssd1 vccd1 vccd1 hold219/A sky130_fd_sc_hd__nand2_1
XFILLER_0_107_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23569_ hold230/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23569_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_37_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16110_ hold428/X vssd1 vssd1 vccd1 vccd1 _16113_/B sky130_fd_sc_hd__inv_2
XFILLER_0_135_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25308_ _26135_/CLK hold124/X vssd1 vssd1 vccd1 vccd1 hold122/A sky130_fd_sc_hd__dfxtp_1
X_13322_ _13322_/A vssd1 vssd1 vccd1 vccd1 _19602_/A sky130_fd_sc_hd__buf_4
XFILLER_0_88_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17090_ _19687_/A _17090_/B vssd1 vssd1 vccd1 vccd1 _17526_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_165_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26288_ _26289_/CLK _26288_/D vssd1 vssd1 vccd1 vccd1 _26288_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_52_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16041_ _16052_/B _16042_/A vssd1 vssd1 vccd1 vccd1 _16041_/X sky130_fd_sc_hd__or2_1
X_13253_ _13253_/A vssd1 vssd1 vccd1 vccd1 _19444_/A sky130_fd_sc_hd__buf_4
X_25239_ _25817_/CLK hold826/X vssd1 vssd1 vccd1 vccd1 hold825/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13184_ _13049_/X _14548_/A _13067_/X _19289_/A vssd1 vssd1 vccd1 vccd1 _13184_/X
+ sky130_fd_sc_hd__a22o_1
X_19800_ _19799_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19801_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17992_ _17992_/A _20546_/A vssd1 vssd1 vccd1 vccd1 _19066_/A sky130_fd_sc_hd__xor2_4
X_16943_ _22680_/A vssd1 vssd1 vccd1 vccd1 _22145_/B sky130_fd_sc_hd__buf_8
X_19731_ _20400_/A _19729_/Y _20405_/C vssd1 vssd1 vccd1 vccd1 _19821_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16874_ _16935_/A _16879_/B vssd1 vssd1 vccd1 vccd1 _16876_/B sky130_fd_sc_hd__nand2_1
X_19662_ _19678_/B _19749_/B vssd1 vssd1 vccd1 vccd1 _19664_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15825_ _15825_/A _15829_/B vssd1 vssd1 vccd1 vccd1 _15828_/A sky130_fd_sc_hd__nand2_1
X_18613_ _18613_/A _18613_/B _18613_/C vssd1 vssd1 vccd1 vccd1 _22299_/A sky130_fd_sc_hd__nand3_1
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19593_ _19593_/A _19593_/B vssd1 vssd1 vccd1 vccd1 _19593_/Y sky130_fd_sc_hd__nand2_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15756_ _23143_/B _15756_/B vssd1 vssd1 vccd1 vccd1 _23140_/B sky130_fd_sc_hd__xor2_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18544_ _18544_/A _18544_/B vssd1 vssd1 vccd1 vccd1 _22207_/A sky130_fd_sc_hd__nand2_1
X_12968_ _26127_/Q _12907_/X _12967_/X vssd1 vssd1 vccd1 vccd1 _12968_/X sky130_fd_sc_hd__a21o_1
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14707_ _21759_/B _15543_/B vssd1 vssd1 vccd1 vccd1 _14907_/B sky130_fd_sc_hd__nand2_1
X_18475_ _18535_/A _18475_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18475_/X sky130_fd_sc_hd__and3_1
X_15687_ _16605_/A _15778_/B vssd1 vssd1 vccd1 vccd1 _16930_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_157_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _26114_/Q _12748_/X _12898_/X vssd1 vssd1 vccd1 vccd1 _12899_/X sky130_fd_sc_hd__a21o_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17426_ _17426_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17426_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14638_ _14638_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14638_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_185_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17357_ _17355_/Y _17356_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _25607_/D sky130_fd_sc_hd__a21oi_1
X_14569_ _14569_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14569_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_56_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16308_ _16333_/A vssd1 vssd1 vccd1 vccd1 _16313_/B sky130_fd_sc_hd__inv_2
X_17288_ _25609_/Q vssd1 vssd1 vccd1 vccd1 _20994_/B sky130_fd_sc_hd__inv_2
XFILLER_0_70_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19027_ _19025_/X _18879_/X _19026_/X vssd1 vssd1 vccd1 vccd1 _19028_/A sky130_fd_sc_hd__a21o_1
X_16239_ _16245_/A _16240_/A vssd1 vssd1 vccd1 vccd1 _16239_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19929_ _19927_/X _19928_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19929_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22940_ _22940_/A _22940_/B vssd1 vssd1 vccd1 vccd1 _22942_/A sky130_fd_sc_hd__nand2_1
X_22871_ _22862_/Y _22870_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22871_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24610_ _24610_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24611_/A sky130_fd_sc_hd__and2_1
X_21822_ _17881_/B _17048_/B _17882_/B vssd1 vssd1 vccd1 vccd1 _21823_/B sky130_fd_sc_hd__o21ai_2
X_25590_ _25594_/CLK _25590_/D vssd1 vssd1 vccd1 vccd1 _25590_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_148_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24541_ hold2696/X _26244_/Q _24587_/S vssd1 vssd1 vccd1 vccd1 _24541_/X sky130_fd_sc_hd__mux2_1
X_21753_ _21754_/A _21754_/B _22745_/A vssd1 vssd1 vccd1 vccd1 _21753_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20704_ _20704_/A _25856_/Q vssd1 vssd1 vccd1 vccd1 _20708_/B sky130_fd_sc_hd__nand2_1
X_24472_ _24472_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24473_/A sky130_fd_sc_hd__and2_1
XFILLER_0_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21684_ _21716_/A _21684_/B _21683_/X vssd1 vssd1 vccd1 vccd1 _21685_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_175_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26211_ _26339_/CLK _26211_/D vssd1 vssd1 vccd1 vccd1 _26211_/Q sky130_fd_sc_hd__dfxtp_1
X_23423_ _24940_/S hold242/A _23422_/X vssd1 vssd1 vccd1 vccd1 _23423_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_188_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20635_ _20635_/A _20635_/B vssd1 vssd1 vccd1 vccd1 _20639_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26142_ _26142_/CLK _26142_/D vssd1 vssd1 vccd1 vccd1 _26142_/Q sky130_fd_sc_hd__dfxtp_1
X_23354_ _23354_/A vssd1 vssd1 vccd1 vccd1 _23356_/B sky130_fd_sc_hd__inv_2
XFILLER_0_150_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20566_ _20566_/A _20566_/B _20566_/C vssd1 vssd1 vccd1 vccd1 _20567_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22305_ _22906_/B _22758_/B vssd1 vssd1 vccd1 vccd1 _22317_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26073_ _26073_/CLK _26073_/D vssd1 vssd1 vccd1 vccd1 _26073_/Q sky130_fd_sc_hd__dfxtp_1
X_23285_ _23293_/B _23307_/A vssd1 vssd1 vccd1 vccd1 _23287_/A sky130_fd_sc_hd__or2_1
XFILLER_0_132_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20497_ _20497_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20502_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_131_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25024_ _25604_/CLK _25024_/D vssd1 vssd1 vccd1 vccd1 _25024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22236_ _22236_/A _25882_/Q vssd1 vssd1 vccd1 vccd1 _22236_/Y sky130_fd_sc_hd__nand2_1
X_22167_ _22168_/A _22168_/C _23106_/A vssd1 vssd1 vccd1 vccd1 _22167_/X sky130_fd_sc_hd__a21o_1
X_21118_ _21118_/A _21118_/B vssd1 vssd1 vccd1 vccd1 _21119_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22098_ _19588_/A _22097_/A _22097_/Y vssd1 vssd1 vccd1 vccd1 _22100_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_22_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25926_ _25939_/CLK _25926_/D vssd1 vssd1 vccd1 vccd1 _25926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13940_ _26288_/Q _13801_/X _13793_/X _13939_/Y vssd1 vssd1 vccd1 vccd1 _13941_/B
+ sky130_fd_sc_hd__a22o_1
X_21049_ _21051_/B _21051_/C vssd1 vssd1 vccd1 vccd1 _21050_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25857_ _26339_/CLK _25857_/D vssd1 vssd1 vccd1 vccd1 _25857_/Q sky130_fd_sc_hd__dfxtp_4
X_13871_ _26277_/Q _13801_/X _13793_/X _13870_/Y vssd1 vssd1 vccd1 vccd1 _13872_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15610_ _15608_/X _15609_/Y _15464_/X vssd1 vssd1 vccd1 vccd1 _15610_/Y sky130_fd_sc_hd__a21oi_1
X_24808_ _26330_/Q hold2693/X _24817_/S vssd1 vssd1 vccd1 vccd1 _24808_/X sky130_fd_sc_hd__mux2_1
X_12822_ _17214_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12822_/X sky130_fd_sc_hd__or2_1
X_16590_ _16574_/B _16589_/Y _16574_/A vssd1 vssd1 vccd1 vccd1 _16591_/B sky130_fd_sc_hd__o21bai_1
X_25788_ _25793_/CLK _25788_/D vssd1 vssd1 vccd1 vccd1 _25788_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_9_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15541_ _22945_/B _15774_/B vssd1 vssd1 vccd1 vccd1 _15542_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12753_ _12726_/B _14292_/A _12752_/X _25583_/Q vssd1 vssd1 vccd1 vccd1 _12753_/X
+ sky130_fd_sc_hd__a22o_1
X_24739_ _24739_/A vssd1 vssd1 vccd1 vccd1 _26308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ _18446_/A _25739_/Q _21716_/A vssd1 vssd1 vccd1 vccd1 _18261_/C sky130_fd_sc_hd__nand3_1
X_15472_ _26025_/Q _25961_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15473_/A sky130_fd_sc_hd__mux2_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12684_ _12684_/A _12684_/B vssd1 vssd1 vccd1 vccd1 _12686_/A sky130_fd_sc_hd__nor2_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17211_ _19816_/A _17211_/B vssd1 vssd1 vccd1 vccd1 _17593_/A sky130_fd_sc_hd__xor2_4
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _14465_/A hold299/X vssd1 vssd1 vccd1 vccd1 hold300/A sky130_fd_sc_hd__nand2_1
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18191_ _18191_/A _20357_/A vssd1 vssd1 vccd1 vccd1 _20349_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17142_ _19257_/A _17142_/B vssd1 vssd1 vccd1 vccd1 _17478_/A sky130_fd_sc_hd__xor2_4
X_14354_ _14352_/Y hold291/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold292/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13305_ _13220_/X _14608_/A _13242_/X _19560_/A vssd1 vssd1 vccd1 vccd1 _13305_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17073_ _20236_/B _25883_/Q _25819_/Q vssd1 vssd1 vccd1 vccd1 _17074_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_12_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14285_ _14588_/A vssd1 vssd1 vccd1 vccd1 _14687_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_0_122_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16024_ _16040_/B _16024_/B vssd1 vssd1 vccd1 vccd1 _16052_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_123_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13236_ _26175_/Q _13065_/X _13235_/X vssd1 vssd1 vccd1 vccd1 _13236_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_20_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13167_ _26164_/Q _13065_/X _13166_/X vssd1 vssd1 vccd1 vccd1 _13167_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13098_ _13018_/X _13095_/X _13096_/X _13097_/X vssd1 vssd1 vccd1 vccd1 _13098_/X
+ sky130_fd_sc_hd__o211a_1
X_17975_ _17976_/B _17976_/A vssd1 vssd1 vccd1 vccd1 _20178_/A sky130_fd_sc_hd__or2_1
X_19714_ _19711_/Y _19714_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19714_/X sky130_fd_sc_hd__and3b_1
X_16926_ _16977_/A _16926_/B vssd1 vssd1 vccd1 vccd1 _16926_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_137_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19645_ _20162_/A _22208_/B _25625_/Q vssd1 vssd1 vccd1 vccd1 _20167_/C sky130_fd_sc_hd__nand3_1
X_16857_ _16857_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16857_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15808_ _15808_/A vssd1 vssd1 vccd1 vccd1 _23191_/B sky130_fd_sc_hd__inv_2
XFILLER_0_133_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16788_ _16786_/X _16711_/X _16787_/Y _25873_/Q _14170_/X vssd1 vssd1 vccd1 vccd1
+ _16789_/A sky130_fd_sc_hd__a32o_1
X_19576_ _21290_/A _19574_/Y _21294_/C vssd1 vssd1 vccd1 vccd1 _19664_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15739_ _23127_/B _15739_/B vssd1 vssd1 vccd1 vccd1 _23124_/B sky130_fd_sc_hd__xor2_1
X_18527_ _18527_/A _25816_/Q _18527_/C vssd1 vssd1 vccd1 vccd1 _20139_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_88_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18458_ _18641_/A _19331_/A vssd1 vssd1 vccd1 vccd1 _18458_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17409_ _25620_/Q vssd1 vssd1 vccd1 vccd1 _21291_/B sky130_fd_sc_hd__inv_2
XFILLER_0_173_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18389_ _21216_/B _21983_/A vssd1 vssd1 vccd1 vccd1 _21210_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_56_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20420_ _26287_/Q _20078_/X hold686/X vssd1 vssd1 vccd1 vccd1 _20423_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20351_ _20354_/A _20354_/C vssd1 vssd1 vccd1 vccd1 _20352_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_125_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23070_ _23068_/X _23069_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _23070_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20282_ _20282_/A _20282_/B vssd1 vssd1 vccd1 vccd1 _21482_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_178_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22021_ _22021_/A _22021_/B vssd1 vssd1 vccd1 vccd1 _22742_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2601 _24495_/X vssd1 vssd1 vccd1 vccd1 _24496_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2612 _26290_/Q vssd1 vssd1 vccd1 vccd1 hold2612/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2623 _15534_/X vssd1 vssd1 vccd1 vccd1 hold2623/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2634 _26271_/Q vssd1 vssd1 vccd1 vccd1 hold2634/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1900 _26014_/Q vssd1 vssd1 vccd1 vccd1 hold1900/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2645 _24760_/X vssd1 vssd1 vccd1 vccd1 _24761_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1911 _26089_/Q vssd1 vssd1 vccd1 vccd1 hold1911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2656 _24781_/X vssd1 vssd1 vccd1 vccd1 _24782_/A sky130_fd_sc_hd__dlygate4sd3_1
X_23972_ _23972_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23973_/A sky130_fd_sc_hd__and2_1
Xhold1922 output8/A vssd1 vssd1 vccd1 vccd1 _23278_/B sky130_fd_sc_hd__buf_2
Xhold2667 _26300_/Q vssd1 vssd1 vccd1 vccd1 hold2667/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1933 _23886_/X vssd1 vssd1 vccd1 vccd1 _23887_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2678 _23238_/Y vssd1 vssd1 vccd1 vccd1 hold2678/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1944 _23815_/X vssd1 vssd1 vccd1 vccd1 _23817_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2689 _26247_/Q vssd1 vssd1 vccd1 vccd1 hold2689/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25711_ _25711_/CLK hold670/X vssd1 vssd1 vccd1 vccd1 hold668/A sky130_fd_sc_hd__dfxtp_1
X_22923_ _22923_/A _22923_/B vssd1 vssd1 vccd1 vccd1 _22925_/A sky130_fd_sc_hd__nand2_1
Xhold1955 _26116_/Q vssd1 vssd1 vccd1 vccd1 hold1955/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1966 _23764_/X vssd1 vssd1 vccd1 vccd1 _23765_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1977 _23920_/X vssd1 vssd1 vccd1 vccd1 _23921_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1988 _26208_/Q vssd1 vssd1 vccd1 vccd1 hold1988/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1999 _26236_/Q vssd1 vssd1 vccd1 vccd1 hold1999/X sky130_fd_sc_hd__dlygate4sd3_1
X_25642_ _26148_/CLK _25642_/D vssd1 vssd1 vccd1 vccd1 _25642_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_168_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22854_ _22844_/Y _22853_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22854_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_79_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21805_ _21806_/B _21806_/A vssd1 vssd1 vccd1 vccd1 _21807_/A sky130_fd_sc_hd__or2_1
X_25573_ _25573_/CLK _25573_/D vssd1 vssd1 vccd1 vccd1 _25573_/Q sky130_fd_sc_hd__dfxtp_1
X_22785_ _16813_/B _22421_/X _22779_/X _22780_/Y _22784_/X vssd1 vssd1 vccd1 vccd1
+ _22787_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24524_ _24524_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24525_/A sky130_fd_sc_hd__and2_1
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21736_ _23056_/A vssd1 vssd1 vccd1 vccd1 _23055_/A sky130_fd_sc_hd__inv_2
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24455_ hold2654/X hold2592/X _24510_/S vssd1 vssd1 vccd1 vccd1 _24456_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_149_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21667_ _21666_/Y _21203_/X _20986_/A _20957_/A vssd1 vssd1 vccd1 vccd1 _21667_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23406_ _23400_/X _23405_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _23406_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20618_ _20617_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20618_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24386_ _24386_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24387_/A sky130_fd_sc_hd__and2_1
X_21598_ _21598_/A _21598_/B vssd1 vssd1 vccd1 vccd1 _21599_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_151_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26125_ _26216_/CLK _26125_/D vssd1 vssd1 vccd1 vccd1 _26125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23337_ _23342_/A vssd1 vssd1 vccd1 vccd1 _23339_/A sky130_fd_sc_hd__inv_2
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20549_ _20549_/A _25852_/Q vssd1 vssd1 vccd1 vccd1 _20554_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26056_ _26057_/CLK _26056_/D vssd1 vssd1 vccd1 vccd1 _26056_/Q sky130_fd_sc_hd__dfxtp_1
X_14070_ _14118_/A hold695/X vssd1 vssd1 vccd1 vccd1 hold696/A sky130_fd_sc_hd__nand2_1
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23268_ _23269_/B _23269_/A vssd1 vssd1 vccd1 vccd1 _23270_/A sky130_fd_sc_hd__or2_1
XFILLER_0_21_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25007_ _25594_/CLK hold994/X vssd1 vssd1 vccd1 vccd1 _25007_/Q sky130_fd_sc_hd__dfxtp_1
X_13021_ _26137_/Q _12907_/X _13020_/X vssd1 vssd1 vccd1 vccd1 _13021_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_123_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22219_ _25789_/Q _22219_/B vssd1 vssd1 vccd1 vccd1 _22219_/Y sky130_fd_sc_hd__nor2_1
X_23199_ _23199_/A _24745_/A _23199_/C vssd1 vssd1 vccd1 vccd1 _23200_/A sky130_fd_sc_hd__and3_4
X_14972_ _14972_/A _25421_/Q vssd1 vssd1 vccd1 vccd1 _14973_/B sky130_fd_sc_hd__nand2_1
X_17760_ _17761_/B _17760_/B _17973_/B vssd1 vssd1 vccd1 vccd1 _18019_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_156_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16711_ _16711_/A vssd1 vssd1 vccd1 vccd1 _16711_/X sky130_fd_sc_hd__buf_12
X_13923_ _13941_/A _13923_/B vssd1 vssd1 vccd1 vccd1 _13923_/Y sky130_fd_sc_hd__nand2_1
X_25909_ _25913_/CLK _25909_/D vssd1 vssd1 vccd1 vccd1 _25909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17691_ _17717_/A _17691_/B _17750_/B vssd1 vssd1 vccd1 vccd1 _17693_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_156_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_210_clk _26093_/CLK vssd1 vssd1 vccd1 vccd1 _26121_/CLK sky130_fd_sc_hd__clkbuf_16
X_16642_ _16642_/A _16642_/B vssd1 vssd1 vccd1 vccd1 _16643_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19430_ _19430_/A _21022_/B vssd1 vssd1 vccd1 vccd1 _19430_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13854_ _13941_/A _13854_/B vssd1 vssd1 vccd1 vccd1 _13854_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12805_ _26096_/Q _12748_/X _12804_/X vssd1 vssd1 vccd1 vccd1 _12805_/X sky130_fd_sc_hd__a21o_1
X_16573_ _16573_/A _16573_/B vssd1 vssd1 vccd1 vccd1 _16574_/B sky130_fd_sc_hd__and2_1
X_19361_ _20882_/A _19359_/Y _20886_/C vssd1 vssd1 vccd1 vccd1 _19449_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_85_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13785_ _13780_/Y _13784_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold848/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15524_ _22931_/B _15524_/B vssd1 vssd1 vccd1 vccd1 _22928_/B sky130_fd_sc_hd__xor2_1
X_18312_ _19066_/A _18312_/B vssd1 vssd1 vccd1 vccd1 _18312_/X sky130_fd_sc_hd__xor2_1
X_12736_ _25581_/Q _13465_/A vssd1 vssd1 vccd1 vccd1 _17008_/A sky130_fd_sc_hd__nor2_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19292_ _19308_/B _19378_/B vssd1 vssd1 vccd1 vccd1 _19294_/A sky130_fd_sc_hd__xnor2_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _18446_/A _18243_/B _18952_/C vssd1 vssd1 vccd1 vccd1 _18244_/C sky130_fd_sc_hd__nand3_1
X_15455_ _22863_/B _16369_/B vssd1 vssd1 vccd1 vccd1 _16424_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_139_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12667_ _12667_/A _24836_/B _12667_/C vssd1 vssd1 vccd1 vccd1 _12667_/X sky130_fd_sc_hd__and3_1
XFILLER_0_127_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14406_ _15464_/A vssd1 vssd1 vccd1 vccd1 _14406_/X sky130_fd_sc_hd__buf_6
X_18174_ _20944_/B _21940_/A vssd1 vssd1 vccd1 vccd1 _20935_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_182_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15386_ _15387_/B _16817_/A vssd1 vssd1 vccd1 vccd1 _15388_/A sky130_fd_sc_hd__nor2_1
X_12598_ _12598_/A vssd1 vssd1 vccd1 vccd1 _24972_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17125_ _17272_/A _17125_/B vssd1 vssd1 vccd1 vccd1 _17125_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_123_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14337_ _14337_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14337_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_41_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold507 hold507/A vssd1 vssd1 vccd1 vccd1 hold507/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold518 hold518/A vssd1 vssd1 vccd1 vccd1 hold518/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold529 hold529/A vssd1 vssd1 vccd1 vccd1 hold529/X sky130_fd_sc_hd__dlygate4sd3_1
X_17056_ _25626_/Q vssd1 vssd1 vccd1 vccd1 _20200_/B sky130_fd_sc_hd__inv_2
X_14268_ _14268_/A vssd1 vssd1 vccd1 vccd1 _14277_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_16007_ _16007_/A _16697_/B _16014_/A vssd1 vssd1 vccd1 vccd1 _16007_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_122_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13219_ _13207_/X _13217_/X _13192_/X _13218_/X vssd1 vssd1 vccd1 vccd1 _13219_/X
+ sky130_fd_sc_hd__o211a_1
X_14199_ _14194_/Y _14198_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold828/A sky130_fd_sc_hd__a21oi_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1207 _25552_/Q vssd1 vssd1 vccd1 vccd1 _16790_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_178_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17958_ _17958_/A _17958_/B _17958_/C vssd1 vssd1 vccd1 vccd1 _21766_/A sky130_fd_sc_hd__nand3_2
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1218 _13129_/X vssd1 vssd1 vccd1 vccd1 _25074_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1229 _13064_/X vssd1 vssd1 vccd1 vccd1 _25062_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16909_ _16935_/A _16914_/B vssd1 vssd1 vccd1 vccd1 _16911_/B sky130_fd_sc_hd__nand2_1
X_17889_ _25850_/Q _22130_/A vssd1 vssd1 vccd1 vccd1 _17898_/A sky130_fd_sc_hd__or2_2
XFILLER_0_75_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_201_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _26232_/CLK sky130_fd_sc_hd__clkbuf_16
X_19628_ _19627_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19629_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19559_ _19556_/Y _19559_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19559_/X sky130_fd_sc_hd__and3b_1
X_22570_ _22570_/A _22570_/B vssd1 vssd1 vccd1 vccd1 _23088_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_180_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21521_ _21520_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21521_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24240_ hold2335/X hold2004/X _24279_/S vssd1 vssd1 vccd1 vccd1 _24241_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_28_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21452_ _21452_/A _21452_/B vssd1 vssd1 vccd1 vccd1 _21453_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_146_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20403_ _20403_/A _25887_/Q vssd1 vssd1 vccd1 vccd1 _20409_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24171_ _24171_/A vssd1 vssd1 vccd1 vccd1 _26123_/D sky130_fd_sc_hd__clkbuf_1
X_21383_ _21433_/A _21386_/A vssd1 vssd1 vccd1 vccd1 _21384_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23122_ _23122_/A _23122_/B vssd1 vssd1 vccd1 vccd1 _23123_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20334_ _21498_/A _21169_/C vssd1 vssd1 vccd1 vccd1 _20335_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_102_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23053_ _23197_/A _23053_/B vssd1 vssd1 vccd1 vccd1 _23053_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_40_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20265_ _26283_/Q hold683/X vssd1 vssd1 vccd1 vccd1 _20265_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_179_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22004_ _22004_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _22004_/X sky130_fd_sc_hd__and2_1
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20196_ _20196_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _20196_/Y sky130_fd_sc_hd__nand2_1
Xhold2420 _26074_/Q vssd1 vssd1 vccd1 vccd1 hold2420/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2431 _25466_/Q vssd1 vssd1 vccd1 vccd1 _15654_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2442 _12682_/X vssd1 vssd1 vccd1 vccd1 _12683_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2453 _15062_/Y vssd1 vssd1 vccd1 vccd1 hold2453/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2464 _26195_/Q vssd1 vssd1 vccd1 vccd1 hold2464/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2475 _25922_/Q vssd1 vssd1 vccd1 vccd1 _23292_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1730 _25635_/Q vssd1 vssd1 vccd1 vccd1 _17583_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1741 _22537_/Y vssd1 vssd1 vccd1 vccd1 _25865_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2486 _24677_/X vssd1 vssd1 vccd1 vccd1 _24678_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23955_ _23955_/A vssd1 vssd1 vccd1 vccd1 _26053_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1752 _14975_/Y vssd1 vssd1 vccd1 vccd1 _14977_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2497 _25694_/Q vssd1 vssd1 vccd1 vccd1 _13371_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1763 _25596_/Q vssd1 vssd1 vccd1 vccd1 _17217_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1774 _22889_/Y vssd1 vssd1 vccd1 vccd1 _25882_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22906_ _22906_/A _22906_/B vssd1 vssd1 vccd1 vccd1 _22908_/A sky130_fd_sc_hd__nand2_1
Xhold1785 _25594_/Q vssd1 vssd1 vccd1 vccd1 _17190_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1796 _25867_/Q vssd1 vssd1 vccd1 vccd1 _22587_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23886_ hold1932/X _26033_/Q _23907_/S vssd1 vssd1 vccd1 vccd1 _23886_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25625_ _26216_/CLK _25625_/D vssd1 vssd1 vccd1 vccd1 _25625_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_168_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22837_ _22827_/Y _22836_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22837_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25556_ _25877_/CLK _25556_/D vssd1 vssd1 vccd1 vccd1 _25556_/Q sky130_fd_sc_hd__dfxtp_1
X_13570_ _26229_/Q _13426_/X _13468_/X _13569_/Y vssd1 vssd1 vccd1 vccd1 _13571_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22768_ _22768_/A _23001_/B _22768_/C vssd1 vssd1 vccd1 vccd1 _22768_/X sky130_fd_sc_hd__and3_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12521_ _13465_/B _14270_/B vssd1 vssd1 vccd1 vccd1 _12724_/B sky130_fd_sc_hd__or2_4
X_24507_ hold2571/X _26233_/Q _24510_/S vssd1 vssd1 vccd1 vccd1 _24507_/X sky130_fd_sc_hd__mux2_1
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21719_ _22058_/A _21719_/B vssd1 vssd1 vccd1 vccd1 _21719_/Y sky130_fd_sc_hd__nand2_1
X_25487_ _25939_/CLK hold773/X vssd1 vssd1 vccd1 vccd1 hold771/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22699_ _23168_/B vssd1 vssd1 vccd1 vccd1 _23167_/B sky130_fd_sc_hd__inv_2
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15240_ _26012_/Q _25948_/Q _15773_/S vssd1 vssd1 vccd1 vccd1 _15241_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_136_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24438_ _24438_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24439_/A sky130_fd_sc_hd__and2_1
XFILLER_0_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15171_ _26008_/Q _25944_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15172_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_152_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24369_ hold2274/X _26188_/Q _24433_/S vssd1 vssd1 vccd1 vccd1 _24369_/X sky130_fd_sc_hd__mux2_1
X_26108_ _26109_/CLK _26108_/D vssd1 vssd1 vccd1 vccd1 _26108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14122_ _26317_/Q _13988_/X _13981_/X _14121_/Y vssd1 vssd1 vccd1 vccd1 _14123_/B
+ sky130_fd_sc_hd__a22o_1
X_26039_ _26079_/CLK _26039_/D vssd1 vssd1 vccd1 vccd1 _26039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18930_ _25900_/Q _22691_/A vssd1 vssd1 vccd1 vccd1 _18938_/A sky130_fd_sc_hd__or2_2
XFILLER_0_31_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14053_ _18264_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14053_/Y sky130_fd_sc_hd__nor2_1
X_13004_ _26134_/Q _12907_/X _13003_/X vssd1 vssd1 vccd1 vccd1 _13004_/X sky130_fd_sc_hd__a21o_1
X_18861_ _18861_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18861_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17812_ _18528_/A _25727_/Q vssd1 vssd1 vccd1 vccd1 _17814_/A sky130_fd_sc_hd__nand2_1
X_18792_ _18792_/A _25765_/Q vssd1 vssd1 vccd1 vccd1 _18794_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14955_ _14955_/A _14955_/B vssd1 vssd1 vccd1 vccd1 _14956_/B sky130_fd_sc_hd__nand2_1
X_17743_ _17743_/A _17773_/B vssd1 vssd1 vccd1 vccd1 _17761_/B sky130_fd_sc_hd__nand2_1
X_13906_ _14000_/A hold683/X vssd1 vssd1 vccd1 vccd1 hold684/A sky130_fd_sc_hd__nand2_1
X_14886_ _22365_/B _15543_/B vssd1 vssd1 vccd1 vccd1 _14887_/A sky130_fd_sc_hd__nand2_1
X_17674_ _17674_/A vssd1 vssd1 vccd1 vccd1 _23208_/B sky130_fd_sc_hd__inv_2
X_19413_ _26234_/Q hold563/X vssd1 vssd1 vccd1 vccd1 _19413_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_186_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16625_ _16676_/A _16625_/B vssd1 vssd1 vccd1 vccd1 _16627_/A sky130_fd_sc_hd__or2_1
XFILLER_0_159_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13837_ hold627/X _13836_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold628/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16556_ _16564_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16556_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_186_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19344_ _19341_/Y _19344_/B _19980_/B vssd1 vssd1 vccd1 vccd1 _19344_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_58_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13768_ _13880_/A hold404/X vssd1 vssd1 vccd1 vccd1 hold405/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12719_ _12717_/X hold411/X _12558_/B vssd1 vssd1 vccd1 vccd1 hold412/A sky130_fd_sc_hd__a21oi_1
X_15507_ _26027_/Q _25963_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15508_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_127_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16487_ _16487_/A _16487_/B vssd1 vssd1 vccd1 vccd1 _16491_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_169_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19275_ _19275_/A _20663_/B vssd1 vssd1 vccd1 vccd1 _19275_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13699_ _13760_/A hold572/X vssd1 vssd1 vccd1 vccd1 hold573/A sky130_fd_sc_hd__nand2_1
XFILLER_0_116_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15438_ _15439_/A _15440_/A vssd1 vssd1 vccd1 vccd1 _15442_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_5_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18226_ _18226_/A _20993_/A vssd1 vssd1 vccd1 vccd1 _18576_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_155_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15369_ _15369_/A vssd1 vssd1 vccd1 vccd1 _16356_/A sky130_fd_sc_hd__inv_2
XFILLER_0_14_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18157_ _18159_/A _18159_/B vssd1 vssd1 vccd1 vccd1 _18158_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17108_ _17652_/A _17108_/B vssd1 vssd1 vccd1 vccd1 _17108_/X sky130_fd_sc_hd__xor2_1
Xhold304 hold304/A vssd1 vssd1 vccd1 vccd1 hold304/X sky130_fd_sc_hd__dlygate4sd3_1
X_18088_ _20630_/B _22250_/A vssd1 vssd1 vccd1 vccd1 _20624_/A sky130_fd_sc_hd__nand2_2
Xhold315 hold315/A vssd1 vssd1 vccd1 vccd1 hold315/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold326 hold326/A vssd1 vssd1 vccd1 vccd1 hold326/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 hold337/A vssd1 vssd1 vccd1 vccd1 hold337/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 hold348/A vssd1 vssd1 vccd1 vccd1 hold348/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17039_ _18212_/B _17039_/B vssd1 vssd1 vccd1 vccd1 _17423_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_111_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold359 hold359/A vssd1 vssd1 vccd1 vccd1 hold359/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20050_ _20050_/A _20050_/B vssd1 vssd1 vccd1 vccd1 _20052_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1004 _13103_/X vssd1 vssd1 vccd1 vccd1 _25069_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 _25064_/Q vssd1 vssd1 vccd1 vccd1 _17646_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1026 _12935_/X vssd1 vssd1 vccd1 vccd1 _25037_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1037 _25035_/Q vssd1 vssd1 vccd1 vccd1 _17435_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 _19668_/Y vssd1 vssd1 vccd1 vccd1 _25748_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 _25791_/Q vssd1 vssd1 vccd1 vccd1 _20699_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23740_ _23740_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23741_/A sky130_fd_sc_hd__and2_1
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20952_ _20952_/A _20952_/B _20952_/C vssd1 vssd1 vccd1 vccd1 _20953_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_96_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23671_ hold2251/X hold2243/X _23677_/S vssd1 vssd1 vccd1 vccd1 _23672_/A sky130_fd_sc_hd__mux2_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20883_ _20883_/A _20883_/B vssd1 vssd1 vccd1 vccd1 _20886_/A sky130_fd_sc_hd__nand2_1
X_25410_ _26001_/CLK _25410_/D vssd1 vssd1 vccd1 vccd1 _25410_/Q sky130_fd_sc_hd__dfxtp_1
X_22622_ _23120_/B vssd1 vssd1 vccd1 vccd1 _23119_/B sky130_fd_sc_hd__inv_2
XFILLER_0_36_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25341_ _26298_/CLK hold268/X vssd1 vssd1 vccd1 vccd1 hold266/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22553_ _15192_/B _22387_/B _14273_/X vssd1 vssd1 vccd1 vccd1 _22553_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21504_ _26327_/Q hold823/X vssd1 vssd1 vccd1 vccd1 _21504_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_134_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25272_ _26103_/CLK hold283/X vssd1 vssd1 vccd1 vccd1 hold281/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22484_ _22475_/Y _22483_/Y _23197_/A vssd1 vssd1 vccd1 vccd1 _22484_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_17_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24223_ _24223_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24224_/A sky130_fd_sc_hd__and2_1
XFILLER_0_161_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21435_ _21435_/A _21435_/B _21435_/C vssd1 vssd1 vccd1 vccd1 _21436_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24154_ hold2281/X _26118_/Q _24203_/S vssd1 vssd1 vccd1 vccd1 _24154_/X sky130_fd_sc_hd__mux2_1
X_21366_ _21418_/A vssd1 vssd1 vccd1 vccd1 _21417_/A sky130_fd_sc_hd__inv_2
XFILLER_0_101_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23105_ _23105_/A _23105_/B vssd1 vssd1 vccd1 vccd1 _23106_/B sky130_fd_sc_hd__nand2_1
X_20317_ _20317_/A vssd1 vssd1 vccd1 vccd1 _20318_/B sky130_fd_sc_hd__inv_2
XFILLER_0_82_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24085_ _24085_/A vssd1 vssd1 vccd1 vccd1 _26095_/D sky130_fd_sc_hd__clkbuf_1
Xhold860 hold860/A vssd1 vssd1 vccd1 vccd1 hold860/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_21297_ _21296_/B _21297_/B _21297_/C vssd1 vssd1 vccd1 vccd1 _21298_/B sky130_fd_sc_hd__nand3b_1
Xhold871 hold871/A vssd1 vssd1 vccd1 vccd1 hold871/X sky130_fd_sc_hd__buf_1
Xhold882 hold882/A vssd1 vssd1 vccd1 vccd1 hold882/X sky130_fd_sc_hd__dlygate4sd3_1
X_23036_ _23027_/Y _23035_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _23036_/X sky130_fd_sc_hd__a21o_1
Xhold893 hold893/A vssd1 vssd1 vccd1 vccd1 hold893/X sky130_fd_sc_hd__dlygate4sd3_1
X_20248_ _20248_/A _20248_/B vssd1 vssd1 vccd1 vccd1 _20251_/A sky130_fd_sc_hd__nand2_1
X_20179_ _20180_/A _20180_/C _20180_/B vssd1 vssd1 vccd1 vccd1 _20181_/A sky130_fd_sc_hd__a21o_1
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2250 _24237_/X vssd1 vssd1 vccd1 vccd1 _24238_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2261 _12628_/Y vssd1 vssd1 vccd1 vccd1 _12630_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2272 _12596_/Y vssd1 vssd1 vccd1 vccd1 _12597_/C sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24987_ _24990_/CLK _24987_/D vssd1 vssd1 vccd1 vccd1 _24987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2283 _25941_/Q vssd1 vssd1 vccd1 vccd1 hold2283/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2294 _26194_/Q vssd1 vssd1 vccd1 vccd1 hold2294/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1560 _13394_/X vssd1 vssd1 vccd1 vccd1 _25117_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ _14900_/A _14740_/B vssd1 vssd1 vccd1 vccd1 _14740_/Y sky130_fd_sc_hd__nand2_1
Xhold1571 _21316_/Y vssd1 vssd1 vccd1 vccd1 _25812_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23938_ hold2507/X hold2471/X _24001_/S vssd1 vssd1 vccd1 vccd1 _23939_/A sky130_fd_sc_hd__mux2_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1582 _25615_/Q vssd1 vssd1 vccd1 vccd1 _17438_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1593 _20308_/Y vssd1 vssd1 vccd1 vccd1 _25781_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ _14669_/Y hold63/X _14646_/X vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__a21oi_1
X_23869_ _23869_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23870_/A sky130_fd_sc_hd__and2_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16410_ hold894/X vssd1 vssd1 vccd1 vccd1 _16413_/B sky130_fd_sc_hd__inv_2
XFILLER_0_39_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25608_ _26240_/CLK _25608_/D vssd1 vssd1 vccd1 vccd1 _25608_/Q sky130_fd_sc_hd__dfxtp_4
X_13622_ _13703_/A _13622_/B vssd1 vssd1 vccd1 vccd1 _13622_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_156_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17390_ _19546_/A _17390_/B vssd1 vssd1 vccd1 vccd1 _17622_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16341_ _16341_/A _16697_/B _16341_/C vssd1 vssd1 vccd1 vccd1 _16341_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_66_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25539_ _25539_/CLK hold577/X vssd1 vssd1 vccd1 vccd1 hold575/A sky130_fd_sc_hd__dfxtp_1
X_13553_ hold582/X _13552_/Y _12558_/B vssd1 vssd1 vccd1 vccd1 hold583/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12504_ _12559_/A hold4/X vssd1 vssd1 vccd1 vccd1 _23597_/A sky130_fd_sc_hd__nor2_1
X_19060_ _19060_/A _19060_/B vssd1 vssd1 vccd1 vccd1 _19060_/X sky130_fd_sc_hd__xor2_1
X_16272_ _16272_/A _16272_/B vssd1 vssd1 vccd1 vccd1 _16273_/A sky130_fd_sc_hd__nor2_1
X_13484_ _13583_/A _13484_/B vssd1 vssd1 vccd1 vccd1 _13484_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_42_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15223_ _26011_/Q _25947_/Q _15773_/S vssd1 vssd1 vccd1 vccd1 _15224_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18011_ _18252_/A _18011_/B vssd1 vssd1 vccd1 vccd1 _18011_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15154_ _22504_/B _15154_/B vssd1 vssd1 vccd1 vccd1 _22501_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_22_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14105_ _14100_/Y _14104_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold795/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15085_ _15085_/A _15085_/B vssd1 vssd1 vccd1 vccd1 _15085_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19962_ _19960_/X _19961_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19962_/Y sky130_fd_sc_hd__a21oi_1
X_14036_ _14061_/A _14036_/B vssd1 vssd1 vccd1 vccd1 _14036_/Y sky130_fd_sc_hd__nand2_1
X_18913_ _18954_/A _25771_/Q vssd1 vssd1 vccd1 vccd1 _18915_/A sky130_fd_sc_hd__nand2_1
X_19893_ _26268_/Q hold677/X vssd1 vssd1 vccd1 vccd1 _19893_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18844_ _25704_/Q _20752_/B vssd1 vssd1 vccd1 vccd1 _18847_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_101_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18775_ _20605_/B _22490_/A vssd1 vssd1 vccd1 vccd1 _20596_/A sky130_fd_sc_hd__nand2_2
X_15987_ _15987_/A _15987_/B vssd1 vssd1 vccd1 vccd1 _15989_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_166_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17726_ _17726_/A _17764_/B _17726_/C vssd1 vssd1 vccd1 vccd1 _17728_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_145_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14938_ _14938_/A _14938_/B vssd1 vssd1 vccd1 vccd1 _14939_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17657_ _17655_/Y _17656_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _17657_/Y sky130_fd_sc_hd__a21oi_1
X_14869_ _14869_/A vssd1 vssd1 vccd1 vccd1 _15058_/A sky130_fd_sc_hd__inv_2
XFILLER_0_175_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16608_ _16608_/A _16608_/B vssd1 vssd1 vccd1 vccd1 _16629_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17588_ _17586_/X _17528_/X _17587_/X vssd1 vssd1 vccd1 vccd1 _17590_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19327_ _26228_/Q _12537_/B hold560/X vssd1 vssd1 vccd1 vccd1 _19327_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16539_ _16698_/A _16539_/B vssd1 vssd1 vccd1 vccd1 _16539_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_128_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19258_ _20624_/A _22248_/B _25598_/Q vssd1 vssd1 vccd1 vccd1 _20628_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_183_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18209_ _18207_/X _17528_/X _18208_/X vssd1 vssd1 vccd1 vccd1 _18211_/A sky130_fd_sc_hd__a21o_1
X_19189_ _20428_/A _17853_/B _20432_/C vssd1 vssd1 vccd1 vccd1 _19280_/B sky130_fd_sc_hd__o21a_4
XFILLER_0_143_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21220_ _21662_/B _21610_/C vssd1 vssd1 vccd1 vccd1 _21222_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_143_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold101 hold101/A vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold112 hold112/A vssd1 vssd1 vccd1 vccd1 hold112/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 hold123/A vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold134 hold134/A vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21151_ _21151_/A _21151_/B vssd1 vssd1 vccd1 vccd1 _21153_/A sky130_fd_sc_hd__nand2_1
Xhold145 hold145/A vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 hold156/A vssd1 vssd1 vccd1 vccd1 hold156/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 hold167/A vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 hold178/A vssd1 vssd1 vccd1 vccd1 hold178/X sky130_fd_sc_hd__dlygate4sd3_1
X_20102_ _25879_/Q _20102_/B _20102_/C vssd1 vssd1 vccd1 vccd1 _20106_/B sky130_fd_sc_hd__nand3b_1
Xhold189 hold189/A vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21082_ _21082_/A _21082_/B vssd1 vssd1 vccd1 vccd1 _21580_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_106_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24910_ _24950_/B _24959_/C _23484_/B _24870_/B vssd1 vssd1 vccd1 vccd1 _24910_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20033_ _22704_/A vssd1 vssd1 vccd1 vccd1 _20730_/B sky130_fd_sc_hd__buf_6
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25890_ _26080_/CLK _25890_/D vssd1 vssd1 vccd1 vccd1 _25890_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24841_ _15198_/A _15213_/B _24860_/S vssd1 vssd1 vccd1 vccd1 _24841_/X sky130_fd_sc_hd__mux2_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24772_ hold2641/X hold2636/X _24817_/S vssd1 vssd1 vccd1 vccd1 _24773_/A sky130_fd_sc_hd__mux2_1
X_21984_ _19532_/A _21983_/A _21983_/Y vssd1 vssd1 vccd1 vccd1 _21986_/A sky130_fd_sc_hd__o21ai_2
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23723_ hold2049/X _25980_/Q _23754_/S vssd1 vssd1 vccd1 vccd1 _23723_/X sky130_fd_sc_hd__mux2_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20935_ _20935_/A _21938_/B vssd1 vssd1 vccd1 vccd1 _20936_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23654_ _23654_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23655_/A sky130_fd_sc_hd__and2_1
XFILLER_0_113_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20866_ _21448_/C _21677_/A vssd1 vssd1 vccd1 vccd1 _20868_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22605_ _26051_/Q vssd1 vssd1 vccd1 vccd1 _22606_/A sky130_fd_sc_hd__inv_2
XFILLER_0_64_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23585_ _25935_/Q _25934_/Q _25933_/Q _25932_/Q vssd1 vssd1 vccd1 vccd1 _23586_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_181_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20797_ _20797_/A _20797_/B vssd1 vssd1 vccd1 vccd1 _20799_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_113_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25324_ _26279_/CLK hold82/X vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22536_ _22561_/A _22536_/B vssd1 vssd1 vccd1 vccd1 _22536_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25255_ _25827_/CLK hold652/X vssd1 vssd1 vccd1 vccd1 hold650/A sky130_fd_sc_hd__dfxtp_1
X_22467_ _22468_/B _22468_/A vssd1 vssd1 vccd1 vccd1 _22469_/A sky130_fd_sc_hd__or2_1
X_24206_ _24835_/S vssd1 vssd1 vccd1 vccd1 _24279_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_122_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21418_ _21418_/A _21466_/A vssd1 vssd1 vccd1 vccd1 _21419_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_60_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25186_ _26269_/CLK hold805/X vssd1 vssd1 vccd1 vccd1 hold803/A sky130_fd_sc_hd__dfxtp_1
X_22398_ _22975_/B vssd1 vssd1 vccd1 vccd1 _22974_/B sky130_fd_sc_hd__inv_2
XFILLER_0_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24137_ _24137_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24138_/A sky130_fd_sc_hd__and2_1
XFILLER_0_32_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21349_ _21710_/B _21402_/A vssd1 vssd1 vccd1 vccd1 _21351_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_102_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24068_ hold1911/X hold992/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24069_/A sky130_fd_sc_hd__mux2_1
Xhold690 hold690/A vssd1 vssd1 vccd1 vccd1 hold690/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15910_ _15921_/A _15911_/A vssd1 vssd1 vccd1 vccd1 _15910_/X sky130_fd_sc_hd__or2_1
X_23019_ _23019_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _23019_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_159_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16890_ _16890_/A _16890_/B vssd1 vssd1 vccd1 vccd1 _16890_/Y sky130_fd_sc_hd__nand2_1
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _16676_/A vssd1 vssd1 vccd1 vccd1 _16401_/C sky130_fd_sc_hd__inv_8
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2080 _26034_/Q vssd1 vssd1 vccd1 vccd1 hold2080/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2091 _24379_/X vssd1 vssd1 vccd1 vccd1 _24380_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18560_ _18641_/A _19402_/A vssd1 vssd1 vccd1 vccd1 _18560_/Y sky130_fd_sc_hd__nand2_1
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ _16970_/B vssd1 vssd1 vccd1 vccd1 _23159_/B sky130_fd_sc_hd__inv_2
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ hold899/X _12907_/X _12983_/X vssd1 vssd1 vccd1 vccd1 hold900/A sky130_fd_sc_hd__a21o_1
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1390 _12829_/X vssd1 vssd1 vccd1 vccd1 _25017_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17511_ _17509_/Y _17510_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _25625_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14723_ _15839_/A _14723_/B vssd1 vssd1 vccd1 vccd1 _21831_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_115_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18491_ _20062_/C _22122_/A vssd1 vssd1 vccd1 vccd1 _20054_/A sky130_fd_sc_hd__nand2_2
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14654_ _14654_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _14654_/Y sky130_fd_sc_hd__nand2_1
X_17442_ _17624_/A _17442_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17442_/X sky130_fd_sc_hd__and3_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13605_ _14170_/A vssd1 vssd1 vccd1 vccd1 _13605_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_185_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17373_ _17393_/A _17373_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17373_/X sky130_fd_sc_hd__and3_1
X_14585_ _14585_/A hold209/X vssd1 vssd1 vccd1 vccd1 hold210/A sky130_fd_sc_hd__nand2_1
XFILLER_0_156_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19112_ _19186_/A _19112_/B vssd1 vssd1 vccd1 vccd1 _19112_/Y sky130_fd_sc_hd__nand2_1
X_16324_ _16324_/A _16336_/B vssd1 vssd1 vccd1 vccd1 _16324_/Y sky130_fd_sc_hd__nand2_1
X_13536_ _13642_/A hold458/X vssd1 vssd1 vccd1 vccd1 hold459/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16255_ _16264_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16255_/Y sky130_fd_sc_hd__nand2_1
X_19043_ _19186_/A _19844_/A vssd1 vssd1 vccd1 vccd1 _19043_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_54_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13467_ _13467_/A vssd1 vssd1 vccd1 vccd1 _14170_/A sky130_fd_sc_hd__clkinv_16
XFILLER_0_36_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ _26010_/Q _25946_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15207_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16186_ _16212_/A hold860/X vssd1 vssd1 vccd1 vccd1 _16186_/Y sky130_fd_sc_hd__nand2_1
X_13398_ _26201_/Q _13239_/X _13397_/X vssd1 vssd1 vccd1 vccd1 _13398_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_26_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15137_ _15137_/A _15776_/B vssd1 vssd1 vccd1 vccd1 _15138_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_50_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15068_ _15067_/X _15068_/B vssd1 vssd1 vccd1 vccd1 _15069_/A sky130_fd_sc_hd__nand2b_1
X_19945_ _19944_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19947_/A
+ sky130_fd_sc_hd__a211o_1
X_14019_ hold504/X _14018_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold505/A sky130_fd_sc_hd__a21oi_1
X_19876_ _19874_/X _19875_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19876_/Y sky130_fd_sc_hd__a21oi_1
X_18827_ _18827_/A _18827_/B vssd1 vssd1 vccd1 vccd1 _22563_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_179_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18758_ _18758_/A _18758_/B vssd1 vssd1 vccd1 vccd1 _18758_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_179_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17709_ _17709_/A _17738_/A _17709_/C vssd1 vssd1 vccd1 vccd1 _17759_/C sky130_fd_sc_hd__nand3_1
X_18689_ _18951_/A _18693_/B vssd1 vssd1 vccd1 vccd1 _18691_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_176_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20720_ _20720_/A _20720_/B _20720_/C vssd1 vssd1 vccd1 vccd1 _20721_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20651_ _20651_/A _21302_/C _20651_/C vssd1 vssd1 vccd1 vccd1 _20652_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_19_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23370_ _23372_/B _23372_/A vssd1 vssd1 vccd1 vccd1 _23376_/A sky130_fd_sc_hd__nor2_1
X_20582_ _20582_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _20582_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_162_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22321_ _22319_/Y _22320_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _22321_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25040_ _26122_/CLK _25040_/D vssd1 vssd1 vccd1 vccd1 _25040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22252_ _25854_/Q _22253_/A vssd1 vssd1 vccd1 vccd1 _22254_/A sky130_fd_sc_hd__or2_1
XFILLER_0_143_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21203_ _21203_/A vssd1 vssd1 vccd1 vccd1 _21203_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_108_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22183_ _25880_/Q _22184_/A vssd1 vssd1 vccd1 vccd1 _22185_/A sky130_fd_sc_hd__or2_1
XFILLER_0_2_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21134_ _21136_/C vssd1 vssd1 vccd1 vccd1 _21135_/B sky130_fd_sc_hd__inv_2
Xclkbuf_2_2_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_25942_ _26073_/CLK _25942_/D vssd1 vssd1 vccd1 vccd1 _25942_/Q sky130_fd_sc_hd__dfxtp_1
X_21065_ _21716_/A vssd1 vssd1 vccd1 vccd1 _21636_/A sky130_fd_sc_hd__buf_6
XFILLER_0_100_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20016_ _20018_/C vssd1 vssd1 vccd1 vccd1 _20017_/B sky130_fd_sc_hd__inv_2
X_25873_ _25877_/CLK _25873_/D vssd1 vssd1 vccd1 vccd1 _25873_/Q sky130_fd_sc_hd__dfxtp_4
X_24824_ _24824_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24825_/A sky130_fd_sc_hd__and2_1
XFILLER_0_119_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24755_ _24755_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24756_/A sky130_fd_sc_hd__and2_1
X_21967_ _22653_/A _21967_/B vssd1 vssd1 vccd1 vccd1 _21967_/X sky130_fd_sc_hd__or2_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23706_ _23706_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23707_/A sky130_fd_sc_hd__and2_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20918_ _21483_/B vssd1 vssd1 vccd1 vccd1 _21480_/C sky130_fd_sc_hd__inv_2
X_24686_ hold2612/X hold2596/X _24740_/S vssd1 vssd1 vccd1 vccd1 _24687_/A sky130_fd_sc_hd__mux2_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21898_ _21895_/Y _21896_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _21898_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23637_ _23637_/A vssd1 vssd1 vccd1 vccd1 _25951_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20849_ _20848_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20849_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14370_ _14370_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14370_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23568_ _24922_/S hold221/A _23567_/X vssd1 vssd1 vccd1 vccd1 _23568_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25307_ _26135_/CLK hold304/X vssd1 vssd1 vccd1 vccd1 hold302/A sky130_fd_sc_hd__dfxtp_1
X_13321_ _13315_/X _13319_/X _13300_/X _13320_/X vssd1 vssd1 vccd1 vccd1 _13321_/X
+ sky130_fd_sc_hd__o211a_1
X_22519_ _22519_/A _22519_/B vssd1 vssd1 vccd1 vccd1 _23056_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_135_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26287_ _26287_/CLK _26287_/D vssd1 vssd1 vccd1 vccd1 _26287_/Q sky130_fd_sc_hd__dfxtp_2
X_23499_ hold131/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23499_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_80_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ _16040_/A _16040_/B vssd1 vssd1 vccd1 vccd1 _16042_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_162_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252_ _13207_/X _13250_/X _13192_/X _13251_/X vssd1 vssd1 vccd1 vccd1 _13252_/X
+ sky130_fd_sc_hd__o211a_1
X_25238_ _25689_/CLK hold436/X vssd1 vssd1 vccd1 vccd1 hold434/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13183_ _26295_/Q _19289_/A vssd1 vssd1 vccd1 vccd1 _14548_/A sky130_fd_sc_hd__xor2_1
X_25169_ _25748_/CLK hold544/X vssd1 vssd1 vccd1 vccd1 hold542/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17991_ _20553_/B _22192_/A vssd1 vssd1 vccd1 vccd1 _20546_/A sky130_fd_sc_hd__nand2_2
X_19730_ _20400_/A _22370_/B _25631_/Q vssd1 vssd1 vccd1 vccd1 _20405_/C sky130_fd_sc_hd__nand3_1
X_16942_ _16939_/Y _16940_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _16942_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19661_ _20199_/A _19659_/Y _20204_/C vssd1 vssd1 vccd1 vccd1 _19749_/B sky130_fd_sc_hd__o21a_2
X_16873_ _16871_/Y _16872_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16873_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18612_ _18612_/A _18612_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18613_/C sky130_fd_sc_hd__nand3_1
X_15824_ _15824_/A _15824_/B vssd1 vssd1 vccd1 vccd1 _15829_/B sky130_fd_sc_hd__and2_1
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19592_ _19593_/B _19593_/A vssd1 vssd1 vccd1 vccd1 _19592_/X sky130_fd_sc_hd__or2_1
XFILLER_0_189_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18543_ _20163_/B _19644_/A vssd1 vssd1 vccd1 vccd1 _18544_/B sky130_fd_sc_hd__nand2_1
X_15755_ _15755_/A _15810_/B vssd1 vssd1 vccd1 vccd1 _15756_/B sky130_fd_sc_hd__nand2_2
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ _12891_/X _14422_/A _12909_/X _25624_/Q vssd1 vssd1 vccd1 vccd1 _12967_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14706_ _14712_/B _21760_/A vssd1 vssd1 vccd1 vccd1 _21759_/B sky130_fd_sc_hd__xnor2_2
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18474_ _18474_/A _18474_/B vssd1 vssd1 vccd1 vccd1 _18474_/X sky130_fd_sc_hd__xor2_1
X_15686_ _15686_/A vssd1 vssd1 vccd1 vccd1 _16605_/A sky130_fd_sc_hd__inv_2
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12898_ _12891_/X _14379_/A _12752_/X _25611_/Q vssd1 vssd1 vccd1 vccd1 _12898_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ _17423_/X _17241_/X _17424_/X vssd1 vssd1 vccd1 vccd1 _17426_/A sky130_fd_sc_hd__a21o_1
X_14637_ _14635_/Y hold450/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold451/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17356_ _17467_/A _17356_/B vssd1 vssd1 vccd1 vccd1 _17356_/Y sky130_fd_sc_hd__nand2_1
X_14568_ _14566_/Y hold306/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold307/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16307_ _16336_/A _16307_/B vssd1 vssd1 vccd1 vccd1 _16333_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13519_ _26221_/Q _13426_/X _13468_/X _13518_/Y vssd1 vssd1 vccd1 vccd1 _13520_/B
+ sky130_fd_sc_hd__a22o_1
X_17287_ _17284_/Y _17286_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _17287_/Y sky130_fd_sc_hd__a21oi_1
X_14499_ _14497_/Y hold249/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold250/A sky130_fd_sc_hd__a21oi_1
X_19026_ _19026_/A _19026_/B _22786_/A vssd1 vssd1 vccd1 vccd1 _19026_/X sky130_fd_sc_hd__and3_1
X_16238_ _16238_/A _16238_/B vssd1 vssd1 vccd1 vccd1 _16240_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16169_ _16182_/B _16169_/B vssd1 vssd1 vccd1 vccd1 _16172_/B sky130_fd_sc_hd__and2_1
XFILLER_0_140_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19928_ _19928_/A _19928_/B vssd1 vssd1 vccd1 vccd1 _19928_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19859_ _20751_/A _18847_/A _20756_/C vssd1 vssd1 vccd1 vccd1 _19937_/A sky130_fd_sc_hd__o21a_1
X_22870_ _22870_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _22870_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21821_ _21821_/A _21821_/B vssd1 vssd1 vccd1 vccd1 _21823_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_167_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24540_ _24540_/A vssd1 vssd1 vccd1 vccd1 _26243_/D sky130_fd_sc_hd__clkbuf_1
X_21752_ _22891_/A vssd1 vssd1 vccd1 vccd1 _22745_/A sky130_fd_sc_hd__inv_2
XFILLER_0_176_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20703_ _20705_/B _20705_/C vssd1 vssd1 vccd1 vccd1 _20704_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_109_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24471_ hold2715/X hold2565/X _24510_/S vssd1 vssd1 vccd1 vccd1 _24472_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_47_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21683_ _21682_/Y _21203_/X _20986_/A _20957_/A vssd1 vssd1 vccd1 vccd1 _21683_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26210_ _26335_/CLK _26210_/D vssd1 vssd1 vccd1 vccd1 _26210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23422_ hold107/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23422_/X sky130_fd_sc_hd__or2b_1
X_20634_ _20634_/A _22513_/B vssd1 vssd1 vccd1 vccd1 _20635_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26141_ _26142_/CLK _26141_/D vssd1 vssd1 vccd1 vccd1 _26141_/Q sky130_fd_sc_hd__dfxtp_1
X_23353_ _23353_/A vssd1 vssd1 vccd1 vccd1 _25933_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20565_ _20565_/A _20565_/B vssd1 vssd1 vccd1 vccd1 _20567_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22304_ _22907_/B vssd1 vssd1 vccd1 vccd1 _22906_/B sky130_fd_sc_hd__inv_2
XFILLER_0_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26072_ _26073_/CLK _26072_/D vssd1 vssd1 vccd1 vccd1 _26072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23284_ _23284_/A hold832/X vssd1 vssd1 vccd1 vccd1 _23307_/A sky130_fd_sc_hd__nor2b_2
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20496_ _20496_/A _20496_/B vssd1 vssd1 vccd1 vccd1 _20497_/A sky130_fd_sc_hd__nand2_1
X_25023_ _26109_/CLK _25023_/D vssd1 vssd1 vccd1 vccd1 _25023_/Q sky130_fd_sc_hd__dfxtp_1
X_22235_ _22235_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _22235_/X sky130_fd_sc_hd__and2_1
XFILLER_0_14_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22166_ _22166_/A _22166_/B vssd1 vssd1 vccd1 vccd1 _23106_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21117_ _21117_/A _21117_/B _21117_/C vssd1 vssd1 vccd1 vccd1 _21118_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_100_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22097_ _22097_/A _22097_/B vssd1 vssd1 vccd1 vccd1 _22097_/Y sky130_fd_sc_hd__nand2_1
X_25925_ _25925_/CLK hold898/X vssd1 vssd1 vccd1 vccd1 hold896/A sky130_fd_sc_hd__dfxtp_1
X_21048_ _21048_/A _21048_/B vssd1 vssd1 vccd1 vccd1 _21051_/B sky130_fd_sc_hd__nand2_1
X_13870_ _17665_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13870_/Y sky130_fd_sc_hd__nor2_1
X_25856_ _26339_/CLK _25856_/D vssd1 vssd1 vccd1 vccd1 _25856_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12821_ _14064_/A vssd1 vssd1 vccd1 vccd1 _12974_/B sky130_fd_sc_hd__buf_8
X_24807_ _24807_/A vssd1 vssd1 vccd1 vccd1 _26330_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22999_ _22999_/A _22999_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _23001_/A sky130_fd_sc_hd__or3_1
X_25787_ _26287_/CLK _25787_/D vssd1 vssd1 vccd1 vccd1 _25787_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_9_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15540_ _22948_/B _15540_/B vssd1 vssd1 vccd1 vccd1 _22945_/B sky130_fd_sc_hd__xor2_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ _13242_/A vssd1 vssd1 vccd1 vccd1 _12752_/X sky130_fd_sc_hd__buf_8
XFILLER_0_55_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24738_ _24738_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24739_/A sky130_fd_sc_hd__and2_1
XFILLER_0_167_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15471_ _16851_/B vssd1 vssd1 vccd1 vccd1 _22882_/B sky130_fd_sc_hd__inv_2
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12683_ _12683_/A vssd1 vssd1 vccd1 vccd1 _24988_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24669_ _24669_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24670_/A sky130_fd_sc_hd__and2_1
XFILLER_0_132_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17210_ _20635_/B _25893_/Q _25829_/Q vssd1 vssd1 vccd1 vccd1 _17211_/B sky130_fd_sc_hd__mux2_2
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _14422_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14422_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_139_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18190_ _18190_/A _25783_/Q _18190_/C vssd1 vssd1 vccd1 vccd1 _20357_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14353_ _14404_/A hold290/X vssd1 vssd1 vccd1 vccd1 hold291/A sky130_fd_sc_hd__nand2_1
X_17141_ _20625_/B _25854_/Q _25790_/Q vssd1 vssd1 vccd1 vccd1 _17142_/B sky130_fd_sc_hd__mux2_2
X_26339_ _26339_/CLK _26339_/D vssd1 vssd1 vccd1 vccd1 _26339_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_123_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13304_ _26314_/Q _19560_/A vssd1 vssd1 vccd1 vccd1 _14608_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_107_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17072_ _25627_/Q vssd1 vssd1 vccd1 vccd1 _20236_/B sky130_fd_sc_hd__inv_2
XFILLER_0_52_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14284_ _14590_/A vssd1 vssd1 vccd1 vccd1 _14588_/A sky130_fd_sc_hd__inv_2
XFILLER_0_123_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16023_ _16023_/A _16023_/B vssd1 vssd1 vccd1 vccd1 _16024_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_122_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13235_ _13220_/X _14572_/A _13067_/X _19402_/A vssd1 vssd1 vccd1 vccd1 _13235_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13166_ _13049_/X _14539_/A _13067_/X _19244_/A vssd1 vssd1 vccd1 vccd1 _13166_/X
+ sky130_fd_sc_hd__a22o_1
X_13097_ _17914_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13097_/X sky130_fd_sc_hd__or2_1
X_17974_ _17974_/A _17974_/B vssd1 vssd1 vccd1 vccd1 _17976_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_100_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19713_ _19712_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19714_/B
+ sky130_fd_sc_hd__a211o_1
X_16925_ _16925_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16925_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_137_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19644_ _19644_/A _20163_/B vssd1 vssd1 vccd1 vccd1 _19644_/Y sky130_fd_sc_hd__nor2_1
X_16856_ _16854_/X _16711_/X _16855_/Y _25883_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16857_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_172_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15807_ _15807_/A vssd1 vssd1 vccd1 vccd1 _15816_/B sky130_fd_sc_hd__inv_2
X_19575_ _21290_/A _22065_/B _25620_/Q vssd1 vssd1 vccd1 vccd1 _21294_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_189_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16787_ _16787_/A _16787_/B vssd1 vssd1 vccd1 vccd1 _16787_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_137_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13999_ hold624/X _13998_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold625/A sky130_fd_sc_hd__a21oi_1
X_18526_ _18529_/A _25752_/Q _18529_/C vssd1 vssd1 vccd1 vccd1 _18527_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_88_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15738_ _15738_/A _15810_/B vssd1 vssd1 vccd1 vccd1 _15739_/B sky130_fd_sc_hd__nand2_2
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18457_ _18457_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18457_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15669_ _23060_/B _15810_/B vssd1 vssd1 vccd1 vccd1 _15670_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17408_ _17406_/Y _17407_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _25612_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18388_ _18388_/A _18388_/B _18388_/C vssd1 vssd1 vccd1 vccd1 _21983_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_172_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17339_ _21102_/B _25869_/Q _21844_/A vssd1 vssd1 vccd1 vccd1 _17340_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20350_ _20350_/A _20350_/B vssd1 vssd1 vccd1 vccd1 _20354_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19009_ _19007_/Y _19008_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25698_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20281_ _20281_/A _20281_/B _20281_/C vssd1 vssd1 vccd1 vccd1 _20282_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22020_ _22020_/A _22756_/B vssd1 vssd1 vccd1 vccd1 _22021_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_144_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2602 _26295_/Q vssd1 vssd1 vccd1 vccd1 hold2602/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2613 _26294_/Q vssd1 vssd1 vccd1 vccd1 hold2613/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2624 _15536_/Y vssd1 vssd1 vccd1 vccd1 _25459_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2635 _24627_/X vssd1 vssd1 vccd1 vccd1 _24628_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1901 _23831_/X vssd1 vssd1 vccd1 vccd1 _23832_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
X_23971_ hold2504/X _26059_/Q _24001_/S vssd1 vssd1 vccd1 vccd1 _23971_/X sky130_fd_sc_hd__mux2_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2646 _26268_/Q vssd1 vssd1 vccd1 vccd1 hold2646/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1912 _26040_/Q vssd1 vssd1 vccd1 vccd1 hold1912/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2657 _26242_/Q vssd1 vssd1 vccd1 vccd1 hold2657/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2668 _25447_/Q vssd1 vssd1 vccd1 vccd1 _15313_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1923 _12519_/X vssd1 vssd1 vccd1 vccd1 _25000_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2679 _23239_/Y vssd1 vssd1 vccd1 vccd1 _25911_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1934 _26041_/Q vssd1 vssd1 vccd1 vccd1 hold1934/X sky130_fd_sc_hd__dlygate4sd3_1
X_22922_ _23074_/A vssd1 vssd1 vccd1 vccd1 _22923_/B sky130_fd_sc_hd__inv_2
Xhold1945 _26279_/Q vssd1 vssd1 vccd1 vccd1 hold1945/X sky130_fd_sc_hd__buf_1
X_25710_ _25711_/CLK _25710_/D vssd1 vssd1 vccd1 vccd1 _25710_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1956 _24151_/X vssd1 vssd1 vccd1 vccd1 _24152_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1967 _26006_/Q vssd1 vssd1 vccd1 vccd1 hold1967/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1978 _26042_/Q vssd1 vssd1 vccd1 vccd1 hold1978/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1989 _26202_/Q vssd1 vssd1 vccd1 vccd1 hold1989/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22853_ _22853_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _22853_/Y sky130_fd_sc_hd__nand2_1
X_25641_ _26148_/CLK _25641_/D vssd1 vssd1 vccd1 vccd1 _25641_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_116_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21804_ _19331_/A _21803_/A _21803_/Y vssd1 vssd1 vccd1 vccd1 _21806_/A sky130_fd_sc_hd__o21ai_1
X_25572_ _25893_/CLK _25572_/D vssd1 vssd1 vccd1 vccd1 _25572_/Q sky130_fd_sc_hd__dfxtp_1
X_22784_ _22784_/A _23001_/B _22784_/C vssd1 vssd1 vccd1 vccd1 _22784_/X sky130_fd_sc_hd__and3_1
XFILLER_0_91_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24523_ hold2687/X hold2660/X _24587_/S vssd1 vssd1 vccd1 vccd1 _24524_/A sky130_fd_sc_hd__mux2_1
X_21735_ _21735_/A _21735_/B vssd1 vssd1 vccd1 vccd1 _23056_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_94_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24454_ _24454_/A vssd1 vssd1 vccd1 vccd1 _26215_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21666_ _26337_/Q hold845/X vssd1 vssd1 vccd1 vccd1 _21666_/Y sky130_fd_sc_hd__nand2_1
X_23405_ _23402_/Y _23404_/Y _24946_/A vssd1 vssd1 vccd1 vccd1 _23405_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_188_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20617_ _26292_/Q hold853/X vssd1 vssd1 vccd1 vccd1 _20617_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_145_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24385_ hold2269/X hold1860/X _24433_/S vssd1 vssd1 vccd1 vccd1 _24386_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_163_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21597_ _21597_/A _21597_/B _21597_/C vssd1 vssd1 vccd1 vccd1 _21598_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_85_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26124_ _26216_/CLK _26124_/D vssd1 vssd1 vccd1 vccd1 _26124_/Q sky130_fd_sc_hd__dfxtp_1
X_23336_ _23336_/A _23336_/B hold952/X vssd1 vssd1 vccd1 vccd1 _23342_/A sky130_fd_sc_hd__and3_1
XFILLER_0_116_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20548_ _20551_/A _20551_/C vssd1 vssd1 vccd1 vccd1 _20549_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26055_ _26060_/CLK _26055_/D vssd1 vssd1 vccd1 vccd1 _26055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23267_ _23275_/A _23267_/B vssd1 vssd1 vccd1 vccd1 _23269_/A sky130_fd_sc_hd__nor2_1
X_20479_ _20479_/A _20479_/B vssd1 vssd1 vccd1 vccd1 _20483_/A sky130_fd_sc_hd__nand2_1
X_25006_ _25587_/CLK hold961/X vssd1 vssd1 vccd1 vccd1 hold960/A sky130_fd_sc_hd__dfxtp_1
X_13020_ _12891_/X _14452_/A _12909_/X _25634_/Q vssd1 vssd1 vccd1 vccd1 _13020_/X
+ sky130_fd_sc_hd__a22o_1
X_22218_ _22218_/A _25853_/Q vssd1 vssd1 vccd1 vccd1 _22218_/Y sky130_fd_sc_hd__nand2_1
X_23198_ _23196_/X _23197_/Y _12702_/A vssd1 vssd1 vccd1 vccd1 _25901_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22149_ _25815_/Q _22149_/B vssd1 vssd1 vccd1 vccd1 _22149_/Y sky130_fd_sc_hd__nor2_1
X_14971_ _25421_/Q _14972_/A vssd1 vssd1 vccd1 vccd1 _14973_/A sky130_fd_sc_hd__or2_1
X_16710_ _16712_/B _16712_/A vssd1 vssd1 vccd1 vccd1 _16710_/X sky130_fd_sc_hd__or2_1
XFILLER_0_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25908_ _25913_/CLK _25908_/D vssd1 vssd1 vccd1 vccd1 _25908_/Q sky130_fd_sc_hd__dfxtp_1
X_13922_ _26285_/Q _13801_/X _13793_/X _13921_/Y vssd1 vssd1 vccd1 vccd1 _13923_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17690_ _17723_/A _17690_/B _17690_/C vssd1 vssd1 vccd1 vccd1 _17699_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16641_ _16639_/Y _16641_/B vssd1 vssd1 vccd1 vccd1 _16647_/B sky130_fd_sc_hd__and2b_1
X_25839_ _25860_/CLK _25839_/D vssd1 vssd1 vccd1 vccd1 _25839_/Q sky130_fd_sc_hd__dfxtp_4
X_13853_ _26274_/Q _13801_/X _13793_/X _13852_/Y vssd1 vssd1 vccd1 vccd1 _13854_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12804_ _12726_/B _14322_/A _12752_/X _25593_/Q vssd1 vssd1 vccd1 vccd1 _12804_/X
+ sky130_fd_sc_hd__a22o_1
X_19360_ _20882_/A _21869_/B _25605_/Q vssd1 vssd1 vccd1 vccd1 _20886_/C sky130_fd_sc_hd__nand3_1
X_16572_ _16573_/B _16573_/A vssd1 vssd1 vccd1 vccd1 _16574_/A sky130_fd_sc_hd__nor2_1
X_13784_ _13823_/A _13784_/B vssd1 vssd1 vccd1 vccd1 _13784_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18311_ _18514_/A _18657_/A vssd1 vssd1 vccd1 vccd1 _18312_/B sky130_fd_sc_hd__xnor2_1
X_15523_ _15523_/A _15812_/B vssd1 vssd1 vccd1 vccd1 _15524_/B sky130_fd_sc_hd__nand2_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12735_ _12527_/A _12496_/A _13465_/B vssd1 vssd1 vccd1 vccd1 _14267_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19291_ _20701_/A _19289_/Y _20705_/C vssd1 vssd1 vccd1 vccd1 _19378_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_155_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ _18445_/A _25738_/Q vssd1 vssd1 vccd1 vccd1 _18244_/A sky130_fd_sc_hd__nand2_1
X_12666_ _12666_/A _12671_/C vssd1 vssd1 vccd1 vccd1 _12674_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_167_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15454_ _22866_/B _15454_/B vssd1 vssd1 vccd1 vccd1 _22863_/B sky130_fd_sc_hd__xor2_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14405_ _23245_/A vssd1 vssd1 vccd1 vccd1 _15464_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18173_ _18173_/A _18173_/B _18173_/C vssd1 vssd1 vccd1 vccd1 _21940_/A sky130_fd_sc_hd__nand3_2
X_15385_ _22796_/B _16369_/B _15778_/B vssd1 vssd1 vccd1 vccd1 _16817_/A sky130_fd_sc_hd__nand3_2
X_12597_ _12601_/A _24836_/B _12597_/C vssd1 vssd1 vccd1 vccd1 _12597_/X sky130_fd_sc_hd__and3_1
XFILLER_0_37_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17124_ _17124_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17124_/Y sky130_fd_sc_hd__nand2_1
X_14336_ _14334_/Y hold246/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold247/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold508 hold508/A vssd1 vssd1 vccd1 vccd1 hold508/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold519 hold519/A vssd1 vssd1 vccd1 vccd1 hold519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14267_ _14267_/A _14267_/B _14266_/Y vssd1 vssd1 vccd1 vccd1 _14268_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17055_ _18232_/B _17055_/B vssd1 vssd1 vccd1 vccd1 _17434_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16006_ _16006_/A _16006_/B vssd1 vssd1 vccd1 vccd1 _16014_/A sky130_fd_sc_hd__nand2_1
X_13218_ _18495_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13218_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14198_ _14264_/A _14198_/B vssd1 vssd1 vccd1 vccd1 _14198_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _26161_/Q _13065_/X _13148_/X vssd1 vssd1 vccd1 vccd1 _13149_/X sky130_fd_sc_hd__a21o_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 _16792_/Y vssd1 vssd1 vccd1 vccd1 _25552_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17957_ _18529_/A _17957_/B _18083_/C vssd1 vssd1 vccd1 vccd1 _17958_/C sky130_fd_sc_hd__nand3_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1219 _25752_/Q vssd1 vssd1 vccd1 vccd1 _19723_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16908_ _16906_/Y _16907_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16908_/Y sky130_fd_sc_hd__a21oi_1
X_17888_ _17888_/A _17888_/B vssd1 vssd1 vccd1 vccd1 _22130_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_189_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19627_ _26249_/Q hold665/X vssd1 vssd1 vccd1 vccd1 _19627_/Y sky130_fd_sc_hd__nand2_1
X_16839_ _16837_/Y _15441_/B _16838_/Y vssd1 vssd1 vccd1 vccd1 _16839_/Y sky130_fd_sc_hd__o21ai_1
X_19558_ _19557_/Y _19272_/X _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19559_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_177_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18509_ _18955_/A _18509_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18510_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19489_ _21128_/A _21878_/B _25614_/Q vssd1 vssd1 vccd1 vccd1 _21132_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_158_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21520_ _26328_/Q hold422/X vssd1 vssd1 vccd1 vccd1 _21520_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_180_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21451_ _21451_/A _21451_/B _21451_/C vssd1 vssd1 vccd1 vccd1 _21452_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_127_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20402_ _20405_/A _20405_/C vssd1 vssd1 vccd1 vccd1 _20403_/A sky130_fd_sc_hd__nand2_1
X_24170_ _24170_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24171_/A sky130_fd_sc_hd__and2_1
XFILLER_0_181_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21382_ _21385_/A _21434_/A vssd1 vssd1 vccd1 vccd1 _21384_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_189_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23121_ _23121_/A _23121_/B vssd1 vssd1 vccd1 vccd1 _23122_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20333_ _21499_/A vssd1 vssd1 vccd1 vccd1 _21498_/A sky130_fd_sc_hd__inv_4
XFILLER_0_141_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23052_ _23043_/Y _23051_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _23052_/X sky130_fd_sc_hd__a21o_1
X_20264_ _26283_/Q _20078_/X hold683/X vssd1 vssd1 vccd1 vccd1 _20267_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22003_ _22001_/X _14270_/A _22002_/Y _14777_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _22004_/A sky130_fd_sc_hd__a32o_1
X_20195_ _20195_/A _20195_/B vssd1 vssd1 vccd1 vccd1 _20196_/A sky130_fd_sc_hd__nand2_1
Xhold2410 _26323_/Q vssd1 vssd1 vccd1 vccd1 hold2410/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2421 _24020_/X vssd1 vssd1 vccd1 vccd1 _24021_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2432 _15676_/X vssd1 vssd1 vccd1 vccd1 _15678_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2443 _25468_/Q vssd1 vssd1 vccd1 vccd1 _15680_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2454 _15063_/Y vssd1 vssd1 vccd1 vccd1 _25431_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1720 _21656_/Y vssd1 vssd1 vccd1 vccd1 _25833_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2465 _24394_/X vssd1 vssd1 vccd1 vccd1 _24395_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1731 _17584_/Y vssd1 vssd1 vccd1 vccd1 _25635_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2476 _26306_/Q vssd1 vssd1 vccd1 vccd1 hold2476/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23954_ _23954_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23955_/A sky130_fd_sc_hd__and2_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2487 _26075_/Q vssd1 vssd1 vccd1 vccd1 hold2487/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1742 _25804_/Q vssd1 vssd1 vccd1 vccd1 _21098_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1753 _14977_/Y vssd1 vssd1 vccd1 vccd1 hold1753/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2498 _25660_/Q vssd1 vssd1 vccd1 vccd1 _13158_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1764 _17218_/Y vssd1 vssd1 vccd1 vccd1 _25596_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1775 _25655_/Q vssd1 vssd1 vccd1 vccd1 _18212_/B sky130_fd_sc_hd__buf_2
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22905_ _23058_/A vssd1 vssd1 vccd1 vccd1 _22906_/A sky130_fd_sc_hd__inv_2
X_23885_ _23885_/A vssd1 vssd1 vccd1 vccd1 _26032_/D sky130_fd_sc_hd__clkbuf_1
Xhold1786 _17191_/Y vssd1 vssd1 vccd1 vccd1 _25594_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1797 _22588_/Y vssd1 vssd1 vccd1 vccd1 _25867_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22836_ _22836_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _22836_/Y sky130_fd_sc_hd__nand2_1
X_25624_ _26130_/CLK _25624_/D vssd1 vssd1 vccd1 vccd1 _25624_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_168_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22767_ _22766_/A _22454_/X _22766_/B vssd1 vssd1 vccd1 vccd1 _22768_/C sky130_fd_sc_hd__o21ai_1
X_25555_ _25878_/CLK _25555_/D vssd1 vssd1 vccd1 vccd1 _25555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _23193_/B vssd1 vssd1 vccd1 vccd1 _13465_/B sky130_fd_sc_hd__inv_2
X_24506_ _24506_/A vssd1 vssd1 vccd1 vccd1 _26232_/D sky130_fd_sc_hd__clkbuf_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21718_ _21718_/A _22902_/B vssd1 vssd1 vccd1 vccd1 _21718_/Y sky130_fd_sc_hd__nand2_1
X_25486_ _25939_/CLK hold811/X vssd1 vssd1 vccd1 vccd1 hold809/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22698_ _22698_/A _22698_/B vssd1 vssd1 vccd1 vccd1 _23168_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24437_ hold1987/X hold1938/X _24510_/S vssd1 vssd1 vccd1 vccd1 _24438_/A sky130_fd_sc_hd__mux2_1
X_21649_ _26336_/Q _19130_/X hold632/X vssd1 vssd1 vccd1 vccd1 _21652_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_164_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15170_ _16736_/B vssd1 vssd1 vccd1 vccd1 _22529_/B sky130_fd_sc_hd__inv_2
XFILLER_0_105_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24368_ _24368_/A vssd1 vssd1 vccd1 vccd1 _26187_/D sky130_fd_sc_hd__clkbuf_1
X_14121_ _18490_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14121_/Y sky130_fd_sc_hd__nor2_1
X_23319_ _23324_/A vssd1 vssd1 vccd1 vccd1 _23321_/A sky130_fd_sc_hd__inv_2
XFILLER_0_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26107_ _26231_/CLK _26107_/D vssd1 vssd1 vccd1 vccd1 _26107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24299_ hold2077/X _26165_/Q _24356_/S vssd1 vssd1 vccd1 vccd1 _24299_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_132_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14052_ _25803_/Q vssd1 vssd1 vccd1 vccd1 _18264_/B sky130_fd_sc_hd__inv_2
X_26038_ _26040_/CLK _26038_/D vssd1 vssd1 vccd1 vccd1 _26038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13003_ _12891_/X _14443_/A _12909_/X _25631_/Q vssd1 vssd1 vccd1 vccd1 _13003_/X
+ sky130_fd_sc_hd__a22o_1
X_18860_ _18858_/X _18269_/X _18859_/X vssd1 vssd1 vccd1 vccd1 _18861_/A sky130_fd_sc_hd__a21o_1
X_17811_ _17811_/A _25791_/Q _17811_/C vssd1 vssd1 vccd1 vccd1 _20668_/B sky130_fd_sc_hd__nand3_1
X_18791_ _18791_/A _25829_/Q _18791_/C vssd1 vssd1 vccd1 vccd1 _20643_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17742_ _17742_/A _20957_/A vssd1 vssd1 vccd1 vccd1 _17773_/B sky130_fd_sc_hd__nand2_2
X_14954_ _14955_/B _14955_/A vssd1 vssd1 vccd1 vccd1 _14956_/A sky130_fd_sc_hd__or2_1
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13905_ hold612/X _13904_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold613/A sky130_fd_sc_hd__a21oi_1
X_17673_ _17688_/A _17707_/B vssd1 vssd1 vccd1 vccd1 _17719_/B sky130_fd_sc_hd__nand2_2
X_14885_ _14891_/B _22366_/A vssd1 vssd1 vccd1 vccd1 _22365_/B sky130_fd_sc_hd__xnor2_2
Xclkbuf_leaf_195_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _26116_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19412_ _26234_/Q _12537_/B hold563/X vssd1 vssd1 vccd1 vccd1 _19412_/Y sky130_fd_sc_hd__a21oi_1
X_16624_ hold948/X vssd1 vssd1 vccd1 vccd1 _16627_/B sky130_fd_sc_hd__inv_2
XFILLER_0_159_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13836_ _13941_/A _13836_/B vssd1 vssd1 vccd1 vccd1 _13836_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_186_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19343_ _19342_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19344_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16555_ _16555_/A _16555_/B vssd1 vssd1 vccd1 vccd1 _16564_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13767_ _14125_/A vssd1 vssd1 vccd1 vccd1 _13880_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_134_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15506_ _16865_/B vssd1 vssd1 vccd1 vccd1 _22914_/B sky130_fd_sc_hd__inv_2
XFILLER_0_85_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12718_ _12718_/A hold410/X vssd1 vssd1 vccd1 vccd1 hold411/A sky130_fd_sc_hd__nand2_1
X_19274_ _19270_/Y _19274_/B _19980_/B vssd1 vssd1 vccd1 vccd1 _19274_/X sky130_fd_sc_hd__and3b_1
X_16486_ _16492_/B _16486_/B vssd1 vssd1 vccd1 vccd1 _16487_/B sky130_fd_sc_hd__nor2_1
X_13698_ hold666/X _13697_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold667/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18225_ _21002_/B _22008_/A vssd1 vssd1 vccd1 vccd1 _20993_/A sky130_fd_sc_hd__nand2_2
X_15437_ _15621_/A _16411_/B vssd1 vssd1 vccd1 vccd1 _15440_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_127_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12649_ _12712_/A _12711_/D vssd1 vssd1 vccd1 vccd1 _12651_/A sky130_fd_sc_hd__and2_1
XFILLER_0_72_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18156_ _18529_/A _18156_/B hold922/A vssd1 vssd1 vccd1 vccd1 _18159_/B sky130_fd_sc_hd__nand3_1
X_15368_ _22779_/B _15812_/B vssd1 vssd1 vccd1 vccd1 _15369_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_124_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17107_ _17456_/A _17534_/A vssd1 vssd1 vccd1 vccd1 _17108_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14319_ _14319_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14319_/Y sky130_fd_sc_hd__nand2_1
Xhold305 hold305/A vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18087_ _18087_/A _18087_/B _18087_/C vssd1 vssd1 vccd1 vccd1 _22250_/A sky130_fd_sc_hd__nand3_2
Xhold316 hold316/A vssd1 vssd1 vccd1 vccd1 hold316/X sky130_fd_sc_hd__dlygate4sd3_1
X_15299_ _15299_/A _15810_/B vssd1 vssd1 vccd1 vccd1 _15300_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_111_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold327 hold327/A vssd1 vssd1 vccd1 vccd1 hold327/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 hold338/A vssd1 vssd1 vccd1 vccd1 hold338/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold349 hold349/A vssd1 vssd1 vccd1 vccd1 hold349/X sky130_fd_sc_hd__dlygate4sd3_1
X_17038_ _20350_/B _25847_/Q _25783_/Q vssd1 vssd1 vccd1 vccd1 _17039_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_180_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ _19039_/A _18989_/B vssd1 vssd1 vccd1 vccd1 _18989_/X sky130_fd_sc_hd__xor2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 _25523_/Q vssd1 vssd1 vccd1 vccd1 _16483_/B sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1016 _13076_/X vssd1 vssd1 vccd1 vccd1 _25064_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1027 _25054_/Q vssd1 vssd1 vccd1 vccd1 _17572_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1038 _12924_/X vssd1 vssd1 vccd1 vccd1 _25035_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 _25129_/Q vssd1 vssd1 vccd1 vccd1 _19082_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20951_ _21451_/B _21497_/C vssd1 vssd1 vccd1 vccd1 _20952_/C sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_186_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _25748_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_178_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23670_ _23670_/A vssd1 vssd1 vccd1 vccd1 _25962_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20882_ _20882_/A _21869_/B vssd1 vssd1 vccd1 vccd1 _20883_/A sky130_fd_sc_hd__nand2_1
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22621_ _22621_/A _22621_/B vssd1 vssd1 vccd1 vccd1 _23120_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_113_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25340_ _26298_/CLK hold97/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__dfxtp_1
X_22552_ _22653_/A _22552_/B vssd1 vssd1 vccd1 vccd1 _22552_/X sky130_fd_sc_hd__or2_1
XFILLER_0_119_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21503_ _26327_/Q _21228_/X hold823/X vssd1 vssd1 vccd1 vccd1 _21506_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_173_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25271_ _26103_/CLK hold190/X vssd1 vssd1 vccd1 vccd1 hold188/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22483_ _22483_/A _22900_/B vssd1 vssd1 vccd1 vccd1 _22483_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24222_ hold1961/X _26140_/Q _24279_/S vssd1 vssd1 vccd1 vccd1 _24222_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21434_ _21434_/A _21482_/A vssd1 vssd1 vccd1 vccd1 _21435_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_133_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24153_ _24153_/A vssd1 vssd1 vccd1 vccd1 _26117_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21365_ _21369_/A _21418_/A vssd1 vssd1 vccd1 vccd1 _21368_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_110_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _25992_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_102_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23104_ _23104_/A _23104_/B vssd1 vssd1 vccd1 vccd1 _23105_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20316_ _20316_/A _20317_/A vssd1 vssd1 vccd1 vccd1 _20319_/A sky130_fd_sc_hd__nand2_1
X_24084_ _24084_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24085_/A sky130_fd_sc_hd__and2_1
XFILLER_0_101_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold850 hold850/A vssd1 vssd1 vccd1 vccd1 hold850/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21296_ _21296_/A _21296_/B vssd1 vssd1 vccd1 vccd1 _21298_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold861 hold861/A vssd1 vssd1 vccd1 vccd1 hold861/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 hold872/A vssd1 vssd1 vccd1 vccd1 hold872/X sky130_fd_sc_hd__dlygate4sd3_1
X_23035_ _23035_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _23035_/Y sky130_fd_sc_hd__nand2_1
Xhold883 hold883/A vssd1 vssd1 vccd1 vccd1 hold883/X sky130_fd_sc_hd__buf_1
X_20247_ _20247_/A _21958_/A vssd1 vssd1 vccd1 vccd1 _20248_/A sky130_fd_sc_hd__nand2_1
Xhold894 hold894/A vssd1 vssd1 vccd1 vccd1 hold894/X sky130_fd_sc_hd__dlygate4sd3_1
X_20178_ _20178_/A vssd1 vssd1 vccd1 vccd1 _20180_/B sky130_fd_sc_hd__inv_2
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2240 _26029_/Q vssd1 vssd1 vccd1 vccd1 hold2240/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2251 _25962_/Q vssd1 vssd1 vccd1 vccd1 hold2251/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2262 _12630_/X vssd1 vssd1 vccd1 vccd1 _12631_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2273 _12597_/X vssd1 vssd1 vccd1 vccd1 _12598_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24986_ _24990_/CLK _24986_/D vssd1 vssd1 vccd1 vccd1 _24986_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2284 _26115_/Q vssd1 vssd1 vccd1 vccd1 hold2284/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1550 _13400_/X vssd1 vssd1 vccd1 vccd1 _25118_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2295 _24391_/X vssd1 vssd1 vccd1 vccd1 _24392_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1561 _25639_/Q vssd1 vssd1 vccd1 vccd1 _17613_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23937_ _23937_/A vssd1 vssd1 vccd1 vccd1 _26047_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_177_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _26239_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1572 _25582_/Q vssd1 vssd1 vccd1 vccd1 _17016_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1583 _17439_/Y vssd1 vssd1 vccd1 vccd1 _25615_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1594 _25259_/Q vssd1 vssd1 vccd1 vccd1 _12482_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14670_ _14688_/A hold62/X vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23868_ hold2043/X _26027_/Q _23907_/S vssd1 vssd1 vccd1 vccd1 _23868_/X sky130_fd_sc_hd__mux2_1
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25607_ _26240_/CLK _25607_/D vssd1 vssd1 vccd1 vccd1 _25607_/Q sky130_fd_sc_hd__dfxtp_2
X_13621_ _26237_/Q _13612_/X _13605_/X _13620_/Y vssd1 vssd1 vccd1 vccd1 _13622_/B
+ sky130_fd_sc_hd__a22o_1
X_22819_ _22819_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _22819_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23799_ _23799_/A vssd1 vssd1 vccd1 vccd1 _26004_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16340_ _16340_/A _16361_/A vssd1 vssd1 vccd1 vccd1 _16341_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_183_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25538_ _25539_/CLK hold610/X vssd1 vssd1 vccd1 vccd1 hold608/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13552_ _13583_/A _13552_/B vssd1 vssd1 vccd1 vccd1 _13552_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12503_ _12503_/A vssd1 vssd1 vccd1 vccd1 _23923_/A sky130_fd_sc_hd__inv_1
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16271_ _16276_/B _16271_/B vssd1 vssd1 vccd1 vccd1 _16272_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_152_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13483_ _26215_/Q _13426_/X _13468_/X _13482_/Y vssd1 vssd1 vccd1 vccd1 _13484_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25469_ _26012_/CLK _25469_/D vssd1 vssd1 vccd1 vccd1 _25469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18010_ _18010_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _18010_/Y sky130_fd_sc_hd__nand2_1
X_15222_ _16757_/B vssd1 vssd1 vccd1 vccd1 _22606_/B sky130_fd_sc_hd__inv_2
XFILLER_0_180_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15153_ _15153_/A _15776_/B vssd1 vssd1 vccd1 vccd1 _15154_/B sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_101_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _25933_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_164_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14104_ _14180_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14104_/Y sky130_fd_sc_hd__nand2_1
X_15084_ _15084_/A _15084_/B vssd1 vssd1 vccd1 vccd1 _15106_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19961_ _19961_/A _19961_/B vssd1 vssd1 vccd1 vccd1 _19961_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14035_ _26303_/Q _13988_/X _13981_/X _14034_/Y vssd1 vssd1 vccd1 vccd1 _14036_/B
+ sky130_fd_sc_hd__a22o_1
X_18912_ _18912_/A _25835_/Q _18912_/C vssd1 vssd1 vccd1 vccd1 _20006_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19892_ _19890_/Y _19891_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19892_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18843_ _18841_/Y _18842_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25686_/D sky130_fd_sc_hd__a21oi_1
X_18774_ _18774_/A _18774_/B _18774_/C vssd1 vssd1 vccd1 vccd1 _22490_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_98_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15986_ _15986_/A _15986_/B vssd1 vssd1 vccd1 vccd1 _15999_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17725_ _17725_/A _17725_/B _17725_/C vssd1 vssd1 vccd1 vccd1 _17728_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_171_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14937_ _14938_/B _14938_/A vssd1 vssd1 vccd1 vccd1 _14939_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_168_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _25794_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_145_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17656_ _18252_/A _17656_/B vssd1 vssd1 vccd1 vccd1 _17656_/Y sky130_fd_sc_hd__nand2_1
X_14868_ _22322_/B _15543_/B vssd1 vssd1 vccd1 vccd1 _14869_/A sky130_fd_sc_hd__nand2_1
X_16607_ _16607_/A vssd1 vssd1 vccd1 vccd1 _16629_/B sky130_fd_sc_hd__inv_2
XFILLER_0_175_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13819_ _13880_/A hold803/X vssd1 vssd1 vccd1 vccd1 hold804/A sky130_fd_sc_hd__nand2_1
X_17587_ _17624_/A _17587_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _17587_/X sky130_fd_sc_hd__and3_1
X_14799_ _22090_/B _15778_/B vssd1 vssd1 vccd1 vccd1 _14800_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19326_ _19324_/Y _19325_/Y _19086_/X vssd1 vssd1 vccd1 vccd1 _19326_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16538_ _16536_/X _16537_/Y _16231_/A vssd1 vssd1 vccd1 vccd1 _16538_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_161_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19257_ _19257_/A _20625_/B vssd1 vssd1 vccd1 vccd1 _19257_/Y sky130_fd_sc_hd__nor2_1
X_16469_ _16486_/B vssd1 vssd1 vccd1 vccd1 _16470_/B sky130_fd_sc_hd__inv_2
XFILLER_0_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18208_ _18535_/A _18208_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _18208_/X sky130_fd_sc_hd__and3_1
X_19188_ _20428_/A _22106_/A _25593_/Q vssd1 vssd1 vccd1 vccd1 _20432_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_182_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18139_ _18139_/A _18139_/B _18139_/C vssd1 vssd1 vccd1 vccd1 _21906_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_5_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold102 hold102/A vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 hold113/A vssd1 vssd1 vccd1 vccd1 hold113/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold124 hold124/A vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold135 hold135/A vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
X_21150_ _21636_/A _21150_/B _21149_/X vssd1 vssd1 vccd1 vccd1 _21151_/B sky130_fd_sc_hd__or3b_1
Xhold146 hold146/A vssd1 vssd1 vccd1 vccd1 hold146/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold157 hold157/A vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 hold168/A vssd1 vssd1 vccd1 vccd1 hold168/X sky130_fd_sc_hd__dlygate4sd3_1
X_20101_ _20101_/A _25879_/Q vssd1 vssd1 vccd1 vccd1 _20106_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold179 hold179/A vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__dlygate4sd3_1
X_21081_ _21080_/B _21081_/B _21081_/C vssd1 vssd1 vccd1 vccd1 _21082_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_186_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20032_ _20032_/A _20032_/B vssd1 vssd1 vccd1 vccd1 _20034_/A sky130_fd_sc_hd__nand2_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24840_ _24838_/X _24839_/X _24858_/S vssd1 vssd1 vccd1 vccd1 _24840_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_119_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_159_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _26297_/CLK sky130_fd_sc_hd__clkbuf_16
X_21983_ _21983_/A _21983_/B vssd1 vssd1 vccd1 vccd1 _21983_/Y sky130_fd_sc_hd__nand2_1
X_24771_ _24771_/A vssd1 vssd1 vccd1 vccd1 _26318_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23722_ _23722_/A vssd1 vssd1 vccd1 vccd1 _25979_/D sky130_fd_sc_hd__clkbuf_1
X_20934_ _20932_/Y _20933_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _20934_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23653_ hold2133/X hold2092/X _23677_/S vssd1 vssd1 vccd1 vccd1 _23654_/A sky130_fd_sc_hd__mux2_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20865_ _21451_/B vssd1 vssd1 vccd1 vccd1 _21448_/C sky130_fd_sc_hd__inv_2
XFILLER_0_77_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22604_ _15225_/B _22387_/B _14273_/X vssd1 vssd1 vccd1 vccd1 _22604_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23584_ hold476/X _25938_/Q _25937_/Q _25936_/Q vssd1 vssd1 vccd1 vccd1 _23586_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_0_119_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20796_ _20798_/B _20798_/C vssd1 vssd1 vccd1 vccd1 _20797_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22535_ _22525_/Y _22533_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22535_/X sky130_fd_sc_hd__a21o_1
X_25323_ _26148_/CLK hold313/X vssd1 vssd1 vccd1 vccd1 hold311/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25254_ _25864_/CLK hold846/X vssd1 vssd1 vccd1 vccd1 hold845/A sky130_fd_sc_hd__dfxtp_1
X_22466_ _19788_/A _22465_/A _22465_/Y vssd1 vssd1 vccd1 vccd1 _22468_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_106_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24205_ _24205_/A vssd1 vssd1 vccd1 vccd1 _26134_/D sky130_fd_sc_hd__clkbuf_1
X_21417_ _21417_/A _21465_/A vssd1 vssd1 vccd1 vccd1 _21419_/A sky130_fd_sc_hd__nand2_1
X_25185_ _26269_/CLK hold679/X vssd1 vssd1 vccd1 vccd1 hold677/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22397_ _22397_/A _22397_/B vssd1 vssd1 vccd1 vccd1 _22975_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_103_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24136_ hold2135/X hold1972/X _24203_/S vssd1 vssd1 vccd1 vccd1 _24137_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21348_ _21346_/Y _21347_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21348_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24067_ _24067_/A vssd1 vssd1 vccd1 vccd1 _26089_/D sky130_fd_sc_hd__clkbuf_1
X_21279_ _21279_/A _21279_/B _21279_/C vssd1 vssd1 vccd1 vccd1 _21280_/B sky130_fd_sc_hd__nand3_1
Xhold680 hold680/A vssd1 vssd1 vccd1 vccd1 hold680/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold691 hold691/A vssd1 vssd1 vccd1 vccd1 hold691/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23018_ hold1551/X _22421_/X _23012_/X _23013_/Y _23017_/X vssd1 vssd1 vccd1 vccd1
+ _23018_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_60_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ _15840_/A vssd1 vssd1 vccd1 vccd1 _16676_/A sky130_fd_sc_hd__buf_12
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2070 _26021_/Q vssd1 vssd1 vccd1 vccd1 hold2070/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2081 _23892_/X vssd1 vssd1 vccd1 vccd1 _23893_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2092 _25957_/Q vssd1 vssd1 vccd1 vccd1 hold2092/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _25473_/Q vssd1 vssd1 vccd1 vccd1 _15780_/B sky130_fd_sc_hd__inv_2
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24969_ _25378_/CLK _24969_/D vssd1 vssd1 vccd1 vccd1 _24969_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ _12891_/X _14431_/A _12909_/X _25627_/Q vssd1 vssd1 vccd1 vccd1 _12983_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1380 _20545_/Y vssd1 vssd1 vccd1 vccd1 _25787_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17510_ _17605_/A _17510_/B vssd1 vssd1 vccd1 vccd1 _17510_/Y sky130_fd_sc_hd__nand2_1
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14722_ _14720_/Y _14721_/Y _14646_/X vssd1 vssd1 vccd1 vccd1 _14722_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1391 _25123_/Q vssd1 vssd1 vccd1 vccd1 _19040_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18490_ _18490_/A _18490_/B _18490_/C vssd1 vssd1 vccd1 vccd1 _22122_/A sky130_fd_sc_hd__nand3_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _17441_/A _17441_/B vssd1 vssd1 vccd1 vccd1 _17441_/X sky130_fd_sc_hd__xor2_1
X_14653_ _14651_/Y hold174/X _14646_/X vssd1 vssd1 vccd1 vccd1 hold175/A sky130_fd_sc_hd__a21oi_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _13642_/A hold641/X vssd1 vssd1 vccd1 vccd1 hold642/A sky130_fd_sc_hd__nand2_1
X_17372_ _17638_/A _17372_/B vssd1 vssd1 vccd1 vccd1 _17372_/X sky130_fd_sc_hd__xor2_1
X_14584_ _14584_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14584_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_83_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19111_ _19111_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _19111_/Y sky130_fd_sc_hd__nand2_1
X_16323_ _16336_/B _16324_/A vssd1 vssd1 vccd1 vccd1 _16323_/X sky130_fd_sc_hd__or2_1
XFILLER_0_172_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13535_ hold510/X _13534_/Y _12558_/B vssd1 vssd1 vccd1 vccd1 hold511/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19042_ _19042_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _19042_/Y sky130_fd_sc_hd__nand2_1
X_16254_ _16254_/A _16254_/B vssd1 vssd1 vccd1 vccd1 _16264_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_153_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13466_ _13466_/A _17008_/B vssd1 vssd1 vccd1 vccd1 _13467_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_125_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15205_ _16750_/B vssd1 vssd1 vccd1 vccd1 _22580_/B sky130_fd_sc_hd__inv_2
XFILLER_0_51_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16185_ _16183_/X _16184_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _16185_/X sky130_fd_sc_hd__a21o_1
X_13397_ _13220_/X _14654_/A _13242_/X _19774_/A vssd1 vssd1 vccd1 vccd1 _13397_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15136_ _15774_/B vssd1 vssd1 vccd1 vccd1 _15776_/B sky130_fd_sc_hd__buf_8
XFILLER_0_121_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15067_ _15067_/A _15067_/B vssd1 vssd1 vccd1 vccd1 _15067_/X sky130_fd_sc_hd__or2_1
X_19944_ _26272_/Q hold812/X vssd1 vssd1 vccd1 vccd1 _19944_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_120_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14018_ _14061_/A _14018_/B vssd1 vssd1 vccd1 vccd1 _14018_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_103_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19875_ _19875_/A _19875_/B vssd1 vssd1 vccd1 vccd1 _19875_/Y sky130_fd_sc_hd__nand2_1
X_18826_ _20712_/B _19844_/A vssd1 vssd1 vccd1 vccd1 _18827_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18757_ _18960_/A _19010_/A vssd1 vssd1 vccd1 vccd1 _18758_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15969_ _22060_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _15971_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17708_ _17708_/A _17750_/B vssd1 vssd1 vccd1 vccd1 _17709_/C sky130_fd_sc_hd__nand2_1
X_18688_ _25888_/Q _22390_/A vssd1 vssd1 vccd1 vccd1 _18696_/A sky130_fd_sc_hd__or2_2
XFILLER_0_187_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17639_ _18535_/A _17639_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _17639_/X sky130_fd_sc_hd__and3_1
XFILLER_0_176_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20650_ _21351_/C _21629_/B vssd1 vssd1 vccd1 vccd1 _20651_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_176_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19309_ _19307_/X _19308_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19309_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20581_ _20581_/A _20581_/B vssd1 vssd1 vccd1 vccd1 _20582_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_144_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22320_ _22561_/A _22320_/B vssd1 vssd1 vccd1 vccd1 _22320_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_144_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22251_ _19257_/A _22250_/A _22250_/Y vssd1 vssd1 vccd1 vccd1 _22253_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21202_ _26311_/Q hold789/X vssd1 vssd1 vccd1 vccd1 _21202_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_103_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22182_ _19630_/A _22181_/A _22181_/Y vssd1 vssd1 vccd1 vccd1 _22184_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_112_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21133_ _21136_/A _21136_/B vssd1 vssd1 vccd1 vccd1 _21135_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25941_ _26040_/CLK _25941_/D vssd1 vssd1 vccd1 vccd1 _25941_/Q sky130_fd_sc_hd__dfxtp_1
X_21064_ _21064_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _21070_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20015_ _20018_/A _20018_/B vssd1 vssd1 vccd1 vccd1 _20017_/A sky130_fd_sc_hd__nand2_1
X_25872_ _25883_/CLK _25872_/D vssd1 vssd1 vccd1 vccd1 _25872_/Q sky130_fd_sc_hd__dfxtp_2
X_24823_ hold2659/X hold2366/X _24835_/S vssd1 vssd1 vccd1 vccd1 _24824_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24754_ hold2746/X hold2730/X _24817_/S vssd1 vssd1 vccd1 vccd1 _24755_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_96_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21966_ _21964_/Y _21965_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _21966_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23705_ hold2128/X hold1957/X _23754_/S vssd1 vssd1 vccd1 vccd1 _23706_/A sky130_fd_sc_hd__mux2_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20917_ _20917_/A _20917_/B vssd1 vssd1 vccd1 vccd1 _21483_/B sky130_fd_sc_hd__nand2_4
X_21897_ _23245_/A vssd1 vssd1 vccd1 vccd1 _21897_/X sky130_fd_sc_hd__clkbuf_8
X_24685_ _24685_/A vssd1 vssd1 vccd1 vccd1 _26290_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23636_ _23636_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23637_/A sky130_fd_sc_hd__and2_1
X_20848_ _26298_/Q hold554/X vssd1 vssd1 vccd1 vccd1 _20848_/Y sky130_fd_sc_hd__nand2_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23567_ hold62/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23567_/X sky130_fd_sc_hd__or2b_1
X_20779_ _20779_/A _21764_/B vssd1 vssd1 vccd1 vccd1 _20780_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25306_ _25636_/CLK hold172/X vssd1 vssd1 vccd1 vccd1 hold170/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13320_ _18819_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13320_/X sky130_fd_sc_hd__or2_1
X_22518_ _22518_/A _22518_/B vssd1 vssd1 vccd1 vccd1 _22519_/B sky130_fd_sc_hd__nand2_1
X_26286_ _26286_/CLK _26286_/D vssd1 vssd1 vccd1 vccd1 _26286_/Q sky130_fd_sc_hd__dfxtp_2
X_23498_ _24940_/S hold179/A _23497_/X vssd1 vssd1 vccd1 vccd1 _23498_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22449_ _22653_/A _22449_/B vssd1 vssd1 vccd1 vccd1 _22449_/X sky130_fd_sc_hd__or2_1
X_13251_ _18597_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13251_/X sky130_fd_sc_hd__or2_1
X_25237_ _25817_/CLK hold750/X vssd1 vssd1 vccd1 vccd1 hold748/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13182_ _13182_/A vssd1 vssd1 vccd1 vccd1 _19289_/A sky130_fd_sc_hd__buf_4
XFILLER_0_60_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25168_ _25752_/CLK hold379/X vssd1 vssd1 vccd1 vccd1 hold377/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24119_ _24119_/A vssd1 vssd1 vccd1 vccd1 _26106_/D sky130_fd_sc_hd__clkbuf_1
X_17990_ _17990_/A _17990_/B _17990_/C vssd1 vssd1 vccd1 vccd1 _22192_/A sky130_fd_sc_hd__nand3_2
X_25099_ _26184_/CLK _25099_/D vssd1 vssd1 vccd1 vccd1 _25099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16941_ _17568_/A vssd1 vssd1 vccd1 vccd1 _16941_/X sky130_fd_sc_hd__buf_8
X_19660_ _20199_/A _22237_/B _25626_/Q vssd1 vssd1 vccd1 vccd1 _20204_/C sky130_fd_sc_hd__nand3_1
X_16872_ _16977_/A _16872_/B vssd1 vssd1 vccd1 vccd1 _16872_/Y sky130_fd_sc_hd__nand2_1
X_18611_ _18611_/A _25756_/Q vssd1 vssd1 vccd1 vccd1 _18613_/A sky130_fd_sc_hd__nand2_1
X_15823_ _15823_/A _15830_/B _15830_/A vssd1 vssd1 vccd1 vccd1 _15824_/A sky130_fd_sc_hd__and3_1
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19591_ _19607_/B _19678_/B vssd1 vssd1 vccd1 vccd1 _19593_/A sky130_fd_sc_hd__xnor2_1
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18542_ _22208_/B _25625_/Q vssd1 vssd1 vccd1 vccd1 _18544_/A sky130_fd_sc_hd__nand2_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _26041_/Q _25977_/Q _15773_/S vssd1 vssd1 vccd1 vccd1 _15755_/A sky130_fd_sc_hd__mux2_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12966_ _26255_/Q _25624_/Q vssd1 vssd1 vccd1 vccd1 _14422_/A sky130_fd_sc_hd__xor2_1
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _15839_/A _14705_/B vssd1 vssd1 vccd1 vccd1 _21760_/A sky130_fd_sc_hd__nand2_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18473_ _18678_/A _18818_/A vssd1 vssd1 vccd1 vccd1 _18474_/B sky130_fd_sc_hd__xnor2_1
X_15685_ _23076_/B _15776_/B vssd1 vssd1 vccd1 vccd1 _15686_/A sky130_fd_sc_hd__nand2_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _26242_/Q _25611_/Q vssd1 vssd1 vccd1 vccd1 _14379_/A sky130_fd_sc_hd__xor2_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17424_ _17624_/A _17424_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17424_/X sky130_fd_sc_hd__and3_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _14645_/A hold449/X vssd1 vssd1 vccd1 vccd1 hold450/A sky130_fd_sc_hd__nand2_1
XFILLER_0_185_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _17355_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17355_/Y sky130_fd_sc_hd__nand2_1
X_14567_ _14585_/A hold305/X vssd1 vssd1 vccd1 vccd1 hold306/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16306_ _16306_/A _16306_/B vssd1 vssd1 vccd1 vccd1 _16307_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13518_ _18155_/B _13518_/B vssd1 vssd1 vccd1 vccd1 _13518_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_153_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17286_ _17467_/A _17286_/B vssd1 vssd1 vccd1 vccd1 _17286_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14498_ _14525_/A hold248/X vssd1 vssd1 vccd1 vccd1 hold249/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19025_ _19025_/A _19025_/B vssd1 vssd1 vccd1 vccd1 _19025_/X sky130_fd_sc_hd__xor2_1
X_16237_ _16237_/A vssd1 vssd1 vccd1 vccd1 _16245_/A sky130_fd_sc_hd__inv_2
X_13449_ _13220_/A _14681_/A _13242_/A _25707_/Q vssd1 vssd1 vccd1 vccd1 _13449_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_180_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16168_ _16168_/A _16168_/B vssd1 vssd1 vccd1 vccd1 _16169_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15119_ _15621_/A _16165_/B vssd1 vssd1 vccd1 vccd1 _15122_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_121_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16099_ _16099_/A _16103_/B vssd1 vssd1 vccd1 vccd1 _16099_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_11_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19927_ _19928_/B _19928_/A vssd1 vssd1 vccd1 vccd1 _19927_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19858_ _20751_/A _22590_/B _25640_/Q vssd1 vssd1 vccd1 vccd1 _20756_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_78_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18809_ _18951_/A _18813_/B vssd1 vssd1 vccd1 vccd1 _18811_/A sky130_fd_sc_hd__nand2_1
X_19789_ _20557_/A _22463_/B _25635_/Q vssd1 vssd1 vccd1 vccd1 _20562_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21820_ _25840_/Q _25776_/Q vssd1 vssd1 vccd1 vccd1 _21821_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_92_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21751_ _21751_/A _21751_/B vssd1 vssd1 vccd1 vccd1 _22891_/A sky130_fd_sc_hd__xor2_4
Xclkbuf_leaf_90_clk clkbuf_leaf_95_clk/A vssd1 vssd1 vccd1 vccd1 _25501_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20702_ _20702_/A _20702_/B vssd1 vssd1 vccd1 vccd1 _20705_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24470_ _24470_/A vssd1 vssd1 vccd1 vccd1 _26220_/D sky130_fd_sc_hd__clkbuf_1
X_21682_ _26338_/Q hold650/X vssd1 vssd1 vccd1 vccd1 _21682_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23421_ _24940_/S hold164/A _23420_/X vssd1 vssd1 vccd1 vccd1 _23421_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_4_9__f_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_9__f_clk/X
+ sky130_fd_sc_hd__clkbuf_16
X_20633_ _21351_/C vssd1 vssd1 vccd1 vccd1 _21354_/B sky130_fd_sc_hd__inv_2
XFILLER_0_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23352_ _23352_/A _23377_/B _23356_/A vssd1 vssd1 vccd1 vccd1 _23352_/X sky130_fd_sc_hd__and3_1
XFILLER_0_34_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26140_ _26142_/CLK _26140_/D vssd1 vssd1 vccd1 vccd1 _26140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20564_ _20566_/B vssd1 vssd1 vccd1 vccd1 _20565_/B sky130_fd_sc_hd__inv_2
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22303_ _22303_/A _22303_/B vssd1 vssd1 vccd1 vccd1 _22907_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23283_ _23281_/X hold833/X _12702_/A vssd1 vssd1 vccd1 vccd1 hold834/A sky130_fd_sc_hd__a21oi_1
X_26071_ _26073_/CLK _26071_/D vssd1 vssd1 vccd1 vccd1 _26071_/Q sky130_fd_sc_hd__dfxtp_1
X_20495_ _20495_/A _21198_/B _20495_/C vssd1 vssd1 vccd1 vccd1 _20496_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_171_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22234_ _22232_/X _15839_/B _22233_/Y _14844_/A _21725_/X vssd1 vssd1 vccd1 vccd1
+ _22235_/A sky130_fd_sc_hd__a32o_1
X_25022_ _26231_/CLK _25022_/D vssd1 vssd1 vccd1 vccd1 _25022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22165_ _22165_/A _22165_/B vssd1 vssd1 vccd1 vccd1 _22166_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21116_ _21548_/B _21594_/C vssd1 vssd1 vccd1 vccd1 _21117_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_160_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22096_ _18472_/A _25813_/Q _22094_/Y _22095_/Y vssd1 vssd1 vccd1 vccd1 _22097_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_121_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25924_ _25925_/CLK _25924_/D vssd1 vssd1 vccd1 vccd1 _25924_/Q sky130_fd_sc_hd__dfxtp_1
X_21047_ _21047_/A _21773_/B vssd1 vssd1 vccd1 vccd1 _21048_/A sky130_fd_sc_hd__nand2_1
X_25855_ _26339_/CLK _25855_/D vssd1 vssd1 vccd1 vccd1 _25855_/Q sky130_fd_sc_hd__dfxtp_4
X_24806_ _24806_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24807_/A sky130_fd_sc_hd__and2_1
X_12820_ _26099_/Q _12748_/X _12819_/X vssd1 vssd1 vccd1 vccd1 _12820_/X sky130_fd_sc_hd__a21o_1
X_25786_ _26287_/CLK _25786_/D vssd1 vssd1 vccd1 vccd1 _25786_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_97_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22998_ _26072_/Q vssd1 vssd1 vccd1 vccd1 _22999_/A sky130_fd_sc_hd__inv_2
XFILLER_0_16_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _12751_/A vssd1 vssd1 vccd1 vccd1 _13242_/A sky130_fd_sc_hd__buf_8
XFILLER_0_16_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24737_ hold2745/X hold2648/X _24740_/S vssd1 vssd1 vccd1 vccd1 _24738_/A sky130_fd_sc_hd__mux2_1
X_21949_ _21949_/A _21949_/B vssd1 vssd1 vccd1 vccd1 _21949_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_179_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_81_clk clkbuf_leaf_82_clk/A vssd1 vssd1 vccd1 vccd1 _25859_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _15414_/A _15552_/A _15469_/Y vssd1 vssd1 vccd1 vccd1 _15470_/X sky130_fd_sc_hd__a21o_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12682_ _12682_/A _24836_/B _12691_/B vssd1 vssd1 vccd1 vccd1 _12682_/X sky130_fd_sc_hd__and3_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24668_ hold2372/X _26285_/Q _24740_/S vssd1 vssd1 vccd1 vccd1 _24668_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _14419_/Y hold15/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__a21oi_1
X_23619_ hold2292/X hold1991/X _23677_/S vssd1 vssd1 vccd1 vccd1 _23620_/A sky130_fd_sc_hd__mux2_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24599_ _24599_/A vssd1 vssd1 vccd1 vccd1 _26262_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17140_ _25598_/Q vssd1 vssd1 vccd1 vccd1 _20625_/B sky130_fd_sc_hd__inv_2
XFILLER_0_107_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26338_ _26339_/CLK _26338_/D vssd1 vssd1 vccd1 vccd1 _26338_/Q sky130_fd_sc_hd__dfxtp_2
X_14352_ _14352_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14352_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_53_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13303_ _13303_/A vssd1 vssd1 vccd1 vccd1 _19560_/A sky130_fd_sc_hd__clkbuf_8
X_17071_ _25657_/Q _17071_/B vssd1 vssd1 vccd1 vccd1 _17441_/A sky130_fd_sc_hd__xor2_4
X_14283_ _25581_/Q _21228_/A vssd1 vssd1 vccd1 vccd1 _14590_/A sky130_fd_sc_hd__nand2_8
X_26269_ _26269_/CLK _26269_/D vssd1 vssd1 vccd1 vccd1 _26269_/Q sky130_fd_sc_hd__dfxtp_2
X_16022_ _16023_/B _16023_/A vssd1 vssd1 vccd1 vccd1 _16040_/B sky130_fd_sc_hd__or2_1
XFILLER_0_165_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13234_ _26303_/Q _19402_/A vssd1 vssd1 vccd1 vccd1 _14572_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_66_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13165_ _26292_/Q _19244_/A vssd1 vssd1 vccd1 vccd1 _14539_/A sky130_fd_sc_hd__xor2_1
X_13096_ _23377_/B vssd1 vssd1 vccd1 vccd1 _13096_/X sky130_fd_sc_hd__buf_6
X_17973_ _17973_/A _17973_/B vssd1 vssd1 vccd1 vccd1 _17974_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_137_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16924_ _16922_/X _16711_/X _16923_/Y _25893_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16925_/A sky130_fd_sc_hd__a32o_1
X_19712_ _26255_/Q hold380/X vssd1 vssd1 vccd1 vccd1 _19712_/Y sky130_fd_sc_hd__nand2_1
X_16855_ _16855_/A _16855_/B vssd1 vssd1 vccd1 vccd1 _16855_/Y sky130_fd_sc_hd__nand2_1
X_19643_ _19640_/Y _19643_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19643_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_189_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15806_ _15802_/Y _15803_/Y _15805_/X vssd1 vssd1 vccd1 vccd1 hold903/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19574_ _19574_/A _21291_/B vssd1 vssd1 vccd1 vccd1 _19574_/Y sky130_fd_sc_hd__nor2_1
X_16786_ _16787_/B _16787_/A vssd1 vssd1 vccd1 vccd1 _16786_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13998_ _14061_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13998_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_189_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18525_ _18528_/A _18529_/B vssd1 vssd1 vccd1 vccd1 _18527_/A sky130_fd_sc_hd__nand2_1
X_15737_ _26040_/Q _25976_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15738_/A sky130_fd_sc_hd__mux2_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12949_ _17471_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12949_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_72_clk _25759_/CLK vssd1 vssd1 vccd1 vccd1 _25901_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_157_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18456_ _18454_/X _18269_/X _18455_/X vssd1 vssd1 vccd1 vccd1 _18457_/A sky130_fd_sc_hd__a21o_1
X_15668_ _23063_/B _15668_/B vssd1 vssd1 vccd1 vccd1 _23060_/B sky130_fd_sc_hd__xor2_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_1_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_17407_ _17467_/A _17407_/B vssd1 vssd1 vccd1 vccd1 _17407_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_56_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14619_ _14617_/Y hold315/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold316/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18387_ _18952_/A _18387_/B _18952_/C vssd1 vssd1 vccd1 vccd1 _18388_/C sky130_fd_sc_hd__nand3_1
X_15599_ _22996_/B _16369_/B vssd1 vssd1 vccd1 vccd1 _16532_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_157_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17338_ _25613_/Q vssd1 vssd1 vccd1 vccd1 _21102_/B sky130_fd_sc_hd__inv_2
XFILLER_0_16_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17269_ _17393_/A _17269_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17269_/X sky130_fd_sc_hd__and3_1
XFILLER_0_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19008_ _19186_/A _19774_/A vssd1 vssd1 vccd1 vccd1 _19008_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20280_ _20280_/A _20280_/B vssd1 vssd1 vccd1 vccd1 _20282_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2603 _24701_/X vssd1 vssd1 vccd1 vccd1 _24702_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2614 _25437_/Q vssd1 vssd1 vccd1 vccd1 _15133_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2625 _26309_/Q vssd1 vssd1 vccd1 vccd1 hold2625/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2636 _26319_/Q vssd1 vssd1 vccd1 vccd1 hold2636/X sky130_fd_sc_hd__dlygate4sd3_1
X_23970_ _23970_/A vssd1 vssd1 vccd1 vccd1 _26058_/D sky130_fd_sc_hd__clkbuf_1
Xhold1902 _25707_/Q vssd1 vssd1 vccd1 vccd1 _19071_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2647 _26245_/Q vssd1 vssd1 vccd1 vccd1 hold2647/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1913 _23911_/X vssd1 vssd1 vccd1 vccd1 _23912_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2658 _24538_/X vssd1 vssd1 vccd1 vccd1 _24539_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1924 _26003_/Q vssd1 vssd1 vccd1 vccd1 _14893_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2669 _15324_/Y vssd1 vssd1 vccd1 vccd1 hold2669/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1935 _23914_/X vssd1 vssd1 vccd1 vccd1 _23915_/A sky130_fd_sc_hd__dlygate4sd3_1
X_22921_ _22919_/X _22920_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _22921_/Y sky130_fd_sc_hd__a21oi_1
Xhold1946 _24651_/X vssd1 vssd1 vccd1 vccd1 _24653_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1957 _25974_/Q vssd1 vssd1 vccd1 vccd1 hold1957/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1968 _23806_/X vssd1 vssd1 vccd1 vccd1 _23807_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1979 _23917_/X vssd1 vssd1 vccd1 vccd1 _23918_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25640_ _26146_/CLK _25640_/D vssd1 vssd1 vccd1 vccd1 _25640_/Q sky130_fd_sc_hd__dfxtp_2
X_22852_ _16837_/B _22421_/X _22845_/X _22846_/Y _22851_/X vssd1 vssd1 vccd1 vccd1
+ _22853_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_116_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21803_ _21803_/A _21803_/B vssd1 vssd1 vccd1 vccd1 _21803_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_149_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25571_ _26066_/CLK _25571_/D vssd1 vssd1 vccd1 vccd1 _25571_/Q sky130_fd_sc_hd__dfxtp_1
X_22783_ _22782_/A _22454_/X _22782_/B vssd1 vssd1 vccd1 vccd1 _22784_/C sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_63_clk clkbuf_leaf_95_clk/A vssd1 vssd1 vccd1 vccd1 _25511_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24522_ _24522_/A vssd1 vssd1 vccd1 vccd1 _26237_/D sky130_fd_sc_hd__clkbuf_1
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21734_ _21734_/A _21734_/B vssd1 vssd1 vccd1 vccd1 _21735_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24453_ _24453_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24454_/A sky130_fd_sc_hd__and2_1
X_21665_ _26337_/Q _19130_/X hold845/X vssd1 vssd1 vccd1 vccd1 _21668_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23404_ _24940_/S hold332/A _23403_/X vssd1 vssd1 vccd1 vccd1 _23404_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_164_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20616_ _26292_/Q _20078_/X hold853/X vssd1 vssd1 vccd1 vccd1 _20619_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21596_ _21596_/A _21645_/B vssd1 vssd1 vccd1 vccd1 _21597_/C sky130_fd_sc_hd__nand2_1
X_24384_ _24384_/A vssd1 vssd1 vccd1 vccd1 _26192_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26123_ _26216_/CLK _26123_/D vssd1 vssd1 vccd1 vccd1 _26123_/Q sky130_fd_sc_hd__dfxtp_1
X_23335_ _23333_/X hold953/X _12702_/A vssd1 vssd1 vccd1 vccd1 hold954/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_144_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20547_ _20547_/A _20547_/B vssd1 vssd1 vccd1 vccd1 _20551_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26054_ _26057_/CLK _26054_/D vssd1 vssd1 vccd1 vccd1 _26054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23266_ hold875/X _23581_/B vssd1 vssd1 vccd1 vccd1 _23275_/A sky130_fd_sc_hd__nand2_1
X_20478_ _20478_/A _22408_/B vssd1 vssd1 vccd1 vccd1 _20479_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_162_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25005_ _26121_/CLK hold989/X vssd1 vssd1 vccd1 vccd1 hold988/A sky130_fd_sc_hd__dfxtp_1
X_22217_ _22703_/A _22858_/B vssd1 vssd1 vccd1 vccd1 _22227_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_123_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23197_ _23197_/A _23197_/B vssd1 vssd1 vccd1 vccd1 _23197_/Y sky130_fd_sc_hd__nand2_1
X_22148_ _22148_/A _25879_/Q vssd1 vssd1 vccd1 vccd1 _22148_/Y sky130_fd_sc_hd__nand2_1
X_14970_ _14968_/X _14969_/Y _14928_/X vssd1 vssd1 vccd1 vccd1 _25420_/D sky130_fd_sc_hd__a21oi_1
X_22079_ _25656_/Q _22078_/A _22078_/Y vssd1 vssd1 vccd1 vccd1 _22081_/A sky130_fd_sc_hd__o21ai_1
X_25907_ _26004_/CLK _25907_/D vssd1 vssd1 vccd1 vccd1 _25907_/Q sky130_fd_sc_hd__dfxtp_1
X_13921_ _18158_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13921_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_92_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16640_ _16640_/A hold920/X vssd1 vssd1 vccd1 vccd1 _16641_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25838_ _25838_/CLK _25838_/D vssd1 vssd1 vccd1 vccd1 _25838_/Q sky130_fd_sc_hd__dfxtp_4
X_13852_ _18914_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13852_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12803_ _26224_/Q _25593_/Q vssd1 vssd1 vccd1 vccd1 _14322_/A sky130_fd_sc_hd__xor2_2
X_16571_ _16676_/A _16571_/B vssd1 vssd1 vccd1 vccd1 _16573_/A sky130_fd_sc_hd__or2_1
XFILLER_0_97_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13783_ _26263_/Q _13612_/X _13605_/X _13782_/Y vssd1 vssd1 vccd1 vccd1 _13784_/B
+ sky130_fd_sc_hd__a22o_1
X_25769_ _25770_/CLK _25769_/D vssd1 vssd1 vccd1 vccd1 _25769_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_54_clk _25472_/CLK vssd1 vssd1 vccd1 vccd1 _26069_/CLK sky130_fd_sc_hd__clkbuf_16
X_18310_ _18310_/A _21101_/A vssd1 vssd1 vccd1 vccd1 _18657_/A sky130_fd_sc_hd__xor2_4
X_15522_ _26028_/Q _25964_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15523_/A sky130_fd_sc_hd__mux2_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12734_ _14279_/B _14277_/B _25259_/Q _23199_/C vssd1 vssd1 vccd1 vccd1 _14266_/A
+ sky130_fd_sc_hd__a31o_1
X_19290_ _20701_/A _22308_/B _25600_/Q vssd1 vssd1 vccd1 vccd1 _20705_/C sky130_fd_sc_hd__nand3_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ _18241_/A _21045_/B _18241_/C vssd1 vssd1 vccd1 vccd1 _21027_/B sky130_fd_sc_hd__nand3_2
X_15453_ _15453_/A _15776_/B vssd1 vssd1 vccd1 vccd1 _15454_/B sky130_fd_sc_hd__nand2_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _12671_/C _12666_/A vssd1 vssd1 vccd1 vccd1 _12667_/A sky130_fd_sc_hd__or2_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14404_ _14404_/A hold329/X vssd1 vssd1 vccd1 vccd1 hold330/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18172_ _18955_/A _18172_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18173_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_65_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15384_ _22799_/B _15384_/B vssd1 vssd1 vccd1 vccd1 _22796_/B sky130_fd_sc_hd__xor2_1
X_12596_ _12646_/A _12644_/B vssd1 vssd1 vccd1 vccd1 _12596_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_26_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17123_ _17121_/X _23187_/B _17122_/X vssd1 vssd1 vccd1 vccd1 _17124_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14335_ _14344_/A hold245/X vssd1 vssd1 vccd1 vccd1 hold246/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold509 hold509/A vssd1 vssd1 vccd1 vccd1 hold509/X sky130_fd_sc_hd__dlygate4sd3_1
X_17054_ _20390_/B _25848_/Q _20426_/B vssd1 vssd1 vccd1 vccd1 _17055_/B sky130_fd_sc_hd__mux2_2
X_14266_ _14266_/A _15839_/B vssd1 vssd1 vccd1 vccd1 _14266_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_122_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16005_ _16006_/B _16006_/A vssd1 vssd1 vccd1 vccd1 _16007_/A sky130_fd_sc_hd__or2_1
X_13217_ _26172_/Q _13065_/X _13216_/X vssd1 vssd1 vccd1 vccd1 _13217_/X sky130_fd_sc_hd__a21o_1
X_14197_ _26329_/Q _13518_/B _14170_/X _14196_/Y vssd1 vssd1 vccd1 vccd1 _14198_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _13049_/X _14529_/A _13067_/X _19206_/A vssd1 vssd1 vccd1 vccd1 _13148_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17956_ _18528_/A _25730_/Q vssd1 vssd1 vccd1 vccd1 _17958_/A sky130_fd_sc_hd__nand2_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _26148_/Q _13065_/X _13078_/X vssd1 vssd1 vccd1 vccd1 _13079_/X sky130_fd_sc_hd__a21o_1
Xhold1209 _25081_/Q vssd1 vssd1 vccd1 vccd1 _18333_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16907_ _16977_/A _25569_/Q vssd1 vssd1 vccd1 vccd1 _16907_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_139_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17887_ _20468_/B _19206_/A vssd1 vssd1 vccd1 vccd1 _17888_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19626_ _26249_/Q _19483_/X hold665/X vssd1 vssd1 vccd1 vccd1 _19626_/Y sky130_fd_sc_hd__a21oi_1
X_16838_ _16411_/B _16837_/Y _15621_/A vssd1 vssd1 vccd1 vccd1 _16838_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_189_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16769_ _16767_/X _16711_/X _16768_/Y _25870_/Q _14170_/X vssd1 vssd1 vccd1 vccd1
+ _16770_/A sky130_fd_sc_hd__a32o_1
X_19557_ _26244_/Q hold674/X vssd1 vssd1 vccd1 vccd1 _19557_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_189_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_45_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _26073_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18508_ _18954_/A _25751_/Q vssd1 vssd1 vccd1 vccd1 _18510_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19488_ _19488_/A _21129_/B vssd1 vssd1 vccd1 vccd1 _19488_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18439_ _18437_/Y _18438_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25666_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21450_ _21450_/A _21499_/A vssd1 vssd1 vccd1 vccd1 _21451_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_185_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20401_ _20401_/A _20401_/B vssd1 vssd1 vccd1 vccd1 _20405_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21381_ _21379_/Y _21380_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21381_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_160_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23120_ _23120_/A _23120_/B vssd1 vssd1 vccd1 vccd1 _23121_/B sky130_fd_sc_hd__nand2_1
X_20332_ _21172_/B _21499_/A vssd1 vssd1 vccd1 vccd1 _20335_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_114_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23051_ _23051_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _23051_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20263_ _20263_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20268_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22002_ _22002_/A _22145_/B vssd1 vssd1 vccd1 vccd1 _22002_/Y sky130_fd_sc_hd__nand2_1
X_20194_ _21042_/A _20194_/B _20193_/X vssd1 vssd1 vccd1 vccd1 _20195_/B sky130_fd_sc_hd__or3b_1
Xhold2400 _26174_/Q vssd1 vssd1 vccd1 vccd1 hold2400/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2411 _25666_/Q vssd1 vssd1 vccd1 vccd1 _13195_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2422 _26061_/Q vssd1 vssd1 vccd1 vccd1 hold2422/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2433 _15678_/Y vssd1 vssd1 vccd1 vccd1 hold2433/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2444 _15701_/Y vssd1 vssd1 vccd1 vccd1 hold2444/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2455 _25674_/Q vssd1 vssd1 vccd1 vccd1 _13247_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1710 _25638_/Q vssd1 vssd1 vccd1 vccd1 _17605_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2466 _26063_/Q vssd1 vssd1 vccd1 vccd1 hold2466/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1721 _25611_/Q vssd1 vssd1 vccd1 vccd1 _17396_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23953_ hold2368/X hold1799/X _24001_/S vssd1 vssd1 vccd1 vccd1 _23954_/A sky130_fd_sc_hd__mux2_1
Xhold1732 _25587_/Q vssd1 vssd1 vccd1 vccd1 _17096_/B sky130_fd_sc_hd__clkbuf_2
Xhold2477 _24734_/X vssd1 vssd1 vccd1 vccd1 _24735_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1743 _21100_/Y vssd1 vssd1 vccd1 vccd1 _25804_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2488 _25465_/Q vssd1 vssd1 vccd1 vccd1 _15631_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2499 _24986_/Q vssd1 vssd1 vccd1 vccd1 _12671_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1754 _14978_/Y vssd1 vssd1 vccd1 vccd1 _25421_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22904_ _22902_/Y _22903_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _22904_/Y sky130_fd_sc_hd__a21oi_1
Xhold1765 _25637_/Q vssd1 vssd1 vccd1 vccd1 _17598_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1776 _25864_/Q vssd1 vssd1 vccd1 vccd1 _22510_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1787 _25870_/Q vssd1 vssd1 vccd1 vccd1 _22662_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_23884_ _23884_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23885_/A sky130_fd_sc_hd__and2_1
Xhold1798 _25657_/Q vssd1 vssd1 vccd1 vccd1 _18252_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25623_ _26216_/CLK _25623_/D vssd1 vssd1 vccd1 vccd1 _25623_/Q sky130_fd_sc_hd__dfxtp_4
X_22835_ _16834_/B _22421_/X _22828_/X _22830_/Y _22834_/X vssd1 vssd1 vccd1 vccd1
+ _22836_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_6_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_clk _25184_/CLK vssd1 vssd1 vccd1 vccd1 _25770_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25554_ _25877_/CLK _25554_/D vssd1 vssd1 vccd1 vccd1 _25554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22766_ _22766_/A _22766_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22768_/A sky130_fd_sc_hd__or3_1
XFILLER_0_94_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24505_ _24505_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24506_/A sky130_fd_sc_hd__and2_1
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21717_ _21717_/A _21717_/B vssd1 vssd1 vccd1 vccd1 _21718_/A sky130_fd_sc_hd__nand2_1
X_25485_ _25925_/CLK hold930/X vssd1 vssd1 vccd1 vccd1 hold929/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22697_ _22697_/A _22697_/B vssd1 vssd1 vccd1 vccd1 _22698_/B sky130_fd_sc_hd__nand2_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24436_ _24835_/S vssd1 vssd1 vccd1 vccd1 _24510_/S sky130_fd_sc_hd__buf_12
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21648_ _21648_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _21653_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24367_ _24367_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24368_/A sky130_fd_sc_hd__and2_1
XFILLER_0_117_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_80 _25837_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21579_ _21579_/A _21629_/B vssd1 vssd1 vccd1 vccd1 _21580_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_105_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14120_ _14120_/A vssd1 vssd1 vccd1 vccd1 _14232_/B sky130_fd_sc_hd__buf_4
X_26106_ _26231_/CLK _26106_/D vssd1 vssd1 vccd1 vccd1 _26106_/Q sky130_fd_sc_hd__dfxtp_1
X_23318_ _23320_/B _23320_/A vssd1 vssd1 vccd1 vccd1 _23324_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_22_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24298_ _24298_/A vssd1 vssd1 vccd1 vccd1 _26164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26037_ _26041_/CLK _26037_/D vssd1 vssd1 vccd1 vccd1 _26037_/Q sky130_fd_sc_hd__dfxtp_1
X_14051_ _14118_/A hold512/X vssd1 vssd1 vccd1 vccd1 hold513/A sky130_fd_sc_hd__nand2_1
X_23249_ _23249_/A _24870_/B vssd1 vssd1 vccd1 vccd1 _23249_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13002_ _26262_/Q _25631_/Q vssd1 vssd1 vccd1 vccd1 _14443_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_120_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17810_ _18612_/A _25727_/Q _18083_/C vssd1 vssd1 vccd1 vccd1 _17811_/C sky130_fd_sc_hd__nand3_1
X_18790_ _18952_/A _25765_/Q _18891_/C vssd1 vssd1 vccd1 vccd1 _18791_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17741_ _17771_/A _17745_/B vssd1 vssd1 vccd1 vccd1 _17743_/A sky130_fd_sc_hd__nand2_1
X_14953_ _14951_/X hold2338/X _14928_/X vssd1 vssd1 vccd1 vccd1 _14953_/Y sky130_fd_sc_hd__a21oi_1
X_13904_ _13941_/A _13904_/B vssd1 vssd1 vccd1 vccd1 _13904_/Y sky130_fd_sc_hd__nand2_1
X_17672_ _25848_/Q _22075_/A vssd1 vssd1 vccd1 vccd1 _17803_/A sky130_fd_sc_hd__or2_2
X_14884_ _15839_/A _14884_/B vssd1 vssd1 vccd1 vccd1 _22366_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_89_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16623_ _16621_/X _16622_/Y _16594_/X vssd1 vssd1 vccd1 vccd1 hold888/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19411_ _19409_/Y _19410_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19411_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_173_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13835_ _26271_/Q _13801_/X _13793_/X _13834_/Y vssd1 vssd1 vccd1 vccd1 _13836_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_187_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_27_clk _25759_/CLK vssd1 vssd1 vccd1 vccd1 _25756_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_187_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16554_ _16554_/A _16554_/B vssd1 vssd1 vccd1 vccd1 _16555_/A sky130_fd_sc_hd__nand2_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19342_ _26229_/Q hold849/X vssd1 vssd1 vccd1 vccd1 _19342_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13766_ hold672/X _13765_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold673/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15505_ _15551_/B _15503_/Y _15504_/Y vssd1 vssd1 vccd1 vccd1 _15505_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_57_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12717_ hold410/X _12718_/A vssd1 vssd1 vccd1 vccd1 _12717_/X sky130_fd_sc_hd__or2_1
X_19273_ _19271_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19274_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16485_ _16485_/A vssd1 vssd1 vccd1 vccd1 _16492_/B sky130_fd_sc_hd__inv_2
XFILLER_0_57_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13697_ _13703_/A _13697_/B vssd1 vssd1 vccd1 vccd1 _13697_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_85_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18224_ _18224_/A _18224_/B _18224_/C vssd1 vssd1 vccd1 vccd1 _22008_/A sky130_fd_sc_hd__nand3_2
X_15436_ _22845_/B _16369_/B vssd1 vssd1 vccd1 vccd1 _16411_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_66_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12648_ _12648_/A vssd1 vssd1 vccd1 vccd1 _12711_/D sky130_fd_sc_hd__inv_2
XFILLER_0_182_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18155_ _18155_/A _18155_/B vssd1 vssd1 vccd1 vccd1 _18159_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15367_ _22782_/B _15367_/B vssd1 vssd1 vccd1 vccd1 _22779_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12579_ _23924_/A _12582_/A vssd1 vssd1 vccd1 vccd1 _12587_/A sky130_fd_sc_hd__or2_1
XFILLER_0_0_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17106_ _19701_/A _17106_/B vssd1 vssd1 vccd1 vccd1 _17534_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14318_ _14316_/Y hold204/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold205/A sky130_fd_sc_hd__a21oi_1
X_18086_ _18529_/A _18086_/B _18529_/C vssd1 vssd1 vccd1 vccd1 _18087_/C sky130_fd_sc_hd__nand3_1
X_15298_ _26015_/Q _25951_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15299_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold306 hold306/A vssd1 vssd1 vccd1 vccd1 hold306/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 hold317/A vssd1 vssd1 vccd1 vccd1 hold317/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold328 hold328/A vssd1 vssd1 vccd1 vccd1 hold328/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold339 hold339/A vssd1 vssd1 vccd1 vccd1 hold339/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17037_ _25591_/Q vssd1 vssd1 vccd1 vccd1 _20350_/B sky130_fd_sc_hd__inv_2
XFILLER_0_123_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14249_ _25835_/Q vssd1 vssd1 vccd1 vccd1 _18915_/B sky130_fd_sc_hd__inv_2
XFILLER_0_159_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _18988_/A _19059_/B vssd1 vssd1 vccd1 vccd1 _18989_/B sky130_fd_sc_hd__xnor2_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1006 _16484_/Y vssd1 vssd1 vccd1 vccd1 _25523_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1017 _25038_/Q vssd1 vssd1 vccd1 vccd1 _17457_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ _25851_/Q _22159_/A vssd1 vssd1 vccd1 vccd1 _17947_/A sky130_fd_sc_hd__or2_2
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1028 _13023_/X vssd1 vssd1 vccd1 vccd1 _25054_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 _25003_/Q vssd1 vssd1 vccd1 vccd1 _17029_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20950_ _21448_/C _21500_/B vssd1 vssd1 vccd1 vccd1 _20952_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19609_ _19601_/X _19608_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19609_/Y sky130_fd_sc_hd__o21ai_1
X_20881_ _20879_/Y _20880_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _20881_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_18_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _26151_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22620_ _22620_/A _22620_/B vssd1 vssd1 vccd1 vccd1 _22621_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22551_ _22551_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _22551_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_118_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21502_ _21502_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21507_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_119_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25270_ _26103_/CLK hold205/X vssd1 vssd1 vccd1 vccd1 hold203/A sky130_fd_sc_hd__dfxtp_1
X_22482_ _16722_/B _22421_/X _22476_/X _22477_/Y _22481_/X vssd1 vssd1 vccd1 vccd1
+ _22483_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_17_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24221_ _24221_/A vssd1 vssd1 vccd1 vccd1 _26139_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21433_ _21433_/A _21481_/A vssd1 vssd1 vccd1 vccd1 _21435_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24152_ _24152_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24153_/A sky130_fd_sc_hd__and2_1
X_21364_ _21362_/Y _21363_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21364_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23103_ _23103_/A _23103_/B vssd1 vssd1 vccd1 vccd1 _23105_/A sky130_fd_sc_hd__nand2_1
X_20315_ _20318_/A _20318_/C vssd1 vssd1 vccd1 vccd1 _20316_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24083_ hold721/X hold2185/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24084_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21295_ _21297_/B _21297_/C vssd1 vssd1 vccd1 vccd1 _21296_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold840 hold840/A vssd1 vssd1 vccd1 vccd1 hold840/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 hold851/A vssd1 vssd1 vccd1 vccd1 hold851/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold862 hold862/A vssd1 vssd1 vccd1 vccd1 hold862/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 hold873/A vssd1 vssd1 vccd1 vccd1 hold873/X sky130_fd_sc_hd__dlygate4sd3_1
X_23034_ _16914_/B _22421_/A _23028_/X _23029_/Y _23033_/X vssd1 vssd1 vccd1 vccd1
+ _23035_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_130_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20246_ _21466_/A vssd1 vssd1 vccd1 vccd1 _21465_/A sky130_fd_sc_hd__inv_2
XFILLER_0_101_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold884 hold884/A vssd1 vssd1 vccd1 vccd1 hold884/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold895 hold895/A vssd1 vssd1 vccd1 vccd1 hold895/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20177_ _20177_/A _25842_/Q vssd1 vssd1 vccd1 vccd1 _20180_/C sky130_fd_sc_hd__nand2_1
Xhold2230 _25422_/Q vssd1 vssd1 vccd1 vccd1 _14980_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2241 _26186_/Q vssd1 vssd1 vccd1 vccd1 hold2241/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2252 _26110_/Q vssd1 vssd1 vccd1 vccd1 hold2252/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24985_ _24990_/CLK _24985_/D vssd1 vssd1 vccd1 vccd1 _24985_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2263 _26141_/Q vssd1 vssd1 vccd1 vccd1 hold2263/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2274 _26187_/Q vssd1 vssd1 vccd1 vccd1 hold2274/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2285 _25699_/Q vssd1 vssd1 vccd1 vccd1 _13401_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1540 _19340_/Y vssd1 vssd1 vccd1 vccd1 _25725_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2296 _25424_/Q vssd1 vssd1 vccd1 vccd1 _14996_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1551 _25569_/Q vssd1 vssd1 vccd1 vccd1 hold1551/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23936_ _23936_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23937_/A sky130_fd_sc_hd__and2_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1562 _25540_/Q vssd1 vssd1 vccd1 vccd1 _22423_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_157_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1573 _17017_/Y vssd1 vssd1 vccd1 vccd1 _25582_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1584 _25825_/Q vssd1 vssd1 vccd1 vccd1 _21525_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1595 _14276_/X vssd1 vssd1 vccd1 vccd1 _25259_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23867_ _23867_/A vssd1 vssd1 vccd1 vccd1 _26026_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25606_ _26240_/CLK _25606_/D vssd1 vssd1 vccd1 vccd1 _25606_/Q sky130_fd_sc_hd__dfxtp_4
X_13620_ _18138_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13620_/Y sky130_fd_sc_hd__nor2_1
X_22818_ _16827_/B _22421_/X _22812_/X _22813_/Y _22817_/X vssd1 vssd1 vccd1 vccd1
+ _22819_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23798_ _23798_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23799_/A sky130_fd_sc_hd__and2_1
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25537_ _25537_/CLK hold691/X vssd1 vssd1 vccd1 vccd1 hold689/A sky130_fd_sc_hd__dfxtp_1
X_13551_ _26226_/Q _13426_/X _13468_/X _13550_/Y vssd1 vssd1 vccd1 vccd1 _13552_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22749_ _26057_/Q vssd1 vssd1 vccd1 vccd1 _22750_/A sky130_fd_sc_hd__inv_2
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xascon_wrapper_20 vssd1 vssd1 vccd1 vccd1 io_oeb[6] ascon_wrapper_20/LO sky130_fd_sc_hd__conb_1
XFILLER_0_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ input7/X vssd1 vssd1 vccd1 vccd1 _23245_/A sky130_fd_sc_hd__buf_12
X_16270_ _16269_/X _16270_/B vssd1 vssd1 vccd1 vccd1 _16276_/B sky130_fd_sc_hd__and2b_1
X_25468_ _25533_/CLK _25468_/D vssd1 vssd1 vccd1 vccd1 _25468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13482_ _17877_/B _13518_/B vssd1 vssd1 vccd1 vccd1 _13482_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_180_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15221_ _15188_/X _15268_/B _15268_/C _15220_/X vssd1 vssd1 vccd1 vccd1 _15221_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_152_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24419_ _24419_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24420_/A sky130_fd_sc_hd__and2_1
XFILLER_0_63_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25399_ _25425_/CLK _25399_/D vssd1 vssd1 vccd1 vccd1 _25399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15152_ _26007_/Q _25943_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15153_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14103_ _26314_/Q _13988_/X _13981_/X _14102_/Y vssd1 vssd1 vccd1 vccd1 _14104_/B
+ sky130_fd_sc_hd__a22o_1
X_15083_ _15083_/A _15083_/B vssd1 vssd1 vccd1 vccd1 _15084_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19960_ _19961_/B _19961_/A vssd1 vssd1 vccd1 vccd1 _19960_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14034_ _18203_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14034_/Y sky130_fd_sc_hd__nor2_1
X_18911_ _18952_/A _25771_/Q _18952_/C vssd1 vssd1 vccd1 vccd1 _18912_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_129_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19891_ _19975_/A _19891_/B vssd1 vssd1 vccd1 vccd1 _19891_/Y sky130_fd_sc_hd__nand2_1
X_18842_ _18986_/A _19602_/A vssd1 vssd1 vccd1 vccd1 _18842_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_98_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15985_ _15985_/A _15985_/B vssd1 vssd1 vccd1 vccd1 _15986_/B sky130_fd_sc_hd__nand2_1
X_18773_ _18955_/A _18773_/B _18894_/C vssd1 vssd1 vccd1 vccd1 _18774_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_175_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14936_ _14934_/X hold2065/X _14928_/X vssd1 vssd1 vccd1 vccd1 _14936_/Y sky130_fd_sc_hd__a21oi_1
X_17724_ _17724_/A _17724_/B _17727_/A vssd1 vssd1 vccd1 vccd1 _17766_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_171_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14867_ _14873_/B _22323_/A vssd1 vssd1 vccd1 vccd1 _22322_/B sky130_fd_sc_hd__xnor2_2
X_17655_ _17655_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _17655_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_159_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16606_ _16608_/B _16608_/A vssd1 vssd1 vccd1 vccd1 _16607_/A sky130_fd_sc_hd__nor2_1
X_13818_ hold678/X _13817_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold679/A sky130_fd_sc_hd__a21oi_1
X_17586_ _17586_/A _17586_/B vssd1 vssd1 vccd1 vccd1 _17586_/X sky130_fd_sc_hd__xor2_2
X_14798_ _14804_/B _22091_/A vssd1 vssd1 vccd1 vccd1 _22090_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_187_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16537_ _16537_/A _16537_/B _16541_/B vssd1 vssd1 vccd1 vccd1 _16537_/Y sky130_fd_sc_hd__nand3_1
X_19325_ _19452_/A _19325_/B vssd1 vssd1 vccd1 vccd1 _19325_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_85_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13749_ _25755_/Q vssd1 vssd1 vccd1 vccd1 _18591_/B sky130_fd_sc_hd__inv_2
XFILLER_0_18_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16468_ _16468_/A _16468_/B vssd1 vssd1 vccd1 vccd1 _16470_/A sky130_fd_sc_hd__nand2_1
X_19256_ _19254_/Y hold892/X _19086_/X vssd1 vssd1 vccd1 vccd1 hold893/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_183_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15419_ _15419_/A _15774_/B vssd1 vssd1 vccd1 vccd1 _15420_/B sky130_fd_sc_hd__nand2_2
X_18207_ _19081_/A _18207_/B vssd1 vssd1 vccd1 vccd1 _18207_/X sky130_fd_sc_hd__xor2_1
X_19187_ _19185_/Y hold819/X _19086_/X vssd1 vssd1 vccd1 vccd1 hold820/A sky130_fd_sc_hd__a21oi_1
X_16399_ hold966/X vssd1 vssd1 vccd1 vccd1 _16399_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_182_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18138_ _18955_/A _18138_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18139_/C sky130_fd_sc_hd__nand3_1
Xhold103 hold103/A vssd1 vssd1 vccd1 vccd1 hold103/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 hold114/A vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 hold125/A vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__dlygate4sd3_1
X_18069_ _18071_/A _18118_/A vssd1 vssd1 vccd1 vccd1 _18070_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_7_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _26136_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold136 hold136/A vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 hold147/A vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold158 hold158/A vssd1 vssd1 vccd1 vccd1 hold158/X sky130_fd_sc_hd__dlygate4sd3_1
X_20100_ _20102_/B _20102_/C vssd1 vssd1 vccd1 vccd1 _20101_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_106_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold169 hold169/A vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
X_21080_ _21080_/A _21080_/B vssd1 vssd1 vccd1 vccd1 _21082_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_111_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20031_ _20031_/A _20949_/C _20031_/C vssd1 vssd1 vccd1 vccd1 _20032_/B sky130_fd_sc_hd__nand3_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24770_ _24770_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24771_/A sky130_fd_sc_hd__and2_1
X_21982_ _18390_/A _25809_/Q _21980_/Y _21981_/Y vssd1 vssd1 vccd1 vccd1 _21983_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_179_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23721_ _23721_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23722_/A sky130_fd_sc_hd__and2_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20933_ _21235_/A _20933_/B vssd1 vssd1 vccd1 vccd1 _20933_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_96_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23652_ _23652_/A vssd1 vssd1 vccd1 vccd1 _25956_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20864_ _20864_/A _20864_/B vssd1 vssd1 vccd1 vccd1 _21451_/B sky130_fd_sc_hd__nand2_4
X_22603_ _22653_/A _22603_/B vssd1 vssd1 vccd1 vccd1 _22603_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23583_ _25931_/Q _25930_/Q hold952/X _25928_/Q vssd1 vssd1 vccd1 vccd1 _23587_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_49_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20795_ _20795_/A _22620_/B _20795_/C vssd1 vssd1 vccd1 vccd1 _20798_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_119_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25322_ _26279_/CLK hold61/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22534_ _22586_/A vssd1 vssd1 vccd1 vccd1 _22534_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_107_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25253_ _25864_/CLK hold634/X vssd1 vssd1 vccd1 vccd1 hold632/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22465_ _22465_/A _22465_/B vssd1 vssd1 vccd1 vccd1 _22465_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24204_ _24204_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24205_/A sky130_fd_sc_hd__and2_1
XFILLER_0_134_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21416_ _21416_/A _21416_/B _21416_/C vssd1 vssd1 vccd1 vccd1 _21420_/A sky130_fd_sc_hd__nand3_1
X_25184_ _25184_/CLK hold945/X vssd1 vssd1 vccd1 vccd1 hold944/A sky130_fd_sc_hd__dfxtp_1
X_22396_ _22396_/A _22396_/B vssd1 vssd1 vccd1 vccd1 _22397_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_102_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24135_ _24135_/A vssd1 vssd1 vccd1 vccd1 _26111_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21347_ _21573_/A _21347_/B vssd1 vssd1 vccd1 vccd1 _21347_/Y sky130_fd_sc_hd__nand2_1
X_24066_ _24066_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24067_/A sky130_fd_sc_hd__and2_1
XFILLER_0_60_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21278_ _21643_/C _21691_/C vssd1 vssd1 vccd1 vccd1 _21279_/C sky130_fd_sc_hd__nand2_1
Xhold670 hold670/A vssd1 vssd1 vccd1 vccd1 hold670/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 hold681/A vssd1 vssd1 vccd1 vccd1 hold681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 hold692/A vssd1 vssd1 vccd1 vccd1 hold692/X sky130_fd_sc_hd__dlygate4sd3_1
X_23017_ _23017_/A _23193_/B _23017_/C vssd1 vssd1 vccd1 vccd1 _23017_/X sky130_fd_sc_hd__and3_1
XFILLER_0_120_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20229_ _20228_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20229_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2060 _23754_/X vssd1 vssd1 vccd1 vccd1 _23755_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2071 _25964_/Q vssd1 vssd1 vccd1 vccd1 hold2071/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2082 _25924_/Q vssd1 vssd1 vccd1 vccd1 _23305_/A sky130_fd_sc_hd__dlygate4sd3_1
X_15770_ _15768_/X _15769_/Y _15464_/X vssd1 vssd1 vccd1 vccd1 _25472_/D sky130_fd_sc_hd__a21oi_1
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2093 _23656_/X vssd1 vssd1 vccd1 vccd1 _23657_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24968_ _25378_/CLK _24968_/D vssd1 vssd1 vccd1 vccd1 _24968_/Q sky130_fd_sc_hd__dfxtp_1
X_12982_ _26258_/Q _25627_/Q vssd1 vssd1 vccd1 vccd1 _14431_/A sky130_fd_sc_hd__xor2_1
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1370 _14892_/Y vssd1 vssd1 vccd1 vccd1 _25410_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1381 _25472_/Q vssd1 vssd1 vccd1 vccd1 _15752_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _14900_/A _14721_/B vssd1 vssd1 vccd1 vccd1 _14721_/Y sky130_fd_sc_hd__nand2_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23919_ _23919_/A vssd1 vssd1 vccd1 vccd1 _26043_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1392 _13432_/X vssd1 vssd1 vccd1 vccd1 _25123_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24899_ _24895_/X _24898_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _24899_/X sky130_fd_sc_hd__mux2_2
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17440_ _17491_/A _17607_/B vssd1 vssd1 vccd1 vccd1 _17441_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _14688_/A hold173/X vssd1 vssd1 vccd1 vccd1 hold174/A sky130_fd_sc_hd__nand2_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13603_ hold564/X _13602_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold565/A sky130_fd_sc_hd__a21oi_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17371_ _17556_/A _17607_/B vssd1 vssd1 vccd1 vccd1 _17372_/B sky130_fd_sc_hd__xnor2_1
X_14583_ _14581_/Y hold93/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16322_ _16322_/A _16336_/A vssd1 vssd1 vccd1 vccd1 _16324_/A sky130_fd_sc_hd__nand2_1
X_19110_ _19101_/X _18879_/X _19109_/X vssd1 vssd1 vccd1 vccd1 _19111_/A sky130_fd_sc_hd__a21o_1
X_13534_ _13583_/A _13534_/B vssd1 vssd1 vccd1 vccd1 _13534_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_165_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19041_ _19039_/X _18879_/X _19040_/X vssd1 vssd1 vccd1 vccd1 _19042_/A sky130_fd_sc_hd__a21o_1
X_16253_ _16269_/B vssd1 vssd1 vccd1 vccd1 _16254_/B sky130_fd_sc_hd__inv_2
XFILLER_0_54_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13465_ _13465_/A _13465_/B vssd1 vssd1 vccd1 vccd1 _13466_/A sky130_fd_sc_hd__nand2_8
X_15204_ _15204_/A vssd1 vssd1 vccd1 vccd1 _15213_/B sky130_fd_sc_hd__inv_2
XFILLER_0_129_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16184_ _16184_/A _16189_/A vssd1 vssd1 vccd1 vccd1 _16184_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13396_ _26329_/Q _19774_/A vssd1 vssd1 vccd1 vccd1 _14654_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_51_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15135_ _26006_/Q _25942_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15137_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_51_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15066_ _15066_/A _15066_/B vssd1 vssd1 vccd1 vccd1 _15085_/A sky130_fd_sc_hd__nand2_1
X_19943_ _19941_/Y _19942_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _19943_/Y sky130_fd_sc_hd__a21oi_1
X_14017_ _26300_/Q _13988_/X _13981_/X _14016_/Y vssd1 vssd1 vccd1 vccd1 _14018_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19874_ _19875_/B _19875_/A vssd1 vssd1 vccd1 vccd1 _19874_/X sky130_fd_sc_hd__or2_1
X_18825_ _22564_/B _25639_/Q vssd1 vssd1 vccd1 vccd1 _18827_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_171_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18756_ _18756_/A _20557_/A vssd1 vssd1 vccd1 vccd1 _19010_/A sky130_fd_sc_hd__xor2_4
X_15968_ hold809/X vssd1 vssd1 vccd1 vccd1 _15971_/B sky130_fd_sc_hd__inv_2
XFILLER_0_78_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17707_ _23208_/B _17707_/B _17711_/A vssd1 vssd1 vccd1 vccd1 _17708_/A sky130_fd_sc_hd__or3_1
X_14919_ _14919_/A _14919_/B vssd1 vssd1 vccd1 vccd1 _14925_/A sky130_fd_sc_hd__nand2_1
X_15899_ _15900_/B _15900_/A vssd1 vssd1 vccd1 vccd1 _15901_/A sky130_fd_sc_hd__or2_1
X_18687_ _18687_/A _18687_/B vssd1 vssd1 vccd1 vccd1 _22390_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17638_ _17638_/A _17638_/B vssd1 vssd1 vccd1 vccd1 _17638_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17569_ _17566_/Y _17567_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _17569_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_175_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19308_ _19308_/A _19308_/B vssd1 vssd1 vccd1 vccd1 _19308_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20580_ _21042_/A _20580_/B _20579_/X vssd1 vssd1 vccd1 vccd1 _20581_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_74_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19239_ _19239_/A _19994_/B _19239_/C vssd1 vssd1 vccd1 vccd1 _19239_/X sky130_fd_sc_hd__and3_1
XFILLER_0_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22250_ _22250_/A _22250_/B vssd1 vssd1 vccd1 vccd1 _22250_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_108_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21201_ _26311_/Q _20731_/X hold789/X vssd1 vssd1 vccd1 vccd1 _21205_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22181_ _22181_/A _22181_/B vssd1 vssd1 vccd1 vccd1 _22181_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_83_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21132_ _25870_/Q _21132_/B _21132_/C vssd1 vssd1 vccd1 vccd1 _21136_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25940_ _26341_/CLK _25940_/D vssd1 vssd1 vccd1 vccd1 output9/A sky130_fd_sc_hd__dfxtp_2
X_21063_ _21063_/A _21063_/B vssd1 vssd1 vccd1 vccd1 _21064_/A sky130_fd_sc_hd__nand2_1
X_20014_ _25877_/Q _20014_/B _20014_/C vssd1 vssd1 vccd1 vccd1 _20018_/B sky130_fd_sc_hd__nand3b_1
X_25871_ _25876_/CLK _25871_/D vssd1 vssd1 vccd1 vccd1 _25871_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_119_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24822_ _24822_/A vssd1 vssd1 vccd1 vccd1 _26335_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24753_ _24753_/A vssd1 vssd1 vccd1 vccd1 _26312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21965_ _22058_/A _21965_/B vssd1 vssd1 vccd1 vccd1 _21965_/Y sky130_fd_sc_hd__nand2_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23704_ _23704_/A vssd1 vssd1 vccd1 vccd1 _25973_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ _20915_/B _20916_/B _20916_/C vssd1 vssd1 vccd1 vccd1 _20917_/B sky130_fd_sc_hd__nand3b_1
X_24684_ _24684_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24685_/A sky130_fd_sc_hd__and2_1
XFILLER_0_139_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21896_ _22058_/A _21896_/B vssd1 vssd1 vccd1 vccd1 _21896_/Y sky130_fd_sc_hd__nand2_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23635_ hold1926/X _25951_/Q _23677_/S vssd1 vssd1 vccd1 vccd1 _23635_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_138_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20847_ _26298_/Q _20731_/X hold554/X vssd1 vssd1 vccd1 vccd1 _20850_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23566_ _23560_/X _23565_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _23566_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20778_ _20776_/Y _20777_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _20778_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25305_ _25636_/CLK hold241/X vssd1 vssd1 vccd1 vccd1 hold239/A sky130_fd_sc_hd__dfxtp_1
X_22517_ _22518_/B _22518_/A vssd1 vssd1 vccd1 vccd1 _22519_/A sky130_fd_sc_hd__or2_1
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26285_ _26286_/CLK _26285_/D vssd1 vssd1 vccd1 vccd1 _26285_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_80_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23497_ hold8/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23497_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13250_ _26177_/Q _13239_/X _13249_/X vssd1 vssd1 vccd1 vccd1 _13250_/X sky130_fd_sc_hd__a21o_1
X_25236_ _25689_/CLK hold732/X vssd1 vssd1 vccd1 vccd1 hold731/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22448_ _22448_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _22448_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ _13109_/X _13179_/X _13096_/X _13180_/X vssd1 vssd1 vccd1 vccd1 _13181_/X
+ sky130_fd_sc_hd__o211a_1
X_25167_ _25779_/CLK hold574/X vssd1 vssd1 vccd1 vccd1 hold572/A sky130_fd_sc_hd__dfxtp_1
X_22379_ _22807_/B _22958_/B vssd1 vssd1 vccd1 vccd1 _22381_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_0_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24118_ _24118_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24119_/A sky130_fd_sc_hd__and2_1
XFILLER_0_32_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25098_ _26184_/CLK _25098_/D vssd1 vssd1 vccd1 vccd1 _25098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24049_ _24049_/A vssd1 vssd1 vccd1 vccd1 _26084_/D sky130_fd_sc_hd__clkbuf_1
X_16940_ _16977_/A _16940_/B vssd1 vssd1 vccd1 vccd1 _16940_/Y sky130_fd_sc_hd__nand2_1
X_16871_ _16871_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16871_/Y sky130_fd_sc_hd__nand2_1
X_18610_ _18610_/A _25820_/Q _18610_/C vssd1 vssd1 vccd1 vccd1 _20281_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_189_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15822_ _15822_/A _15822_/B vssd1 vssd1 vccd1 vccd1 _15826_/A sky130_fd_sc_hd__nand2_1
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19590_ _20010_/A _19588_/Y _20014_/C vssd1 vssd1 vccd1 vccd1 _19678_/B sky130_fd_sc_hd__o21a_2
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15753_ _16963_/B vssd1 vssd1 vccd1 vccd1 _23143_/B sky130_fd_sc_hd__inv_2
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18541_ _19644_/A vssd1 vssd1 vccd1 vccd1 _22208_/B sky130_fd_sc_hd__inv_2
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ _12930_/X _12963_/X _12917_/X _12964_/X vssd1 vssd1 vccd1 vccd1 _12965_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14704_ _14701_/Y _14703_/Y _14646_/X vssd1 vssd1 vccd1 vccd1 _14704_/Y sky130_fd_sc_hd__a21oi_1
X_15684_ _23079_/B _15684_/B vssd1 vssd1 vccd1 vccd1 _23076_/B sky130_fd_sc_hd__xor2_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18472_ _18472_/A _20010_/A vssd1 vssd1 vccd1 vccd1 _18818_/A sky130_fd_sc_hd__xor2_4
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _12840_/X _12894_/X _12827_/X _12895_/X vssd1 vssd1 vccd1 vccd1 _12896_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17423_ _17423_/A _17423_/B vssd1 vssd1 vccd1 vccd1 _17423_/X sky130_fd_sc_hd__xor2_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _14635_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14635_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_158_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17354_ _17352_/X _17241_/X _17353_/X vssd1 vssd1 vccd1 vccd1 _17355_/A sky130_fd_sc_hd__a21o_1
X_14566_ _14566_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14566_/Y sky130_fd_sc_hd__nand2_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16305_ _16306_/B _16306_/A vssd1 vssd1 vccd1 vccd1 _16336_/A sky130_fd_sc_hd__or2_1
X_13517_ hold922/A vssd1 vssd1 vccd1 vccd1 _18155_/B sky130_fd_sc_hd__inv_2
X_17285_ _19199_/A vssd1 vssd1 vccd1 vccd1 _17467_/A sky130_fd_sc_hd__clkbuf_8
X_14497_ _14497_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14497_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_153_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16236_ _16236_/A _16236_/B vssd1 vssd1 vccd1 vccd1 _16237_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19024_ _19024_/A _19074_/A vssd1 vssd1 vccd1 vccd1 _19025_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13448_ _26338_/Q _25707_/Q vssd1 vssd1 vccd1 vccd1 _14681_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_181_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16167_ _16167_/A vssd1 vssd1 vccd1 vccd1 _16182_/B sky130_fd_sc_hd__inv_2
XFILLER_0_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13379_ _13220_/X _14644_/A _13242_/X _19729_/A vssd1 vssd1 vccd1 vccd1 _13379_/X
+ sky130_fd_sc_hd__a22o_1
X_15118_ _22449_/B _15812_/B vssd1 vssd1 vccd1 vccd1 _16165_/B sky130_fd_sc_hd__nand2_1
X_16098_ _16103_/B _16099_/A vssd1 vssd1 vccd1 vccd1 _16098_/X sky130_fd_sc_hd__or2_1
X_15049_ _15049_/A _15049_/B vssd1 vssd1 vccd1 vccd1 _15050_/B sky130_fd_sc_hd__nand2_2
X_19926_ _19937_/A _19989_/B vssd1 vssd1 vccd1 vccd1 _19928_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_167_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19857_ _19857_/A _19980_/B _19857_/C vssd1 vssd1 vccd1 vccd1 _19857_/X sky130_fd_sc_hd__and3_1
XFILLER_0_76_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18808_ _25894_/Q _22538_/A vssd1 vssd1 vccd1 vccd1 _18816_/A sky130_fd_sc_hd__or2_2
X_19788_ _19788_/A _20558_/B vssd1 vssd1 vccd1 vccd1 _19788_/Y sky130_fd_sc_hd__nor2_1
X_18739_ _19026_/A _18739_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18739_/X sky130_fd_sc_hd__and3_1
XFILLER_0_92_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21750_ _17665_/B _17016_/B _17666_/B vssd1 vssd1 vccd1 vccd1 _21751_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_188_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20701_ _20701_/A _22308_/B vssd1 vssd1 vccd1 vccd1 _20702_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21681_ _26338_/Q _19130_/X hold650/X vssd1 vssd1 vccd1 vccd1 _21684_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_188_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23420_ hold326/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23420_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_114_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20632_ _20632_/A _20632_/B vssd1 vssd1 vccd1 vccd1 _21351_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23351_ _23351_/A _23351_/B vssd1 vssd1 vccd1 vccd1 _23356_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_149_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20563_ _20566_/A _20566_/C vssd1 vssd1 vccd1 vccd1 _20565_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_144_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22302_ _22302_/A _22302_/B vssd1 vssd1 vccd1 vccd1 _22303_/B sky130_fd_sc_hd__nand2_1
X_26070_ _26073_/CLK _26070_/D vssd1 vssd1 vccd1 vccd1 _26070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23282_ _23284_/A hold832/X vssd1 vssd1 vccd1 vccd1 hold833/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20494_ _21279_/B _21563_/A vssd1 vssd1 vccd1 vccd1 _20495_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_143_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25021_ _26231_/CLK _25021_/D vssd1 vssd1 vccd1 vccd1 _25021_/Q sky130_fd_sc_hd__dfxtp_1
X_22233_ _22233_/A _22387_/B vssd1 vssd1 vccd1 vccd1 _22233_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22164_ _22165_/B _22165_/A vssd1 vssd1 vccd1 vccd1 _22166_/A sky130_fd_sc_hd__or2_1
XFILLER_0_100_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21115_ _21545_/C _21597_/B vssd1 vssd1 vccd1 vccd1 _21117_/A sky130_fd_sc_hd__nand2_1
X_22095_ _25813_/Q _22095_/B vssd1 vssd1 vccd1 vccd1 _22095_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_10_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25923_ _25925_/CLK hold987/X vssd1 vssd1 vccd1 vccd1 hold985/A sky130_fd_sc_hd__dfxtp_1
X_21046_ _21044_/Y _21045_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _21046_/Y sky130_fd_sc_hd__a21oi_1
X_25854_ _26336_/CLK _25854_/D vssd1 vssd1 vccd1 vccd1 _25854_/Q sky130_fd_sc_hd__dfxtp_4
X_24805_ hold2712/X _26330_/Q _24817_/S vssd1 vssd1 vccd1 vccd1 _24805_/X sky130_fd_sc_hd__mux2_1
X_25785_ _25785_/CLK _25785_/D vssd1 vssd1 vccd1 vccd1 _25785_/Q sky130_fd_sc_hd__dfxtp_2
X_22997_ _15598_/B _22893_/A _22829_/X vssd1 vssd1 vccd1 vccd1 _22997_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12750_ _23193_/B _21203_/A _17008_/B vssd1 vssd1 vccd1 vccd1 _12751_/A sky130_fd_sc_hd__or3_1
X_24736_ _24736_/A vssd1 vssd1 vccd1 vccd1 _26307_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21948_ _18370_/A _25808_/Q _21946_/Y _21947_/Y vssd1 vssd1 vccd1 vccd1 _21949_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12681_ _12684_/A _12681_/B _12676_/B vssd1 vssd1 vccd1 vccd1 _12691_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_139_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24667_ _24743_/A vssd1 vssd1 vccd1 vccd1 _24740_/S sky130_fd_sc_hd__buf_12
XFILLER_0_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21879_ _18330_/A _25806_/Q _21877_/Y _21878_/Y vssd1 vssd1 vccd1 vccd1 _21880_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14465_/A hold14/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__nand2_1
X_23618_ _23618_/A vssd1 vssd1 vccd1 vccd1 _25945_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24598_ _24598_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24599_/A sky130_fd_sc_hd__and2_1
XFILLER_0_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26337_ _26339_/CLK _26337_/D vssd1 vssd1 vccd1 vccd1 _26337_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14351_ _14348_/Y hold27/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23549_ hold32/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23549_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_163_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13302_ _13207_/X _13298_/X _13300_/X _13301_/X vssd1 vssd1 vccd1 vccd1 _13302_/X
+ sky130_fd_sc_hd__o211a_1
X_17070_ _20429_/B _25849_/Q _25785_/Q vssd1 vssd1 vccd1 vccd1 _17071_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_165_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14282_ _21203_/A vssd1 vssd1 vccd1 vccd1 _21228_/A sky130_fd_sc_hd__buf_12
X_26268_ _26273_/CLK _26268_/D vssd1 vssd1 vccd1 vccd1 _26268_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_162_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16021_ _22173_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _16023_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_150_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13233_ _13233_/A vssd1 vssd1 vccd1 vccd1 _19402_/A sky130_fd_sc_hd__buf_4
X_25219_ _26303_/CLK hold439/X vssd1 vssd1 vccd1 vccd1 hold437/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26199_ _26200_/CLK _26199_/D vssd1 vssd1 vccd1 vccd1 _26199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13164_ _13164_/A vssd1 vssd1 vccd1 vccd1 _19244_/A sky130_fd_sc_hd__buf_4
XFILLER_0_21_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13095_ _26151_/Q _13065_/X _13094_/X vssd1 vssd1 vccd1 vccd1 _13095_/X sky130_fd_sc_hd__a21o_1
X_17972_ _17759_/A _17759_/C _17925_/B vssd1 vssd1 vccd1 vccd1 _17973_/A sky130_fd_sc_hd__a21o_1
X_19711_ _26255_/Q _19483_/X hold380/X vssd1 vssd1 vccd1 vccd1 _19711_/Y sky130_fd_sc_hd__a21oi_1
X_16923_ _16923_/A _16923_/B vssd1 vssd1 vccd1 vccd1 _16923_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_137_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_213_clk _26093_/CLK vssd1 vssd1 vccd1 vccd1 _26221_/CLK sky130_fd_sc_hd__clkbuf_16
X_19642_ _19641_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19643_/B
+ sky130_fd_sc_hd__a211o_1
X_16854_ _16855_/B _16855_/A vssd1 vssd1 vccd1 vccd1 _16854_/X sky130_fd_sc_hd__or2_1
X_15805_ _17568_/A vssd1 vssd1 vccd1 vccd1 _15805_/X sky130_fd_sc_hd__buf_8
X_19573_ _19570_/Y _19573_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19573_/X sky130_fd_sc_hd__and3b_1
X_16785_ _16980_/A _16790_/B vssd1 vssd1 vccd1 vccd1 _16787_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_137_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13997_ _26297_/Q _13988_/X _13981_/X _13996_/Y vssd1 vssd1 vccd1 vccd1 _13998_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18524_ _25880_/Q _22178_/A vssd1 vssd1 vccd1 vccd1 _18532_/A sky130_fd_sc_hd__or2_2
X_15736_ _16956_/B vssd1 vssd1 vccd1 vccd1 _23127_/B sky130_fd_sc_hd__inv_2
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12948_ _26123_/Q _12907_/X _12947_/X vssd1 vssd1 vccd1 vccd1 _12948_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18455_ _18535_/A _18455_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18455_/X sky130_fd_sc_hd__and3_1
X_15667_ _15667_/A _15774_/B vssd1 vssd1 vccd1 vccd1 _15668_/B sky130_fd_sc_hd__nand2_1
X_12879_ _17353_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12879_/X sky130_fd_sc_hd__or2_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17406_ _17406_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17406_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14618_ _14645_/A hold314/X vssd1 vssd1 vccd1 vccd1 hold315/A sky130_fd_sc_hd__nand2_1
X_15598_ _22999_/B _15598_/B vssd1 vssd1 vccd1 vccd1 _22996_/B sky130_fd_sc_hd__xor2_1
X_18386_ _18951_/A _19624_/B vssd1 vssd1 vccd1 vccd1 _18388_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_157_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14549_ _14585_/A hold344/X vssd1 vssd1 vccd1 vccd1 hold345/A sky130_fd_sc_hd__nand2_1
X_17337_ _17335_/Y _17336_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _17337_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17268_ _17492_/A _17268_/B vssd1 vssd1 vccd1 vccd1 _17268_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19007_ _19007_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _19007_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_24_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16219_ _16276_/A vssd1 vssd1 vccd1 vccd1 _16227_/B sky130_fd_sc_hd__inv_2
XFILLER_0_144_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17199_ _17456_/A _17199_/B vssd1 vssd1 vccd1 vccd1 _17199_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_144_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2604 _26310_/Q vssd1 vssd1 vccd1 vccd1 hold2604/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2615 _26264_/Q vssd1 vssd1 vccd1 vccd1 hold2615/X sky130_fd_sc_hd__dlygate4sd3_1
X_19909_ _19909_/A _19980_/B _19909_/C vssd1 vssd1 vccd1 vccd1 _19909_/X sky130_fd_sc_hd__and3_1
Xhold2626 _26241_/Q vssd1 vssd1 vccd1 vccd1 hold2626/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2637 _24775_/X vssd1 vssd1 vccd1 vccd1 _24776_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1903 _25965_/Q vssd1 vssd1 vccd1 vccd1 hold1903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2648 _26308_/Q vssd1 vssd1 vccd1 vccd1 hold2648/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2659 _26335_/Q vssd1 vssd1 vccd1 vccd1 hold2659/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_204_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _26103_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1914 _25692_/Q vssd1 vssd1 vccd1 vccd1 _13359_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1925 _23797_/X vssd1 vssd1 vccd1 vccd1 _23798_/A sky130_fd_sc_hd__dlygate4sd3_1
X_22920_ _22937_/A _22920_/B vssd1 vssd1 vccd1 vccd1 _22920_/Y sky130_fd_sc_hd__nand2_1
Xhold1936 _25959_/Q vssd1 vssd1 vccd1 vccd1 hold1936/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1947 _25949_/Q vssd1 vssd1 vccd1 vccd1 hold1947/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1958 _23708_/X vssd1 vssd1 vccd1 vccd1 _23709_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1969 _24969_/Q vssd1 vssd1 vccd1 vccd1 _12578_/A sky130_fd_sc_hd__dlygate4sd3_1
X_22851_ _22851_/A _23001_/B _22851_/C vssd1 vssd1 vccd1 vccd1 _22851_/X sky130_fd_sc_hd__and3_1
XFILLER_0_79_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21802_ _18005_/A _25795_/Q _21800_/Y _21801_/Y vssd1 vssd1 vccd1 vccd1 _21803_/B
+ sky130_fd_sc_hd__a31o_1
X_25570_ _25573_/CLK _25570_/D vssd1 vssd1 vccd1 vccd1 _25570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22782_ _22782_/A _22782_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22784_/A sky130_fd_sc_hd__or3_1
XFILLER_0_52_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24521_ _24521_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24522_/A sky130_fd_sc_hd__and2_1
XFILLER_0_176_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21733_ _21734_/B _21734_/A vssd1 vssd1 vccd1 vccd1 _21735_/A sky130_fd_sc_hd__or2_1
XFILLER_0_94_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24452_ hold2726/X hold2654/X _24510_/S vssd1 vssd1 vccd1 vccd1 _24453_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_148_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21664_ _21664_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _21669_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23403_ hold206/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23403_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20615_ _20615_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20620_/A sky130_fd_sc_hd__nand2_1
X_24383_ _24383_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24384_/A sky130_fd_sc_hd__and2_1
X_21595_ _21595_/A _21644_/B vssd1 vssd1 vccd1 vccd1 _21597_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_151_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26122_ _26122_/CLK _26122_/D vssd1 vssd1 vccd1 vccd1 _26122_/Q sky130_fd_sc_hd__dfxtp_1
X_23334_ _23334_/A hold952/X vssd1 vssd1 vccd1 vccd1 hold953/A sky130_fd_sc_hd__nand2_1
X_20546_ _20546_/A _22190_/B vssd1 vssd1 vccd1 vccd1 _20547_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26053_ _26053_/CLK _26053_/D vssd1 vssd1 vccd1 vccd1 _26053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23265_ _23263_/X hold876/X _12702_/A vssd1 vssd1 vccd1 vccd1 hold877/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_160_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20477_ _21279_/B vssd1 vssd1 vccd1 vccd1 _21276_/C sky130_fd_sc_hd__inv_2
XFILLER_0_162_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25004_ _26121_/CLK _25004_/D vssd1 vssd1 vccd1 vccd1 _25004_/Q sky130_fd_sc_hd__dfxtp_1
X_22216_ _22216_/A _22859_/A vssd1 vssd1 vccd1 vccd1 _22227_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_104_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23196_ _23187_/Y _23195_/Y _19199_/A vssd1 vssd1 vccd1 vccd1 _23196_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_113_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22147_ _22147_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _22147_/X sky130_fd_sc_hd__and2_1
XFILLER_0_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22078_ _22078_/A _22078_/B vssd1 vssd1 vccd1 vccd1 _22078_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_100_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25906_ _26269_/CLK _25906_/D vssd1 vssd1 vccd1 vccd1 _25906_/Q sky130_fd_sc_hd__dfxtp_1
X_13920_ _25782_/Q vssd1 vssd1 vccd1 vccd1 _18158_/B sky130_fd_sc_hd__inv_2
X_21029_ _21029_/A _21029_/B vssd1 vssd1 vccd1 vccd1 _21548_/B sky130_fd_sc_hd__nand2_2
X_13851_ _25771_/Q vssd1 vssd1 vccd1 vccd1 _18914_/B sky130_fd_sc_hd__inv_2
X_25837_ _25838_/CLK _25837_/D vssd1 vssd1 vccd1 vccd1 _25837_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_69_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12802_ _12746_/X _12800_/X _14910_/B _12801_/X vssd1 vssd1 vccd1 vccd1 _12802_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16570_ hold918/X vssd1 vssd1 vccd1 vccd1 _16573_/B sky130_fd_sc_hd__inv_2
X_13782_ _18693_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13782_/Y sky130_fd_sc_hd__nor2_1
X_25768_ _26275_/CLK _25768_/D vssd1 vssd1 vccd1 vccd1 _25768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15521_ _16872_/B vssd1 vssd1 vccd1 vccd1 _22931_/B sky130_fd_sc_hd__inv_2
X_12733_ _12733_/A vssd1 vssd1 vccd1 vccd1 _14279_/B sky130_fd_sc_hd__inv_2
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24719_ hold2594/X _26302_/Q _24740_/S vssd1 vssd1 vccd1 vccd1 _24719_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25699_ _25708_/CLK _25699_/D vssd1 vssd1 vccd1 vccd1 _25699_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15452_ _26024_/Q _25960_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15453_/A sky130_fd_sc_hd__mux2_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18240_ _18446_/A _25738_/Q _21716_/A vssd1 vssd1 vccd1 vccd1 _18241_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_84_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12664_ _12664_/A _12664_/B vssd1 vssd1 vccd1 vccd1 _12666_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_155_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14403_ _14403_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14403_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_167_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15383_ _15383_/A _15776_/B vssd1 vssd1 vccd1 vccd1 _15384_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18171_ _18954_/A _25735_/Q vssd1 vssd1 vccd1 vccd1 _18173_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_170_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12595_ _12644_/B _12646_/A vssd1 vssd1 vccd1 vccd1 _12601_/A sky130_fd_sc_hd__or2_1
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17122_ _17393_/A _17122_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17122_/X sky130_fd_sc_hd__and3_1
X_14334_ _14334_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14334_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_107_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17053_ _25592_/Q vssd1 vssd1 vccd1 vccd1 _20390_/B sky130_fd_sc_hd__inv_2
X_14265_ hold426/X _14264_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold427/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16004_ _16001_/Y _15953_/B _16056_/B vssd1 vssd1 vccd1 vccd1 _16006_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_123_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13216_ _13049_/X _14563_/A _13067_/X _19359_/A vssd1 vssd1 vccd1 vccd1 _13216_/X
+ sky130_fd_sc_hd__a22o_1
X_14196_ _18734_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14196_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _26289_/Q _19206_/A vssd1 vssd1 vccd1 vccd1 _14529_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17955_ _17955_/A _20815_/B _17955_/C vssd1 vssd1 vccd1 vccd1 _20786_/B sky130_fd_sc_hd__nand3_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _13049_/X _14488_/A _13067_/X _25645_/Q vssd1 vssd1 vccd1 vccd1 _13078_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16906_ _16906_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16906_/Y sky130_fd_sc_hd__nand2_1
X_17886_ _22131_/B _25594_/Q vssd1 vssd1 vccd1 vccd1 _17888_/A sky130_fd_sc_hd__nand2_1
X_19625_ _19623_/Y _19624_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19625_/Y sky130_fd_sc_hd__a21oi_1
X_16837_ _16980_/A _16837_/B vssd1 vssd1 vccd1 vccd1 _16837_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_178_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19556_ _26244_/Q _19483_/X hold674/X vssd1 vssd1 vccd1 vccd1 _19556_/Y sky130_fd_sc_hd__a21oi_1
X_16768_ _16768_/A _16768_/B vssd1 vssd1 vccd1 vccd1 _16768_/Y sky130_fd_sc_hd__nand2_1
X_18507_ _18507_/A _25815_/Q _18507_/C vssd1 vssd1 vccd1 vccd1 _20106_/C sky130_fd_sc_hd__nand3_2
X_15719_ _15691_/A _15718_/B _15713_/A vssd1 vssd1 vccd1 vccd1 _15719_/X sky130_fd_sc_hd__o21a_1
X_19487_ _19484_/Y _19487_/B _19980_/B vssd1 vssd1 vccd1 vccd1 _19487_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_88_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16699_ _16697_/Y hold576/X _16594_/X vssd1 vssd1 vccd1 vccd1 hold577/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18438_ _18641_/A _19317_/A vssd1 vssd1 vccd1 vccd1 _18438_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_91_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18369_ _21189_/B _21949_/A vssd1 vssd1 vccd1 vccd1 _21183_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_145_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20400_ _20400_/A _22370_/B vssd1 vssd1 vccd1 vccd1 _20401_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_114_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21380_ _21573_/A _21380_/B vssd1 vssd1 vccd1 vccd1 _21380_/Y sky130_fd_sc_hd__nand2_1
X_20331_ _20331_/A _20331_/B vssd1 vssd1 vccd1 vccd1 _21499_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_109_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23050_ _15647_/A _22421_/A _23044_/X _23045_/Y _23049_/X vssd1 vssd1 vccd1 vccd1
+ _23050_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_4_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20262_ _20262_/A _20262_/B vssd1 vssd1 vccd1 vccd1 _20263_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_113_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22001_ _22653_/A _22001_/B vssd1 vssd1 vccd1 vccd1 _22001_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20193_ _20191_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20193_/X
+ sky130_fd_sc_hd__a211o_1
Xhold2401 _26050_/Q vssd1 vssd1 vccd1 vccd1 hold2401/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2412 _26176_/Q vssd1 vssd1 vccd1 vccd1 hold2412/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2423 _23977_/X vssd1 vssd1 vccd1 vccd1 _23978_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2434 _15679_/Y vssd1 vssd1 vccd1 vccd1 _25467_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2445 _15702_/Y vssd1 vssd1 vccd1 vccd1 _25468_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1700 _25612_/Q vssd1 vssd1 vccd1 vccd1 _17407_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1711 _25828_/Q vssd1 vssd1 vccd1 vccd1 _21573_/B sky130_fd_sc_hd__dlygate4sd3_1
X_23952_ _23952_/A vssd1 vssd1 vccd1 vccd1 _26052_/D sky130_fd_sc_hd__clkbuf_1
Xhold2456 _26045_/Q vssd1 vssd1 vccd1 vccd1 hold2456/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1722 _17397_/Y vssd1 vssd1 vccd1 vccd1 _25611_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2467 _25679_/Q vssd1 vssd1 vccd1 vccd1 _13277_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2478 _26067_/Q vssd1 vssd1 vccd1 vccd1 hold2478/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1733 _17097_/Y vssd1 vssd1 vccd1 vccd1 _25587_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2489 _15644_/X vssd1 vssd1 vccd1 vccd1 hold2489/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1744 _25872_/Q vssd1 vssd1 vccd1 vccd1 _22715_/B sky130_fd_sc_hd__buf_1
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22903_ _22937_/A _22903_/B vssd1 vssd1 vccd1 vccd1 _22903_/Y sky130_fd_sc_hd__nand2_1
Xhold1755 _25624_/Q vssd1 vssd1 vccd1 vccd1 _17503_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1766 _25866_/Q vssd1 vssd1 vccd1 vccd1 _22561_/B sky130_fd_sc_hd__buf_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23883_ hold2177/X hold1932/X _23907_/S vssd1 vssd1 vccd1 vccd1 _23884_/A sky130_fd_sc_hd__mux2_1
Xhold1777 _22511_/Y vssd1 vssd1 vccd1 vccd1 _25864_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1788 _22663_/Y vssd1 vssd1 vccd1 vccd1 _25870_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1799 _26053_/Q vssd1 vssd1 vccd1 vccd1 hold1799/X sky130_fd_sc_hd__dlygate4sd3_1
X_22834_ _22834_/A _23001_/B _22834_/C vssd1 vssd1 vccd1 vccd1 _22834_/X sky130_fd_sc_hd__and3_1
X_25622_ _25716_/CLK _25622_/D vssd1 vssd1 vccd1 vccd1 _25622_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25553_ _25877_/CLK _25553_/D vssd1 vssd1 vccd1 vccd1 _25553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22765_ _26058_/Q vssd1 vssd1 vccd1 vccd1 _22766_/A sky130_fd_sc_hd__inv_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24504_ hold2599/X hold2571/X _24510_/S vssd1 vssd1 vccd1 vccd1 _24505_/A sky130_fd_sc_hd__mux2_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21716_ _21716_/A _21716_/B _21715_/X vssd1 vssd1 vccd1 vccd1 _21717_/B sky130_fd_sc_hd__or3b_1
X_25484_ _25495_/CLK hold881/X vssd1 vssd1 vccd1 vccd1 hold880/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22696_ _22697_/B _22697_/A vssd1 vssd1 vccd1 vccd1 _22698_/A sky130_fd_sc_hd__or2_1
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24435_ _24435_/A vssd1 vssd1 vccd1 vccd1 _26209_/D sky130_fd_sc_hd__clkbuf_1
X_21647_ _21647_/A _21647_/B vssd1 vssd1 vccd1 vccd1 _21648_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24366_ hold2241/X _26187_/Q _24433_/S vssd1 vssd1 vccd1 vccd1 _24366_/X sky130_fd_sc_hd__mux2_1
XANTENNA_70 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21578_ _21578_/A _21628_/B vssd1 vssd1 vccd1 vccd1 _21580_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26105_ _26231_/CLK _26105_/D vssd1 vssd1 vccd1 vccd1 _26105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23317_ _23317_/A hold896/X vssd1 vssd1 vccd1 vccd1 _23320_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_104_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20529_ _21579_/A vssd1 vssd1 vccd1 vccd1 _21578_/A sky130_fd_sc_hd__inv_2
X_24297_ _24297_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24298_/A sky130_fd_sc_hd__and2_1
XFILLER_0_104_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26036_ _26041_/CLK _26036_/D vssd1 vssd1 vccd1 vccd1 _26036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14050_ hold483/X _14049_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold484/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23248_ _24870_/B _23249_/A vssd1 vssd1 vccd1 vccd1 _23248_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13001_ _12930_/X _12999_/X _12917_/X _13000_/X vssd1 vssd1 vccd1 vccd1 _13001_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23179_ _23179_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _23179_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_0_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17740_ _17740_/A _17740_/B vssd1 vssd1 vccd1 vccd1 _17745_/B sky130_fd_sc_hd__nand2_1
X_14952_ _14965_/A _14964_/A vssd1 vssd1 vccd1 vccd1 _14952_/Y sky130_fd_sc_hd__nand2_1
X_13903_ _26282_/Q _13801_/X _13793_/X _13902_/Y vssd1 vssd1 vccd1 vccd1 _13904_/B
+ sky130_fd_sc_hd__a22o_1
X_17671_ _17671_/A _17671_/B vssd1 vssd1 vccd1 vccd1 _22075_/A sky130_fd_sc_hd__or2_1
X_14883_ _14881_/Y _14882_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14883_/Y sky130_fd_sc_hd__a21oi_1
X_19410_ _19452_/A _19410_/B vssd1 vssd1 vccd1 vccd1 _19410_/Y sky130_fd_sc_hd__nand2_1
X_16622_ _16698_/A hold887/X vssd1 vssd1 vccd1 vccd1 _16622_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_187_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13834_ _18853_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13834_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19341_ _26229_/Q _12537_/B hold849/X vssd1 vssd1 vccd1 vccd1 _19341_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16553_ _16555_/B vssd1 vssd1 vccd1 vccd1 _16575_/B sky130_fd_sc_hd__inv_2
XFILLER_0_168_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13765_ _13823_/A _13765_/B vssd1 vssd1 vccd1 vccd1 _13765_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_69_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15504_ _15502_/A _15481_/B _15496_/A vssd1 vssd1 vccd1 vccd1 _15504_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12716_ _12716_/A vssd1 vssd1 vccd1 vccd1 _24994_/D sky130_fd_sc_hd__clkbuf_1
X_19272_ _21203_/A vssd1 vssd1 vccd1 vccd1 _19272_/X sky130_fd_sc_hd__buf_12
X_16484_ _16482_/Y _16483_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 _16484_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13696_ _26249_/Q _13612_/X _13605_/X _13695_/Y vssd1 vssd1 vccd1 vccd1 _13697_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18223_ _18612_/A _18223_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18224_/C sky130_fd_sc_hd__nand3_1
X_12647_ _12654_/C _24980_/Q vssd1 vssd1 vccd1 vccd1 _12648_/A sky130_fd_sc_hd__nand2_1
X_15435_ _22848_/B _15435_/B vssd1 vssd1 vccd1 vccd1 _22845_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15366_ _15366_/A _15810_/B vssd1 vssd1 vccd1 vccd1 _15367_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_143_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18154_ _18529_/A _18156_/B vssd1 vssd1 vccd1 vccd1 _18155_/A sky130_fd_sc_hd__nand2_1
X_12578_ _12578_/A vssd1 vssd1 vccd1 vccd1 _23924_/A sky130_fd_sc_hd__inv_2
XFILLER_0_68_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17105_ _20322_/B _25885_/Q _25821_/Q vssd1 vssd1 vccd1 vccd1 _17106_/B sky130_fd_sc_hd__mux2_2
X_14317_ _14344_/A hold203/X vssd1 vssd1 vccd1 vccd1 hold204/A sky130_fd_sc_hd__nand2_1
X_15297_ _16781_/B vssd1 vssd1 vccd1 vccd1 _22709_/B sky130_fd_sc_hd__inv_2
XFILLER_0_29_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18085_ _18528_/A _25726_/Q vssd1 vssd1 vccd1 vccd1 _18087_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold307 hold307/A vssd1 vssd1 vccd1 vccd1 hold307/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 hold318/A vssd1 vssd1 vccd1 vccd1 hold318/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold329 hold329/A vssd1 vssd1 vccd1 vccd1 hold329/X sky130_fd_sc_hd__dlygate4sd3_1
X_17036_ _17917_/B _17036_/B vssd1 vssd1 vccd1 vccd1 _17623_/A sky130_fd_sc_hd__xor2_4
X_14248_ _14260_/A hold650/X vssd1 vssd1 vccd1 vccd1 hold651/A sky130_fd_sc_hd__nand2_1
XFILLER_0_159_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14179_ _26326_/Q _13518_/B _14170_/X _14178_/Y vssd1 vssd1 vccd1 vccd1 _14180_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ _18985_/Y _18986_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25695_/D sky130_fd_sc_hd__a21oi_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1007 _25093_/Q vssd1 vssd1 vccd1 vccd1 _18577_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17938_ _17938_/A _17938_/B vssd1 vssd1 vccd1 vccd1 _22159_/A sky130_fd_sc_hd__nand2_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1018 _12940_/X vssd1 vssd1 vccd1 vccd1 _25038_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1029 _25546_/Q vssd1 vssd1 vccd1 vccd1 _16750_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_79_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17869_ _19115_/B _25648_/Q vssd1 vssd1 vccd1 vccd1 _17873_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19608_ _19606_/X _19607_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19608_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20880_ _21235_/A _20880_/B vssd1 vssd1 vccd1 vccd1 _20880_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_177_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19539_ _19531_/X _19538_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19539_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22550_ _22550_/A _22550_/B vssd1 vssd1 vccd1 vccd1 _22551_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21501_ _21501_/A _21501_/B vssd1 vssd1 vccd1 vccd1 _21502_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_173_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22481_ _22481_/A _23001_/B _22481_/C vssd1 vssd1 vccd1 vccd1 _22481_/X sky130_fd_sc_hd__and3_1
XFILLER_0_12_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24220_ _24220_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24221_/A sky130_fd_sc_hd__and2_1
XFILLER_0_16_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21432_ _21432_/A _21432_/B _21432_/C vssd1 vssd1 vccd1 vccd1 _21436_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_146_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24151_ hold1955/X _26117_/Q _24203_/S vssd1 vssd1 vccd1 vccd1 _24151_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21363_ _21573_/A _21363_/B vssd1 vssd1 vccd1 vccd1 _21363_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23102_ _23100_/X _23101_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _23102_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20314_ _20314_/A _20314_/B _20314_/C vssd1 vssd1 vccd1 vccd1 _20318_/C sky130_fd_sc_hd__nand3_1
X_24082_ _24082_/A vssd1 vssd1 vccd1 vccd1 _26094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold830 hold830/A vssd1 vssd1 vccd1 vccd1 hold830/X sky130_fd_sc_hd__dlygate4sd3_1
X_21294_ _25876_/Q _21294_/B _21294_/C vssd1 vssd1 vccd1 vccd1 _21297_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold841 hold841/A vssd1 vssd1 vccd1 vccd1 hold841/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold852 hold852/A vssd1 vssd1 vccd1 vccd1 hold852/X sky130_fd_sc_hd__dlygate4sd3_1
X_23033_ _23033_/A _23193_/B _23033_/C vssd1 vssd1 vccd1 vccd1 _23033_/X sky130_fd_sc_hd__and3_1
Xhold863 hold863/A vssd1 vssd1 vccd1 vccd1 hold863/X sky130_fd_sc_hd__buf_1
X_20245_ _20245_/A _20245_/B vssd1 vssd1 vccd1 vccd1 _21466_/A sky130_fd_sc_hd__nand2_4
Xhold874 hold874/A vssd1 vssd1 vccd1 vccd1 hold874/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 hold885/A vssd1 vssd1 vccd1 vccd1 hold885/X sky130_fd_sc_hd__buf_1
Xhold896 hold896/A vssd1 vssd1 vccd1 vccd1 hold896/X sky130_fd_sc_hd__buf_1
X_20176_ _25842_/Q _20177_/A vssd1 vssd1 vccd1 vccd1 _20180_/A sky130_fd_sc_hd__or2_1
Xhold2220 _25997_/Q vssd1 vssd1 vccd1 vccd1 _14843_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2231 _14986_/Y vssd1 vssd1 vccd1 vccd1 hold2231/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2242 _24366_/X vssd1 vssd1 vccd1 vccd1 _24367_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2253 _26073_/Q vssd1 vssd1 vccd1 vccd1 hold2253/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24984_ _25422_/CLK _24984_/D vssd1 vssd1 vccd1 vccd1 _24984_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2264 _24228_/X vssd1 vssd1 vccd1 vccd1 _24229_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1530 _21445_/Y vssd1 vssd1 vccd1 vccd1 _25820_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2275 _24369_/X vssd1 vssd1 vccd1 vccd1 _24370_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2286 _26080_/Q vssd1 vssd1 vccd1 vccd1 hold2286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1541 _25814_/Q vssd1 vssd1 vccd1 vccd1 _21347_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2297 _15003_/Y vssd1 vssd1 vccd1 vccd1 hold2297/X sky130_fd_sc_hd__dlygate4sd3_1
X_23935_ hold2126/X _26047_/Q _24001_/S vssd1 vssd1 vccd1 vccd1 _23935_/X sky130_fd_sc_hd__mux2_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1552 _23018_/X vssd1 vssd1 vccd1 vccd1 _23019_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1563 _16707_/Y vssd1 vssd1 vccd1 vccd1 _25540_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1574 _25785_/Q vssd1 vssd1 vccd1 vccd1 _20464_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1585 _21526_/Y vssd1 vssd1 vccd1 vccd1 _25825_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23866_ _23866_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23867_/A sky130_fd_sc_hd__and2_1
Xhold1596 _25742_/Q vssd1 vssd1 vccd1 vccd1 _19582_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22817_ _22817_/A _23001_/B _22817_/C vssd1 vssd1 vccd1 vccd1 _22817_/X sky130_fd_sc_hd__and3_1
X_25605_ _26240_/CLK _25605_/D vssd1 vssd1 vccd1 vccd1 _25605_/Q sky130_fd_sc_hd__dfxtp_2
X_23797_ _14893_/B _26004_/Q _23831_/S vssd1 vssd1 vccd1 vccd1 _23797_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_183_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13550_ _17944_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13550_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_94_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25536_ _25537_/CLK hold943/X vssd1 vssd1 vccd1 vccd1 hold942/A sky130_fd_sc_hd__dfxtp_1
X_22748_ _15335_/B _22680_/X _14273_/X vssd1 vssd1 vccd1 vccd1 _22748_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xascon_wrapper_21 vssd1 vssd1 vccd1 vccd1 io_oeb[7] ascon_wrapper_21/LO sky130_fd_sc_hd__conb_1
XFILLER_0_183_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12501_ _19483_/A vssd1 vssd1 vccd1 vccd1 _12537_/B sky130_fd_sc_hd__buf_8
XFILLER_0_109_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25467_ _26069_/CLK _25467_/D vssd1 vssd1 vccd1 vccd1 _25467_/Q sky130_fd_sc_hd__dfxtp_1
X_13481_ hold605/X vssd1 vssd1 vccd1 vccd1 _17877_/B sky130_fd_sc_hd__inv_2
XFILLER_0_82_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22679_ _23188_/A _22679_/B vssd1 vssd1 vccd1 vccd1 _22679_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15220_ _15268_/C _15199_/B _15214_/A vssd1 vssd1 vccd1 vccd1 _15220_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_165_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24418_ hold2222/X _26204_/Q _24433_/S vssd1 vssd1 vccd1 vccd1 _24418_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_180_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25398_ _25425_/CLK _25398_/D vssd1 vssd1 vccd1 vccd1 _25398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15151_ _16729_/B vssd1 vssd1 vccd1 vccd1 _22504_/B sky130_fd_sc_hd__inv_2
X_24349_ _24349_/A vssd1 vssd1 vccd1 vccd1 _26181_/D sky130_fd_sc_hd__clkbuf_1
X_14102_ _18430_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14102_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_121_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15082_ _15083_/B _15083_/A vssd1 vssd1 vccd1 vccd1 _15084_/A sky130_fd_sc_hd__or2_1
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26019_ _26032_/CLK _26019_/D vssd1 vssd1 vccd1 vccd1 _26019_/Q sky130_fd_sc_hd__dfxtp_1
X_14033_ _25800_/Q vssd1 vssd1 vccd1 vccd1 _18203_/B sky130_fd_sc_hd__inv_2
X_18910_ _18951_/A _18914_/B vssd1 vssd1 vccd1 vccd1 _18912_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19890_ _19883_/X _19889_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19890_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18841_ _18841_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18841_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18772_ _18954_/A _25764_/Q vssd1 vssd1 vccd1 vccd1 _18774_/A sky130_fd_sc_hd__nand2_1
X_15984_ _15985_/B _15985_/A vssd1 vssd1 vccd1 vccd1 _15986_/A sky130_fd_sc_hd__or2_1
XFILLER_0_175_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17723_ _17723_/A _17723_/B vssd1 vssd1 vccd1 vccd1 _17727_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_145_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14935_ _14948_/A _14947_/A vssd1 vssd1 vccd1 vccd1 _14935_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_188_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17654_ _17652_/X _17528_/X _17653_/X vssd1 vssd1 vccd1 vccd1 _17655_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_188_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14866_ _14893_/A _14866_/B vssd1 vssd1 vccd1 vccd1 _22323_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16605_ _16605_/A _16691_/B vssd1 vssd1 vccd1 vccd1 _16608_/A sky130_fd_sc_hd__nand2_1
X_13817_ _13823_/A _13817_/B vssd1 vssd1 vccd1 vccd1 _13817_/Y sky130_fd_sc_hd__nand2_1
X_17585_ _17585_/A _17637_/A vssd1 vssd1 vccd1 vccd1 _17586_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14797_ _15839_/A _14797_/B vssd1 vssd1 vccd1 vccd1 _22091_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_161_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19324_ _19316_/X _19323_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19324_/Y sky130_fd_sc_hd__o21ai_1
X_16536_ _16537_/A _16537_/B _16541_/B vssd1 vssd1 vccd1 vccd1 _16536_/X sky130_fd_sc_hd__a21o_1
X_13748_ _13760_/A hold524/X vssd1 vssd1 vccd1 vccd1 hold525/A sky130_fd_sc_hd__nand2_1
XFILLER_0_156_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19255_ _19452_/A hold891/X vssd1 vssd1 vccd1 vccd1 hold892/A sky130_fd_sc_hd__nand2_1
X_16467_ _16492_/A _16467_/B vssd1 vssd1 vccd1 vccd1 _16486_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_57_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13679_ _14345_/A vssd1 vssd1 vccd1 vccd1 _13679_/X sky130_fd_sc_hd__buf_6
XFILLER_0_171_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18206_ _18413_/A _18555_/A vssd1 vssd1 vccd1 vccd1 _18207_/B sky130_fd_sc_hd__xnor2_1
X_15418_ _26022_/Q _25958_/Q _15773_/S vssd1 vssd1 vccd1 vccd1 _15419_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_5_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19186_ _19186_/A hold818/X vssd1 vssd1 vccd1 vccd1 hold819/A sky130_fd_sc_hd__nand2_1
X_16398_ _16396_/X hold519/X _16343_/X vssd1 vssd1 vccd1 vccd1 hold520/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18137_ _18954_/A _25734_/Q vssd1 vssd1 vccd1 vccd1 _18139_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_182_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15349_ _26018_/Q _25954_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15350_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_26_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold104 hold104/A vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold115 hold115/A vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold126 hold126/A vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
X_18068_ _18118_/B _17775_/C _17775_/A vssd1 vssd1 vccd1 vccd1 _18071_/A sky130_fd_sc_hd__a21o_1
Xhold137 hold137/A vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 hold148/A vssd1 vssd1 vccd1 vccd1 hold148/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold159 hold159/A vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
X_17019_ _20067_/B _25839_/Q _25775_/Q vssd1 vssd1 vccd1 vccd1 _17020_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_112_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20030_ _21677_/A _21370_/A vssd1 vssd1 vccd1 vccd1 _20031_/C sky130_fd_sc_hd__nand2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21981_ _25809_/Q _21981_/B vssd1 vssd1 vccd1 vccd1 _21981_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23720_ hold2079/X hold2049/X _23754_/S vssd1 vssd1 vccd1 vccd1 _23721_/A sky130_fd_sc_hd__mux2_1
X_20932_ _20932_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _20932_/Y sky130_fd_sc_hd__nand2_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23651_ _23651_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23652_/A sky130_fd_sc_hd__and2_1
X_20863_ _20862_/B _20863_/B _20863_/C vssd1 vssd1 vccd1 vccd1 _20864_/B sky130_fd_sc_hd__nand3b_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22602_ _22602_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _22602_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23582_ _25927_/Q _25926_/Q hold896/X _25924_/Q vssd1 vssd1 vccd1 vccd1 _23587_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_0_9_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20794_ _23133_/B vssd1 vssd1 vccd1 vccd1 _22620_/B sky130_fd_sc_hd__inv_2
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25321_ _26252_/CLK hold199/X vssd1 vssd1 vccd1 vccd1 hold197/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22533_ _22533_/A _22900_/B vssd1 vssd1 vccd1 vccd1 _22533_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_119_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25252_ _25257_/CLK hold385/X vssd1 vssd1 vccd1 vccd1 hold383/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22464_ _18756_/A _25827_/Q _22462_/Y _22463_/Y vssd1 vssd1 vccd1 vccd1 _22465_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24203_ hold1930/X _26134_/Q _24203_/S vssd1 vssd1 vccd1 vccd1 _24203_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21415_ _21465_/A _21418_/A vssd1 vssd1 vccd1 vccd1 _21416_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25183_ _26273_/CLK hold619/X vssd1 vssd1 vccd1 vccd1 hold617/A sky130_fd_sc_hd__dfxtp_1
X_22395_ _22396_/B _22396_/A vssd1 vssd1 vccd1 vccd1 _22397_/A sky130_fd_sc_hd__or2_1
X_24134_ _24134_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24135_/A sky130_fd_sc_hd__and2_1
X_21346_ _21346_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21346_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24065_ hold2134/X hold1911/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24066_/A sky130_fd_sc_hd__mux2_1
X_21277_ _21646_/B _21694_/B vssd1 vssd1 vccd1 vccd1 _21279_/A sky130_fd_sc_hd__nand2_1
Xhold660 hold660/A vssd1 vssd1 vccd1 vccd1 hold660/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 hold671/A vssd1 vssd1 vccd1 vccd1 hold671/X sky130_fd_sc_hd__buf_1
XFILLER_0_60_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23016_ _23015_/A _22849_/X _23015_/B vssd1 vssd1 vccd1 vccd1 _23017_/C sky130_fd_sc_hd__o21ai_1
Xhold682 hold682/A vssd1 vssd1 vccd1 vccd1 hold682/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 hold693/A vssd1 vssd1 vccd1 vccd1 hold693/X sky130_fd_sc_hd__dlygate4sd3_1
X_20228_ _26282_/Q hold611/X vssd1 vssd1 vccd1 vccd1 _20228_/Y sky130_fd_sc_hd__nand2_1
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20159_ _20159_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _20159_/Y sky130_fd_sc_hd__nand2_1
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2050 _23723_/X vssd1 vssd1 vccd1 vccd1 _23725_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2061 _26036_/Q vssd1 vssd1 vccd1 vccd1 hold2061/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2072 _25971_/Q vssd1 vssd1 vccd1 vccd1 hold2072/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2083 _23310_/Y vssd1 vssd1 vccd1 vccd1 _23311_/C sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _12930_/X _12978_/X _12917_/X _12980_/X vssd1 vssd1 vccd1 vccd1 _12981_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2094 _25951_/Q vssd1 vssd1 vccd1 vccd1 hold2094/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24967_ _25378_/CLK _24967_/D vssd1 vssd1 vccd1 vccd1 _24967_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1360 _13252_/X vssd1 vssd1 vccd1 vccd1 _25094_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ _14720_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14720_/Y sky130_fd_sc_hd__nand2_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1371 _25099_/Q vssd1 vssd1 vccd1 vccd1 _18699_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1382 _15783_/B vssd1 vssd1 vccd1 vccd1 _15784_/A sky130_fd_sc_hd__dlygate4sd3_1
X_23918_ _23918_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23919_/A sky130_fd_sc_hd__and2_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1393 _25767_/Q vssd1 vssd1 vccd1 vccd1 _19931_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24898_ _24896_/X _24897_/X _24957_/S vssd1 vssd1 vccd1 vccd1 _24898_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_169_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14651_ _14651_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _14651_/Y sky130_fd_sc_hd__nand2_1
X_23849_ _23849_/A vssd1 vssd1 vccd1 vccd1 _26020_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _13703_/A _13602_/B vssd1 vssd1 vccd1 vccd1 _13602_/Y sky130_fd_sc_hd__nand2_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _19518_/A _17370_/B vssd1 vssd1 vccd1 vccd1 _17607_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_170_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14582_ _14585_/A hold92/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16321_ _16321_/A _16321_/B vssd1 vssd1 vccd1 vccd1 _16336_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_82_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25519_ _25535_/CLK hold934/X vssd1 vssd1 vccd1 vccd1 hold933/A sky130_fd_sc_hd__dfxtp_1
X_13533_ _26223_/Q _13426_/X _13468_/X _13532_/Y vssd1 vssd1 vccd1 vccd1 _13534_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19040_ _19082_/A _19040_/B _22786_/A vssd1 vssd1 vccd1 vccd1 _19040_/X sky130_fd_sc_hd__and3_1
X_16252_ _16252_/A _16252_/B vssd1 vssd1 vccd1 vccd1 _16254_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_180_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13464_ _13944_/A vssd1 vssd1 vccd1 vccd1 _13583_/A sky130_fd_sc_hd__buf_8
XFILLER_0_164_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15203_ _15201_/Y _15202_/Y _15090_/X vssd1 vssd1 vccd1 vccd1 hold928/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16183_ _16189_/A _16184_/A vssd1 vssd1 vccd1 vccd1 _16183_/X sky130_fd_sc_hd__or2_1
X_13395_ _13395_/A vssd1 vssd1 vccd1 vccd1 _19774_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15134_ _16722_/B vssd1 vssd1 vccd1 vccd1 _22479_/B sky130_fd_sc_hd__inv_2
XFILLER_0_65_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15065_ _15065_/A _15065_/B vssd1 vssd1 vccd1 vccd1 _15066_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_121_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19942_ _19975_/A _19942_/B vssd1 vssd1 vccd1 vccd1 _19942_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_49_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14016_ _18102_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14016_/Y sky130_fd_sc_hd__nor2_1
X_19873_ _19948_/A _19888_/B vssd1 vssd1 vccd1 vccd1 _19875_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18824_ _19844_/A vssd1 vssd1 vccd1 vccd1 _22564_/B sky130_fd_sc_hd__inv_2
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18755_ _20566_/B _22465_/A vssd1 vssd1 vccd1 vccd1 _20557_/A sky130_fd_sc_hd__nand2_2
X_15967_ _15964_/X _15966_/Y _15805_/X vssd1 vssd1 vccd1 vccd1 hold930/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_164_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17706_ _17706_/A vssd1 vssd1 vccd1 vccd1 _17711_/A sky130_fd_sc_hd__clkinvlp_2
X_14918_ _14919_/B _14919_/A vssd1 vssd1 vccd1 vccd1 _14920_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18686_ _20439_/B _19744_/A vssd1 vssd1 vccd1 vccd1 _18687_/B sky130_fd_sc_hd__nand2_1
X_15898_ _16274_/A _15942_/B _15897_/X vssd1 vssd1 vccd1 vccd1 _15900_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_76_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17637_ _17637_/A _17637_/B vssd1 vssd1 vccd1 vccd1 _17638_/B sky130_fd_sc_hd__xnor2_1
X_14849_ _14842_/Y _14848_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14849_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17568_ _17568_/A vssd1 vssd1 vccd1 vccd1 _17568_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_147_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19307_ _19308_/B _19308_/A vssd1 vssd1 vccd1 vccd1 _19307_/X sky130_fd_sc_hd__or2_1
X_16519_ hold864/X vssd1 vssd1 vccd1 vccd1 _16522_/B sky130_fd_sc_hd__inv_2
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17499_ _17499_/A _17499_/B vssd1 vssd1 vccd1 vccd1 _17499_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19238_ _26221_/Q _19483_/A hold843/X vssd1 vssd1 vccd1 vccd1 _19239_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_128_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19169_ _19157_/X _19168_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19169_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_182_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21200_ _21200_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _21206_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_182_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22180_ _18532_/A _25816_/Q _22178_/Y _22179_/Y vssd1 vssd1 vccd1 vccd1 _22181_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21131_ _21131_/A _25870_/Q vssd1 vssd1 vccd1 vccd1 _21136_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21062_ _21062_/A _21062_/B _21062_/C vssd1 vssd1 vccd1 vccd1 _21063_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_10_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20013_ _20013_/A _25877_/Q vssd1 vssd1 vccd1 vccd1 _20018_/A sky130_fd_sc_hd__nand2_1
X_25870_ _25875_/CLK _25870_/D vssd1 vssd1 vccd1 vccd1 _25870_/Q sky130_fd_sc_hd__dfxtp_4
X_24821_ _24821_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24822_/A sky130_fd_sc_hd__and2_1
X_21964_ _21936_/X _21963_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _21964_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24752_ _24752_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24753_/A sky130_fd_sc_hd__and2_1
XFILLER_0_94_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23703_ _23703_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23704_/A sky130_fd_sc_hd__and2_1
X_20915_ _20915_/A _20915_/B vssd1 vssd1 vccd1 vccd1 _20917_/A sky130_fd_sc_hd__nand2_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24683_ hold2495/X _26290_/Q _24740_/S vssd1 vssd1 vccd1 vccd1 _24683_/X sky130_fd_sc_hd__mux2_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21895_ _21867_/X _21894_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _21895_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23634_ _23634_/A vssd1 vssd1 vccd1 vccd1 _25950_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20846_ _20846_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _20851_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23565_ _23562_/Y _23564_/Y _24957_/S vssd1 vssd1 vccd1 vccd1 _23565_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20777_ _21235_/A _20777_/B vssd1 vssd1 vccd1 vccd1 _20777_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_119_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22516_ _19816_/A _22515_/A _22515_/Y vssd1 vssd1 vccd1 vccd1 _22518_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25304_ _26135_/CLK hold217/X vssd1 vssd1 vccd1 vccd1 hold215/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26284_ _26284_/CLK _26284_/D vssd1 vssd1 vccd1 vccd1 _26284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23496_ _23489_/X _23495_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _23496_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_146_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22447_ _23136_/A _22447_/B vssd1 vssd1 vccd1 vccd1 _22448_/A sky130_fd_sc_hd__xor2_1
X_25235_ _25689_/CLK hold759/X vssd1 vssd1 vccd1 vccd1 hold757/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13180_ _18373_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13180_/X sky130_fd_sc_hd__or2_1
X_25166_ _25779_/CLK hold667/X vssd1 vssd1 vccd1 vccd1 hold665/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22378_ _22808_/A _22957_/B vssd1 vssd1 vccd1 vccd1 _22381_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24117_ hold2512/X hold2451/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24118_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_32_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21329_ _21329_/A _21329_/B vssd1 vssd1 vccd1 vccd1 _21330_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_130_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25097_ _26184_/CLK _25097_/D vssd1 vssd1 vccd1 vccd1 _25097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24048_ _24048_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24049_/A sky130_fd_sc_hd__and2_1
Xhold490 hold490/A vssd1 vssd1 vccd1 vccd1 hold490/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16870_ _16868_/X _16711_/X _16869_/Y _25885_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16871_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_159_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15821_ _15819_/X hold2681/X _15805_/X vssd1 vssd1 vccd1 vccd1 _15821_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25999_ _25999_/CLK _25999_/D vssd1 vssd1 vccd1 vccd1 _25999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18540_ _18537_/Y _18538_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25671_/D sky130_fd_sc_hd__a21oi_1
X_15752_ _15752_/A vssd1 vssd1 vccd1 vccd1 _15761_/B sky130_fd_sc_hd__inv_2
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _17493_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12964_/X sky130_fd_sc_hd__or2_1
XFILLER_0_172_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1190 _16950_/Y vssd1 vssd1 vccd1 vccd1 _25575_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ _14900_/A _14703_/B vssd1 vssd1 vccd1 vccd1 _14703_/Y sky130_fd_sc_hd__nand2_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18471_ _20018_/C _22097_/A vssd1 vssd1 vccd1 vccd1 _20010_/A sky130_fd_sc_hd__nand2_2
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ _15683_/A _15774_/B vssd1 vssd1 vccd1 vccd1 _15684_/B sky130_fd_sc_hd__nand2_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _17383_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12895_/X sky130_fd_sc_hd__or2_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _17594_/A _17644_/B vssd1 vssd1 vccd1 vccd1 _17423_/B sky130_fd_sc_hd__xnor2_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ _14632_/Y hold144/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold145/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _17393_/A _17353_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17353_/X sky130_fd_sc_hd__and3_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14565_ _14563_/Y hold162/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold163/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16304_ _16304_/A _16691_/B vssd1 vssd1 vccd1 vccd1 _16306_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_165_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13516_ _13522_/A hold843/X vssd1 vssd1 vccd1 vccd1 _13516_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17284_ _17284_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17284_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14496_ _14494_/Y hold111/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold112/A sky130_fd_sc_hd__a21oi_1
X_19023_ _19021_/Y _19022_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25700_/D sky130_fd_sc_hd__a21oi_1
X_16235_ _16235_/A hold972/X _16401_/C vssd1 vssd1 vccd1 vccd1 _16236_/B sky130_fd_sc_hd__and3_1
XFILLER_0_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13447_ _13522_/A _13445_/X _23629_/B _13446_/X vssd1 vssd1 vccd1 vccd1 _13447_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16166_ _16168_/B _16168_/A vssd1 vssd1 vccd1 vccd1 _16167_/A sky130_fd_sc_hd__nor2_1
X_13378_ _26326_/Q _19729_/A vssd1 vssd1 vccd1 vccd1 _14644_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15117_ _15810_/B vssd1 vssd1 vccd1 vccd1 _15812_/B sky130_fd_sc_hd__buf_8
XFILLER_0_140_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16097_ _16097_/A _16097_/B vssd1 vssd1 vccd1 vccd1 _16099_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15048_ _15049_/B _15049_/A vssd1 vssd1 vccd1 vccd1 _15050_/A sky130_fd_sc_hd__or2_1
X_19925_ _20087_/A _18949_/A _20092_/C vssd1 vssd1 vccd1 vccd1 _19989_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_167_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19856_ _26265_/Q _19134_/X hold733/X vssd1 vssd1 vccd1 vccd1 _19857_/C sky130_fd_sc_hd__a21o_1
X_18807_ _18807_/A _18807_/B vssd1 vssd1 vccd1 vccd1 _22538_/A sky130_fd_sc_hd__nand2_1
X_19787_ _19784_/Y _19787_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19787_/X sky130_fd_sc_hd__and3b_1
X_16999_ _21716_/A vssd1 vssd1 vccd1 vccd1 _21042_/A sky130_fd_sc_hd__buf_12
X_18738_ _18738_/A _18738_/B vssd1 vssd1 vccd1 vccd1 _18738_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_183_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18669_ _18951_/A _18673_/B vssd1 vssd1 vccd1 vccd1 _18671_/A sky130_fd_sc_hd__nand2_1
X_20700_ _20697_/Y _20699_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _20700_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21680_ _21680_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _21685_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_114_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20631_ _20630_/B _20631_/B _20631_/C vssd1 vssd1 vccd1 vccd1 _20632_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_110_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23350_ _23351_/B _23351_/A vssd1 vssd1 vccd1 vccd1 _23350_/X sky130_fd_sc_hd__or2_1
XFILLER_0_144_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20562_ _20562_/A _22468_/B _20562_/C vssd1 vssd1 vccd1 vccd1 _20566_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22301_ _22302_/B _22302_/A vssd1 vssd1 vccd1 vccd1 _22303_/A sky130_fd_sc_hd__or2_1
X_23281_ hold832/X _23284_/A vssd1 vssd1 vccd1 vccd1 _23281_/X sky130_fd_sc_hd__or2_1
XFILLER_0_117_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20493_ _21276_/C _21562_/A vssd1 vssd1 vccd1 vccd1 _20495_/A sky130_fd_sc_hd__nand2_1
X_25020_ _26231_/CLK _25020_/D vssd1 vssd1 vccd1 vccd1 _25020_/Q sky130_fd_sc_hd__dfxtp_1
X_22232_ _22653_/A _22232_/B vssd1 vssd1 vccd1 vccd1 _22232_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22163_ _19216_/A _22162_/A _22162_/Y vssd1 vssd1 vccd1 vccd1 _22165_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21114_ _21114_/A _21114_/B _21114_/C vssd1 vssd1 vccd1 vccd1 _21118_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_100_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22094_ _22094_/A _25877_/Q vssd1 vssd1 vccd1 vccd1 _22094_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25922_ _25925_/CLK _25922_/D vssd1 vssd1 vccd1 vccd1 _25922_/Q sky130_fd_sc_hd__dfxtp_1
X_21045_ _21235_/A _21045_/B vssd1 vssd1 vccd1 vccd1 _21045_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25853_ _26207_/CLK _25853_/D vssd1 vssd1 vccd1 vccd1 _25853_/Q sky130_fd_sc_hd__dfxtp_4
X_24804_ _24804_/A vssd1 vssd1 vccd1 vccd1 _26329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25784_ _25784_/CLK _25784_/D vssd1 vssd1 vccd1 vccd1 _25784_/Q sky130_fd_sc_hd__dfxtp_1
X_22996_ _23188_/A _22996_/B vssd1 vssd1 vccd1 vccd1 _22996_/X sky130_fd_sc_hd__or2_1
XFILLER_0_119_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24735_ _24735_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24736_/A sky130_fd_sc_hd__and2_1
XFILLER_0_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21947_ _25808_/Q _21947_/B vssd1 vssd1 vccd1 vccd1 _21947_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_97_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12680_ _12680_/A _12684_/A vssd1 vssd1 vccd1 vccd1 _12680_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_139_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24666_ _24666_/A vssd1 vssd1 vccd1 vccd1 _26284_/D sky130_fd_sc_hd__clkbuf_1
X_21878_ _25806_/Q _21878_/B vssd1 vssd1 vccd1 vccd1 _21878_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_132_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23617_ _23617_/A _23629_/B vssd1 vssd1 vccd1 vccd1 _23618_/A sky130_fd_sc_hd__and2_1
X_20829_ _20829_/A _20829_/B vssd1 vssd1 vccd1 vccd1 _20833_/A sky130_fd_sc_hd__nand2_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24597_ hold2738/X hold2329/X _24664_/S vssd1 vssd1 vccd1 vccd1 _24598_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_107_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26336_ _26336_/CLK _26336_/D vssd1 vssd1 vccd1 vccd1 _26336_/Q sky130_fd_sc_hd__dfxtp_2
X_14350_ _14404_/A hold26/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__nand2_1
X_23548_ _23545_/Y _23547_/Y _24858_/S vssd1 vssd1 vccd1 vccd1 _23548_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_135_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13301_ _18759_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13301_/X sky130_fd_sc_hd__or2_1
X_14281_ _14278_/X hold1941/X _14280_/X vssd1 vssd1 vccd1 vccd1 _14281_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23479_ _23476_/Y _23478_/Y _24946_/A vssd1 vssd1 vccd1 vccd1 _23479_/X sky130_fd_sc_hd__mux2_1
X_26267_ _26267_/CLK _26267_/D vssd1 vssd1 vccd1 vccd1 _26267_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_80_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16020_ hold662/X vssd1 vssd1 vccd1 vccd1 _16023_/B sky130_fd_sc_hd__inv_2
X_13232_ _13207_/X _13230_/X _13192_/X _13231_/X vssd1 vssd1 vccd1 vccd1 _13232_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25218_ _25797_/CLK hold637/X vssd1 vssd1 vccd1 vccd1 hold635/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26198_ _26198_/CLK _26198_/D vssd1 vssd1 vccd1 vccd1 _26198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13163_ _13109_/X _13161_/X _13096_/X _13162_/X vssd1 vssd1 vccd1 vccd1 _13163_/X
+ sky130_fd_sc_hd__o211a_1
X_25149_ _26226_/CLK hold592/X vssd1 vssd1 vccd1 vccd1 hold590/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13094_ _13049_/X _14497_/A _13067_/X _25648_/Q vssd1 vssd1 vccd1 vccd1 _13094_/X
+ sky130_fd_sc_hd__a22o_1
X_17971_ _25842_/Q _17971_/B _17971_/C vssd1 vssd1 vccd1 vccd1 _17978_/A sky130_fd_sc_hd__and3b_2
X_19710_ _19708_/Y _19709_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19710_/Y sky130_fd_sc_hd__a21oi_1
X_16922_ _16923_/B _16923_/A vssd1 vssd1 vccd1 vccd1 _16922_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19641_ _26250_/Q hold572/X vssd1 vssd1 vccd1 vccd1 _19641_/Y sky130_fd_sc_hd__nand2_1
X_16853_ _16935_/A _16858_/B vssd1 vssd1 vccd1 vccd1 _16855_/B sky130_fd_sc_hd__nand2_1
X_15804_ _23245_/A vssd1 vssd1 vccd1 vccd1 _17568_/A sky130_fd_sc_hd__buf_6
XFILLER_0_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19572_ _19571_/Y _19272_/X _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19573_/B
+ sky130_fd_sc_hd__a211o_1
X_16784_ _22709_/B _16977_/A _16780_/Y _16783_/Y _12702_/A vssd1 vssd1 vccd1 vccd1
+ _16784_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_0_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13996_ _17958_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13996_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_87_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18523_ _18523_/A _18523_/B vssd1 vssd1 vccd1 vccd1 _22178_/A sky130_fd_sc_hd__nand2_1
X_15735_ _15733_/Y _15734_/Y _15464_/X vssd1 vssd1 vccd1 vccd1 hold884/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ _12891_/X _14409_/A _12909_/X _25620_/Q vssd1 vssd1 vccd1 vccd1 _12947_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18454_ _18454_/A _18454_/B vssd1 vssd1 vccd1 vccd1 _18454_/X sky130_fd_sc_hd__xor2_1
X_15666_ _26036_/Q _25972_/Q _15773_/S vssd1 vssd1 vccd1 vccd1 _15667_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_87_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _26110_/Q _12748_/X _12877_/X vssd1 vssd1 vccd1 vccd1 _12878_/X sky130_fd_sc_hd__a21o_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ _17402_/X _17241_/X _17404_/X vssd1 vssd1 vccd1 vccd1 _17406_/A sky130_fd_sc_hd__a21o_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14617_ _14617_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14617_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_173_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18385_ _18385_/A _25809_/Q _18385_/C vssd1 vssd1 vccd1 vccd1 _21216_/B sky130_fd_sc_hd__nand3_2
X_15597_ _15597_/A _15776_/B vssd1 vssd1 vccd1 vccd1 _15598_/B sky130_fd_sc_hd__nand2_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17336_ _17467_/A _17336_/B vssd1 vssd1 vccd1 vccd1 _17336_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_173_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14548_ _14548_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14548_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_83_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17267_ _17542_/A _17622_/A vssd1 vssd1 vccd1 vccd1 _17268_/B sky130_fd_sc_hd__xnor2_2
X_14479_ _14479_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14479_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_148_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19006_ _19004_/X _18879_/X _19005_/X vssd1 vssd1 vccd1 vccd1 _19007_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_102_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16218_ _16208_/B _16214_/B _16188_/Y _16217_/Y _16206_/B vssd1 vssd1 vccd1 vccd1
+ _16276_/A sky130_fd_sc_hd__o221ai_4
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17198_ _17506_/A _17585_/A vssd1 vssd1 vccd1 vccd1 _17199_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16149_ _16149_/A _16149_/B vssd1 vssd1 vccd1 vccd1 _16156_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2605 _24748_/X vssd1 vssd1 vccd1 vccd1 _24749_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2616 _24606_/X vssd1 vssd1 vccd1 vccd1 _24607_/A sky130_fd_sc_hd__dlygate4sd3_1
X_19908_ _26269_/Q _19134_/X hold803/X vssd1 vssd1 vccd1 vccd1 _19909_/C sky130_fd_sc_hd__a21o_1
Xhold2627 _24535_/X vssd1 vssd1 vccd1 vccd1 _24536_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2638 _26293_/Q vssd1 vssd1 vccd1 vccd1 hold2638/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2649 _25441_/Q vssd1 vssd1 vccd1 vccd1 _15204_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1904 _23681_/X vssd1 vssd1 vccd1 vccd1 _23682_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1915 _25913_/Q vssd1 vssd1 vccd1 vccd1 _23254_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1926 _25950_/Q vssd1 vssd1 vccd1 vccd1 hold1926/X sky130_fd_sc_hd__dlygate4sd3_1
X_19839_ _19837_/Y _19838_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19839_/Y sky130_fd_sc_hd__a21oi_1
Xhold1937 _23662_/X vssd1 vssd1 vccd1 vccd1 _23663_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1948 _24971_/Q vssd1 vssd1 vccd1 vccd1 _12503_/A sky130_fd_sc_hd__buf_1
Xhold1959 _26305_/Q vssd1 vssd1 vccd1 vccd1 hold1959/X sky130_fd_sc_hd__dlygate4sd3_1
X_22850_ _22848_/A _22849_/X _22848_/B vssd1 vssd1 vccd1 vccd1 _22851_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21801_ _25795_/Q _21801_/B vssd1 vssd1 vccd1 vccd1 _21801_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_91_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22781_ _26059_/Q vssd1 vssd1 vccd1 vccd1 _22782_/A sky130_fd_sc_hd__inv_2
XFILLER_0_151_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24520_ hold1999/X _26237_/Q _24587_/S vssd1 vssd1 vccd1 vccd1 _24520_/X sky130_fd_sc_hd__mux2_1
X_21732_ _19303_/A _21731_/A _21731_/Y vssd1 vssd1 vccd1 vccd1 _21734_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24451_ _24451_/A vssd1 vssd1 vccd1 vccd1 _26214_/D sky130_fd_sc_hd__clkbuf_1
X_21663_ _21663_/A _21663_/B vssd1 vssd1 vccd1 vccd1 _21664_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_143_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23402_ _24942_/S hold335/A _23401_/X vssd1 vssd1 vccd1 vccd1 _23402_/Y sky130_fd_sc_hd__o21ai_1
X_20614_ _20614_/A _20614_/B vssd1 vssd1 vccd1 vccd1 _20615_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24382_ hold2331/X hold2269/X _24433_/S vssd1 vssd1 vccd1 vccd1 _24383_/A sky130_fd_sc_hd__mux2_1
X_21594_ _21594_/A _21594_/B _21594_/C vssd1 vssd1 vccd1 vccd1 _21598_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23333_ hold952/X _23334_/A vssd1 vssd1 vccd1 vccd1 _23333_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26121_ _26121_/CLK _26121_/D vssd1 vssd1 vccd1 vccd1 _26121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20545_ _20543_/Y _20544_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _20545_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_140_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _25803_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_172_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23264_ _23264_/A hold875/X vssd1 vssd1 vccd1 vccd1 hold876/A sky130_fd_sc_hd__nand2_1
X_26052_ _26052_/CLK _26052_/D vssd1 vssd1 vccd1 vccd1 _26052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20476_ _20476_/A _20476_/B vssd1 vssd1 vccd1 vccd1 _21279_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_85_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22215_ _22858_/B vssd1 vssd1 vccd1 vccd1 _22859_/A sky130_fd_sc_hd__inv_2
X_25003_ _26121_/CLK _25003_/D vssd1 vssd1 vccd1 vccd1 _25003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23195_ _23195_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _23195_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_131_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22146_ _22144_/X _15839_/B _22145_/Y _14822_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _22147_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_125_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22077_ _17803_/A _25784_/Q _22075_/Y _22076_/Y vssd1 vssd1 vccd1 vccd1 _22078_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25905_ _26269_/CLK _25905_/D vssd1 vssd1 vccd1 vccd1 _25905_/Q sky130_fd_sc_hd__dfxtp_1
X_21028_ _21027_/B _21028_/B _21028_/C vssd1 vssd1 vccd1 vccd1 _21029_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_96_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25836_ _25838_/CLK _25836_/D vssd1 vssd1 vccd1 vccd1 _25836_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13850_ _13880_/A hold680/X vssd1 vssd1 vccd1 vccd1 hold681/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12801_ _17161_/B _14264_/A vssd1 vssd1 vccd1 vccd1 _12801_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13781_ _25760_/Q vssd1 vssd1 vccd1 vccd1 _18693_/B sky130_fd_sc_hd__inv_2
X_25767_ _25770_/CLK _25767_/D vssd1 vssd1 vccd1 vccd1 _25767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22979_ _23188_/A _22979_/B vssd1 vssd1 vccd1 vccd1 _22979_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15520_ _15518_/Y _15519_/Y _15464_/X vssd1 vssd1 vccd1 vccd1 hold879/A sky130_fd_sc_hd__a21oi_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _15543_/B vssd1 vssd1 vccd1 vccd1 _16711_/A sky130_fd_sc_hd__clkbuf_16
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24718_ _24718_/A vssd1 vssd1 vccd1 vccd1 _26301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25698_ _26334_/CLK _25698_/D vssd1 vssd1 vccd1 vccd1 _25698_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _16842_/B vssd1 vssd1 vccd1 vccd1 _22866_/B sky130_fd_sc_hd__inv_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12663_ _12663_/A vssd1 vssd1 vccd1 vccd1 _24984_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24649_ _24649_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24650_/A sky130_fd_sc_hd__and2_1
XFILLER_0_155_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _14400_/Y hold201/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold202/A sky130_fd_sc_hd__a21oi_1
X_18170_ _18170_/A _20962_/B _18170_/C vssd1 vssd1 vccd1 vccd1 _20944_/B sky130_fd_sc_hd__nand3_2
X_15382_ _26020_/Q _25956_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15383_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_136_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12594_ _12594_/A vssd1 vssd1 vccd1 vccd1 _12644_/B sky130_fd_sc_hd__inv_2
XFILLER_0_136_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17121_ _17402_/A _17121_/B vssd1 vssd1 vccd1 vccd1 _17121_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_182_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14333_ _14331_/Y hold336/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold337/A sky130_fd_sc_hd__a21oi_1
X_26319_ _26325_/CLK _26319_/D vssd1 vssd1 vccd1 vccd1 _26319_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_53_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_131_clk clkbuf_leaf_82_clk/A vssd1 vssd1 vccd1 vccd1 _25249_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_151_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17052_ _17966_/B _17052_/B vssd1 vssd1 vccd1 vccd1 _17630_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_162_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14264_ _14264_/A _14264_/B vssd1 vssd1 vccd1 vccd1 _14264_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16003_ _15975_/A _16054_/C _16002_/Y vssd1 vssd1 vccd1 vccd1 _16056_/B sky130_fd_sc_hd__a21o_1
X_13215_ _26300_/Q _19359_/A vssd1 vssd1 vccd1 vccd1 _14563_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_122_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14195_ _25826_/Q vssd1 vssd1 vccd1 vccd1 _18734_/B sky130_fd_sc_hd__inv_2
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13146_ _13146_/A vssd1 vssd1 vccd1 vccd1 _19206_/A sky130_fd_sc_hd__buf_4
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17954_ _18612_/A _25730_/Q _18083_/C vssd1 vssd1 vccd1 vccd1 _17955_/C sky130_fd_sc_hd__nand3_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13077_ _26276_/Q _25645_/Q vssd1 vssd1 vccd1 vccd1 _14488_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16905_ _16903_/X _16711_/X _16904_/Y _23021_/B _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16905_/X sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_198_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _26240_/CLK sky130_fd_sc_hd__clkbuf_16
X_17885_ _19206_/A vssd1 vssd1 vccd1 vccd1 _22131_/B sky130_fd_sc_hd__inv_2
XFILLER_0_164_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16836_ _25880_/Q _13468_/X _16774_/Y vssd1 vssd1 vccd1 vccd1 _16836_/Y sky130_fd_sc_hd__a21oi_1
X_19624_ _19723_/A _19624_/B vssd1 vssd1 vccd1 vccd1 _19624_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19555_ _19553_/Y _19554_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19555_/Y sky130_fd_sc_hd__a21oi_1
X_16767_ _16768_/B _16768_/A vssd1 vssd1 vccd1 vccd1 _16767_/X sky130_fd_sc_hd__or2_1
XFILLER_0_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13979_ hold761/X _13978_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold762/A sky130_fd_sc_hd__a21oi_1
X_18506_ _18793_/A _25751_/Q _18891_/C vssd1 vssd1 vccd1 vccd1 _18507_/C sky130_fd_sc_hd__nand3_1
X_15718_ _15718_/A _15718_/B vssd1 vssd1 vccd1 vccd1 _15763_/A sky130_fd_sc_hd__nor2_1
X_19486_ _19485_/Y _19272_/X _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19487_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16698_ _16698_/A hold575/X vssd1 vssd1 vccd1 vccd1 hold576/A sky130_fd_sc_hd__nand2_1
XFILLER_0_119_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18437_ _18437_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18437_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_185_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15649_ _15649_/A _15774_/B vssd1 vssd1 vccd1 vccd1 _15650_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_146_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18368_ _18368_/A _18368_/B _18368_/C vssd1 vssd1 vccd1 vccd1 _21949_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_145_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17319_ _25709_/Q _17319_/B vssd1 vssd1 vccd1 vccd1 _17651_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18299_ _21844_/B _25613_/Q vssd1 vssd1 vccd1 vccd1 _18301_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_122_clk clkbuf_4_11__f_clk/X vssd1 vssd1 vccd1 vccd1 _26193_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20330_ _20330_/A _20330_/B _20330_/C vssd1 vssd1 vccd1 vccd1 _20331_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_109_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20261_ _20261_/A _20261_/B _21036_/B vssd1 vssd1 vccd1 vccd1 _20262_/B sky130_fd_sc_hd__nand3_1
X_22000_ _21998_/Y _21999_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _22000_/Y sky130_fd_sc_hd__a21oi_1
X_20192_ _21203_/A vssd1 vssd1 vccd1 vccd1 _20192_/X sky130_fd_sc_hd__buf_12
XFILLER_0_45_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2402 _26077_/Q vssd1 vssd1 vccd1 vccd1 hold2402/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2413 _25444_/Q vssd1 vssd1 vccd1 vccd1 _15261_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2424 _25689_/Q vssd1 vssd1 vccd1 vccd1 _13341_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2435 _26124_/Q vssd1 vssd1 vccd1 vccd1 hold2435/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2446 _24967_/Q vssd1 vssd1 vccd1 vccd1 _12567_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1701 _25788_/Q vssd1 vssd1 vccd1 vccd1 _20583_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2457 _25469_/Q vssd1 vssd1 vccd1 vccd1 _15703_/A sky130_fd_sc_hd__dlygate4sd3_1
X_23951_ _23951_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23952_/A sky130_fd_sc_hd__and2_1
Xhold1712 _21574_/Y vssd1 vssd1 vccd1 vccd1 _25828_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_189_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _26248_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1723 _25652_/Q vssd1 vssd1 vccd1 vccd1 _18110_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2468 _25684_/Q vssd1 vssd1 vccd1 vccd1 _13309_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1734 _25881_/Q vssd1 vssd1 vccd1 vccd1 _22872_/B sky130_fd_sc_hd__buf_1
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2479 _23995_/X vssd1 vssd1 vccd1 vccd1 _23996_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1745 _22716_/Y vssd1 vssd1 vccd1 vccd1 _25872_/D sky130_fd_sc_hd__dlygate4sd3_1
X_22902_ _22902_/A _22902_/B vssd1 vssd1 vccd1 vccd1 _22902_/Y sky130_fd_sc_hd__nand2_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1756 _25598_/Q vssd1 vssd1 vccd1 vccd1 _17246_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23882_ _23882_/A vssd1 vssd1 vccd1 vccd1 _26031_/D sky130_fd_sc_hd__clkbuf_1
Xhold1767 _22562_/Y vssd1 vssd1 vccd1 vccd1 _25866_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1778 _25868_/Q vssd1 vssd1 vccd1 vccd1 _22612_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1789 _25860_/Q vssd1 vssd1 vccd1 vccd1 _22405_/B sky130_fd_sc_hd__dlygate4sd3_1
X_25621_ _26122_/CLK _25621_/D vssd1 vssd1 vccd1 vccd1 _25621_/Q sky130_fd_sc_hd__dfxtp_4
X_22833_ _22832_/A _22454_/X _22832_/B vssd1 vssd1 vccd1 vccd1 _22834_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_168_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25552_ _25877_/CLK _25552_/D vssd1 vssd1 vccd1 vccd1 _25552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22764_ _15351_/B _22680_/X _14273_/X vssd1 vssd1 vccd1 vccd1 _22764_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24503_ _24503_/A vssd1 vssd1 vccd1 vccd1 _26231_/D sky130_fd_sc_hd__clkbuf_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21715_ _21714_/Y _21203_/X _20986_/A _20957_/A vssd1 vssd1 vccd1 vccd1 _21715_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25483_ _25483_/CLK hold445/X vssd1 vssd1 vccd1 vccd1 hold443/A sky130_fd_sc_hd__dfxtp_1
X_22695_ _25708_/Q _22694_/A _22694_/Y vssd1 vssd1 vccd1 vccd1 _22697_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24434_ _24434_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24435_/A sky130_fd_sc_hd__and2_1
X_21646_ _21646_/A _21646_/B _21646_/C vssd1 vssd1 vccd1 vccd1 _21647_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_47_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_113_clk clkbuf_4_14__f_clk/X vssd1 vssd1 vccd1 vccd1 _26207_/CLK sky130_fd_sc_hd__clkbuf_16
X_24365_ _24365_/A vssd1 vssd1 vccd1 vccd1 _26186_/D sky130_fd_sc_hd__clkbuf_1
X_21577_ _21577_/A _21577_/B _21577_/C vssd1 vssd1 vccd1 vccd1 _21581_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_133_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_60 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_71 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26104_ _26231_/CLK _26104_/D vssd1 vssd1 vccd1 vccd1 _26104_/Q sky130_fd_sc_hd__dfxtp_1
X_23316_ _23316_/A vssd1 vssd1 vccd1 vccd1 _23320_/B sky130_fd_sc_hd__inv_2
XFILLER_0_90_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20528_ _21302_/C _21579_/A vssd1 vssd1 vccd1 vccd1 _20531_/A sky130_fd_sc_hd__nand2_1
X_24296_ hold2171/X hold2077/X _24356_/S vssd1 vssd1 vccd1 vccd1 _24297_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26035_ _26041_/CLK _26035_/D vssd1 vssd1 vccd1 vccd1 _26035_/Q sky130_fd_sc_hd__dfxtp_1
X_23247_ _23254_/A vssd1 vssd1 vccd1 vccd1 _24870_/B sky130_fd_sc_hd__inv_2
XFILLER_0_127_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20459_ _26288_/Q hold485/X vssd1 vssd1 vccd1 vccd1 _20459_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13000_ _17543_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13000_/X sky130_fd_sc_hd__or2_1
X_23178_ _16977_/B _22421_/A _23172_/X _23173_/Y _23177_/X vssd1 vssd1 vccd1 vccd1
+ _23179_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_63_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22129_ _22626_/A _22807_/B vssd1 vssd1 vccd1 vccd1 _22139_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14951_ _14964_/A _14965_/A vssd1 vssd1 vccd1 vccd1 _14951_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13902_ _18022_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13902_/Y sky130_fd_sc_hd__nor2_1
X_17670_ _25592_/Q _22076_/B vssd1 vssd1 vccd1 vccd1 _17671_/B sky130_fd_sc_hd__nor2_1
X_14882_ _14900_/A _14882_/B vssd1 vssd1 vccd1 vccd1 _14882_/Y sky130_fd_sc_hd__nand2_1
X_16621_ _16619_/X _16620_/Y _16231_/A vssd1 vssd1 vccd1 vccd1 _16621_/X sky130_fd_sc_hd__a21o_1
X_13833_ _25768_/Q vssd1 vssd1 vccd1 vccd1 _18853_/B sky130_fd_sc_hd__inv_2
X_25819_ _25822_/CLK _25819_/D vssd1 vssd1 vccd1 vccd1 _25819_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19340_ _19338_/Y _19339_/Y _19086_/X vssd1 vssd1 vccd1 vccd1 _19340_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16552_ _16564_/B _16552_/B vssd1 vssd1 vccd1 vccd1 _16555_/B sky130_fd_sc_hd__and2_1
XFILLER_0_134_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13764_ _26260_/Q _13612_/X _13605_/X _13763_/Y vssd1 vssd1 vccd1 vccd1 _13765_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15503_ _15414_/A _15552_/A _15469_/Y vssd1 vssd1 vccd1 vccd1 _15503_/Y sky130_fd_sc_hd__a21oi_1
X_12715_ _12715_/A _24836_/B _12718_/A vssd1 vssd1 vccd1 vccd1 _12715_/X sky130_fd_sc_hd__and3_1
X_19271_ _26224_/Q hold458/X vssd1 vssd1 vccd1 vccd1 _19271_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_35_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16483_ _16698_/A _16483_/B vssd1 vssd1 vccd1 vccd1 _16483_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13695_ _18408_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13695_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_167_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18222_ _18611_/A _25737_/Q vssd1 vssd1 vccd1 vccd1 _18224_/A sky130_fd_sc_hd__nand2_1
X_15434_ _15434_/A _15776_/B vssd1 vssd1 vccd1 vccd1 _15435_/B sky130_fd_sc_hd__nand2_2
X_12646_ _12646_/A _12646_/B vssd1 vssd1 vccd1 vccd1 _12712_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_143_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18153_ _18153_/A _18153_/B _18153_/C vssd1 vssd1 vccd1 vccd1 _18156_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_81_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_104_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _24990_/CLK sky130_fd_sc_hd__clkbuf_16
X_15365_ _26019_/Q _25955_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15366_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12577_ _12577_/A vssd1 vssd1 vccd1 vccd1 _24968_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17104_ _25629_/Q vssd1 vssd1 vccd1 vccd1 _20322_/B sky130_fd_sc_hd__inv_2
X_14316_ _14316_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14316_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18084_ _18084_/A _20660_/B _18084_/C vssd1 vssd1 vccd1 vccd1 _20630_/B sky130_fd_sc_hd__nand3_1
X_15296_ _15296_/A vssd1 vssd1 vccd1 vccd1 _15305_/B sky130_fd_sc_hd__inv_2
XFILLER_0_180_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold308 hold308/A vssd1 vssd1 vccd1 vccd1 hold308/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold319 hold319/A vssd1 vssd1 vccd1 vccd1 hold319/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17035_ _19115_/B _25840_/Q _25776_/Q vssd1 vssd1 vccd1 vccd1 _17036_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_123_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14247_ _14242_/Y _14246_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold846/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14178_ _18674_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14178_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13129_ _13109_/X _13127_/X _13096_/X _13128_/X vssd1 vssd1 vccd1 vccd1 _13129_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _18986_/A _19729_/A vssd1 vssd1 vccd1 vccd1 _18986_/Y sky130_fd_sc_hd__nand2_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1008 _13246_/X vssd1 vssd1 vccd1 vccd1 _25093_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17937_ _20507_/B _19216_/A vssd1 vssd1 vccd1 vccd1 _17938_/B sky130_fd_sc_hd__nand2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1019 _25033_/Q vssd1 vssd1 vccd1 vccd1 _17414_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17868_ _17866_/Y _17867_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _25647_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19607_ _19607_/A _19607_/B vssd1 vssd1 vccd1 vccd1 _19607_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16819_ _16819_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16819_/Y sky130_fd_sc_hd__nand2_1
X_17799_ _18100_/A vssd1 vssd1 vccd1 vccd1 _18529_/A sky130_fd_sc_hd__buf_12
XFILLER_0_49_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19538_ _19536_/X _19537_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19538_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19469_ _26238_/Q _12537_/B hold494/X vssd1 vssd1 vccd1 vccd1 _19469_/Y sky130_fd_sc_hd__a21oi_1
X_21500_ _21500_/A _21500_/B _21500_/C vssd1 vssd1 vccd1 vccd1 _21501_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_119_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22480_ _22479_/A _22454_/X _22479_/B vssd1 vssd1 vccd1 vccd1 _22481_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21431_ _21481_/A _21434_/A vssd1 vssd1 vccd1 vccd1 _21432_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24150_ _24150_/A vssd1 vssd1 vccd1 vccd1 _26116_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21362_ _21362_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21362_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_185_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23101_ _23197_/A _23101_/B vssd1 vssd1 vccd1 vccd1 _23101_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20313_ _25846_/Q vssd1 vssd1 vccd1 vccd1 _20314_/B sky130_fd_sc_hd__inv_2
XFILLER_0_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24081_ _24081_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24082_/A sky130_fd_sc_hd__and2_1
XFILLER_0_47_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold820 hold820/A vssd1 vssd1 vccd1 vccd1 hold820/X sky130_fd_sc_hd__dlygate4sd3_1
X_21293_ _21293_/A _25876_/Q vssd1 vssd1 vccd1 vccd1 _21297_/B sky130_fd_sc_hd__nand2_1
Xhold831 hold831/A vssd1 vssd1 vccd1 vccd1 hold831/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23032_ _23031_/A _22849_/X _23031_/B vssd1 vssd1 vccd1 vccd1 _23033_/C sky130_fd_sc_hd__o21ai_1
Xhold842 hold842/A vssd1 vssd1 vccd1 vccd1 hold842/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 hold853/A vssd1 vssd1 vccd1 vccd1 hold853/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_20244_ _20244_/A _20244_/B _20244_/C vssd1 vssd1 vccd1 vccd1 _20245_/B sky130_fd_sc_hd__nand3_1
Xhold864 hold864/A vssd1 vssd1 vccd1 vccd1 hold864/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 hold875/A vssd1 vssd1 vccd1 vccd1 hold875/X sky130_fd_sc_hd__buf_1
Xhold886 hold886/A vssd1 vssd1 vccd1 vccd1 hold886/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold897 hold897/A vssd1 vssd1 vccd1 vccd1 hold897/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20175_ _20175_/A _20175_/B vssd1 vssd1 vccd1 vccd1 _20177_/A sky130_fd_sc_hd__nand2_1
Xhold2210 _24314_/X vssd1 vssd1 vccd1 vccd1 _24315_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2221 _26154_/Q vssd1 vssd1 vccd1 vccd1 hold2221/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2232 _14987_/Y vssd1 vssd1 vccd1 vccd1 _25422_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2243 _25963_/Q vssd1 vssd1 vccd1 vccd1 hold2243/X sky130_fd_sc_hd__dlygate4sd3_1
X_24983_ _24983_/CLK _24983_/D vssd1 vssd1 vccd1 vccd1 _24983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2254 _24017_/X vssd1 vssd1 vccd1 vccd1 _24018_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1520 _19825_/Y vssd1 vssd1 vccd1 vccd1 _25759_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2265 _26184_/Q vssd1 vssd1 vccd1 vccd1 hold2265/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1531 _25894_/Q vssd1 vssd1 vccd1 vccd1 _23085_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2276 _26201_/Q vssd1 vssd1 vccd1 vccd1 hold2276/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23934_ _23934_/A vssd1 vssd1 vccd1 vccd1 _26046_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2287 _24038_/X vssd1 vssd1 vccd1 vccd1 _24039_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1542 _21348_/Y vssd1 vssd1 vccd1 vccd1 _25814_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1553 _25819_/Q vssd1 vssd1 vccd1 vccd1 _21428_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2298 _15004_/Y vssd1 vssd1 vccd1 vccd1 _25424_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1564 _25776_/Q vssd1 vssd1 vccd1 vccd1 _20129_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1575 _20466_/Y vssd1 vssd1 vccd1 vccd1 _25785_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1586 _25821_/Q vssd1 vssd1 vccd1 vccd1 _21460_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23865_ hold2193/X hold2043/X _23907_/S vssd1 vssd1 vccd1 vccd1 _23866_/A sky130_fd_sc_hd__mux2_1
Xhold1597 _19583_/Y vssd1 vssd1 vccd1 vccd1 _25742_/D sky130_fd_sc_hd__dlygate4sd3_1
X_25604_ _25604_/CLK _25604_/D vssd1 vssd1 vccd1 vccd1 _25604_/Q sky130_fd_sc_hd__dfxtp_2
X_22816_ _22815_/A _22454_/X _22815_/B vssd1 vssd1 vccd1 vccd1 _22817_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23796_ _23796_/A vssd1 vssd1 vccd1 vccd1 _26003_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25535_ _25535_/CLK hold921/X vssd1 vssd1 vccd1 vccd1 hold920/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22747_ _23188_/A _22747_/B vssd1 vssd1 vccd1 vccd1 _22747_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xascon_wrapper_11 vssd1 vssd1 vccd1 vccd1 ascon_wrapper_11/HI io_oeb[8] sky130_fd_sc_hd__conb_1
X_12500_ _21203_/A vssd1 vssd1 vccd1 vccd1 _19483_/A sky130_fd_sc_hd__buf_12
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25466_ _26064_/CLK _25466_/D vssd1 vssd1 vccd1 vccd1 _25466_/Q sky130_fd_sc_hd__dfxtp_1
X_13480_ _13522_/A hold715/X vssd1 vssd1 vccd1 vccd1 hold716/A sky130_fd_sc_hd__nand2_1
X_22678_ _22680_/A vssd1 vssd1 vccd1 vccd1 _23188_/A sky130_fd_sc_hd__buf_8
XFILLER_0_48_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24417_ _24417_/A vssd1 vssd1 vccd1 vccd1 _26203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21629_ _21677_/B _21629_/B vssd1 vssd1 vccd1 vccd1 _21630_/C sky130_fd_sc_hd__nand2_1
X_25397_ _25999_/CLK _25397_/D vssd1 vssd1 vccd1 vccd1 _25397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15150_ _15148_/X _15149_/Y _15090_/X vssd1 vssd1 vccd1 vccd1 _25437_/D sky130_fd_sc_hd__a21oi_1
X_24348_ _24348_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24349_/A sky130_fd_sc_hd__and2_1
XFILLER_0_90_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14101_ _25811_/Q vssd1 vssd1 vccd1 vccd1 _18430_/B sky130_fd_sc_hd__inv_2
XFILLER_0_106_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15081_ _15079_/X hold2116/X _14928_/X vssd1 vssd1 vccd1 vccd1 _15081_/Y sky130_fd_sc_hd__a21oi_1
X_24279_ hold2598/X hold2309/X _24279_/S vssd1 vssd1 vccd1 vccd1 _24280_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_132_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26018_ _26021_/CLK _26018_/D vssd1 vssd1 vccd1 vccd1 _26018_/Q sky130_fd_sc_hd__dfxtp_1
X_14032_ _14118_/A hold710/X vssd1 vssd1 vccd1 vccd1 hold711/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18840_ _18838_/X _18269_/X _18839_/X vssd1 vssd1 vccd1 vccd1 _18841_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_140_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18771_ _18771_/A _25828_/Q _18771_/C vssd1 vssd1 vccd1 vccd1 _20605_/B sky130_fd_sc_hd__nand3_2
X_15983_ _22090_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _15985_/A sky130_fd_sc_hd__nand2_1
X_17722_ _17722_/A _17829_/A vssd1 vssd1 vccd1 vccd1 _17723_/B sky130_fd_sc_hd__nand2_1
X_14934_ _14947_/A _14948_/A vssd1 vssd1 vccd1 vccd1 _14934_/X sky130_fd_sc_hd__or2_1
XFILLER_0_175_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17653_ _18535_/A _17653_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _17653_/X sky130_fd_sc_hd__and3_1
X_14865_ _14858_/Y _14864_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14865_/Y sky130_fd_sc_hd__a21oi_1
X_16604_ hold871/X vssd1 vssd1 vccd1 vccd1 _16608_/B sky130_fd_sc_hd__inv_2
XFILLER_0_98_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13816_ _26268_/Q _13801_/X _13793_/X _13815_/Y vssd1 vssd1 vccd1 vccd1 _13817_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_188_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17584_ _17582_/Y _17583_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _17584_/Y sky130_fd_sc_hd__a21oi_1
X_14796_ _14794_/Y _14795_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14796_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19323_ _19321_/X _19322_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19323_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16535_ _16533_/Y _16535_/B vssd1 vssd1 vccd1 vccd1 _16541_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_161_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13747_ hold585/X _13746_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold586/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19254_ _19254_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _19254_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16466_ _16466_/A _16466_/B vssd1 vssd1 vccd1 vccd1 _16467_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_156_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13678_ _13703_/A _13678_/B vssd1 vssd1 vccd1 vccd1 _13678_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_85_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18205_ _18205_/A _20964_/A vssd1 vssd1 vccd1 vccd1 _18555_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_171_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15417_ _16834_/B vssd1 vssd1 vccd1 vccd1 _22832_/B sky130_fd_sc_hd__inv_2
XFILLER_0_155_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12629_ _12629_/A _12629_/B vssd1 vssd1 vccd1 vccd1 _12635_/A sky130_fd_sc_hd__nand2_1
X_19185_ _19175_/X _19184_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19185_/Y sky130_fd_sc_hd__o21ai_1
X_16397_ _16473_/A hold518/X vssd1 vssd1 vccd1 vccd1 hold519/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18136_ _18136_/A _25798_/Q _18136_/C vssd1 vssd1 vccd1 vccd1 _20915_/B sky130_fd_sc_hd__nand3_2
X_15348_ _16806_/B vssd1 vssd1 vccd1 vccd1 _22766_/B sky130_fd_sc_hd__inv_2
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold105 hold105/A vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__dlygate4sd3_1
X_18067_ _18067_/A _18067_/B _20251_/B vssd1 vssd1 vccd1 vccd1 _18076_/A sky130_fd_sc_hd__and3_2
X_15279_ _15827_/A _15307_/B vssd1 vssd1 vccd1 vccd1 _15279_/Y sky130_fd_sc_hd__nand2_1
Xhold116 hold116/A vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 hold127/A vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 hold138/A vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ _25583_/Q vssd1 vssd1 vccd1 vccd1 _20067_/B sky130_fd_sc_hd__inv_2
Xhold149 hold149/A vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18969_ _18967_/X _18879_/X _18968_/X vssd1 vssd1 vccd1 vccd1 _18971_/A sky130_fd_sc_hd__a21o_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21980_ _21980_/A _25873_/Q vssd1 vssd1 vccd1 vccd1 _21980_/Y sky130_fd_sc_hd__nand2_1
X_20931_ _20931_/A _20931_/B vssd1 vssd1 vccd1 vccd1 _20932_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23650_ hold2068/X _25956_/Q _23677_/S vssd1 vssd1 vccd1 vccd1 _23650_/X sky130_fd_sc_hd__mux2_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20862_ _20862_/A _20862_/B vssd1 vssd1 vccd1 vccd1 _20864_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22601_ _22601_/A _22601_/B vssd1 vssd1 vccd1 vccd1 _22602_/A sky130_fd_sc_hd__xor2_1
X_23581_ _23581_/A _23581_/B vssd1 vssd1 vccd1 vccd1 _23581_/Y sky130_fd_sc_hd__nand2_1
X_20793_ _20793_/A _25897_/Q vssd1 vssd1 vccd1 vccd1 _20798_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25320_ _26252_/CLK hold70/X vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22532_ _16736_/B _22421_/X _22526_/X _22527_/Y _22531_/X vssd1 vssd1 vccd1 vccd1
+ _22533_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25251_ _25864_/CLK hold568/X vssd1 vssd1 vccd1 vccd1 hold566/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22463_ _25827_/Q _22463_/B vssd1 vssd1 vccd1 vccd1 _22463_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_151_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24202_ _24202_/A vssd1 vssd1 vccd1 vccd1 _26133_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21414_ _21417_/A _21466_/A vssd1 vssd1 vccd1 vccd1 _21416_/A sky130_fd_sc_hd__nand2_1
X_22394_ _19744_/A _22393_/A _22393_/Y vssd1 vssd1 vccd1 vccd1 _22396_/A sky130_fd_sc_hd__o21ai_1
X_25182_ _26275_/CLK hold735/X vssd1 vssd1 vccd1 vccd1 hold733/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24133_ hold2252/X hold2135/X _24203_/S vssd1 vssd1 vccd1 vccd1 _24134_/A sky130_fd_sc_hd__mux2_1
X_21345_ _21345_/A _21345_/B vssd1 vssd1 vccd1 vccd1 _21346_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_142_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24064_ _24064_/A vssd1 vssd1 vccd1 vccd1 _26088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21276_ _21276_/A _21276_/B _21276_/C vssd1 vssd1 vccd1 vccd1 _21280_/A sky130_fd_sc_hd__nand3_1
Xhold650 hold650/A vssd1 vssd1 vccd1 vccd1 hold650/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 hold661/A vssd1 vssd1 vccd1 vccd1 hold661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 hold672/A vssd1 vssd1 vccd1 vccd1 hold672/X sky130_fd_sc_hd__dlygate4sd3_1
X_23015_ _23015_/A _23015_/B _23191_/C vssd1 vssd1 vccd1 vccd1 _23017_/A sky130_fd_sc_hd__or3_1
Xhold683 hold683/A vssd1 vssd1 vccd1 vccd1 hold683/X sky130_fd_sc_hd__dlygate4sd3_1
X_20227_ _26282_/Q _20078_/X hold611/X vssd1 vssd1 vccd1 vccd1 _20230_/B sky130_fd_sc_hd__a21oi_1
Xhold694 hold694/A vssd1 vssd1 vccd1 vccd1 hold694/X sky130_fd_sc_hd__dlygate4sd3_1
X_20158_ _20158_/A _20158_/B vssd1 vssd1 vccd1 vccd1 _20159_/A sky130_fd_sc_hd__nand2_1
Xhold2040 _25449_/Q vssd1 vssd1 vccd1 vccd1 _15347_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2051 _26018_/Q vssd1 vssd1 vccd1 vccd1 hold2051/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2062 _23895_/X vssd1 vssd1 vccd1 vccd1 _23896_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24966_ _25418_/CLK _24966_/D vssd1 vssd1 vccd1 vccd1 _24966_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2073 _23699_/X vssd1 vssd1 vccd1 vccd1 _23700_/A sky130_fd_sc_hd__dlygate4sd3_1
X_12980_ _17514_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _12980_/X sky130_fd_sc_hd__or2_1
X_20089_ _20092_/A _20092_/C vssd1 vssd1 vccd1 vccd1 _20091_/A sky130_fd_sc_hd__nand2_1
Xhold2084 _23311_/X vssd1 vssd1 vccd1 vccd1 _23312_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2095 _23638_/X vssd1 vssd1 vccd1 vccd1 _23639_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1350 _19866_/Y vssd1 vssd1 vccd1 vccd1 _25762_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1361 _25396_/Q vssd1 vssd1 vccd1 vccd1 _14768_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23917_ hold1978/X _26043_/Q _23920_/S vssd1 vssd1 vccd1 vccd1 _23917_/X sky130_fd_sc_hd__mux2_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1372 _13282_/X vssd1 vssd1 vccd1 vccd1 _25099_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24897_ _15799_/A _15816_/B _24945_/S vssd1 vssd1 vccd1 vccd1 _24897_/X sky130_fd_sc_hd__mux2_1
Xhold1383 _15784_/Y vssd1 vssd1 vccd1 vccd1 hold1383/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1394 _19932_/Y vssd1 vssd1 vccd1 vccd1 _25767_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _14648_/Y hold288/X _14646_/X vssd1 vssd1 vccd1 vccd1 hold289/A sky130_fd_sc_hd__a21oi_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23848_ _23848_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23849_/A sky130_fd_sc_hd__and2_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _26234_/Q _13426_/X _13468_/X _13600_/Y vssd1 vssd1 vccd1 vccd1 _13602_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14581_ _14581_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14581_/Y sky130_fd_sc_hd__nand2_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23779_ _14843_/B _14851_/B _23831_/S vssd1 vssd1 vccd1 vccd1 _23780_/A sky130_fd_sc_hd__mux2_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16320_ hold873/X _16320_/B vssd1 vssd1 vccd1 vccd1 _16321_/B sky130_fd_sc_hd__or2_1
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25518_ _25539_/CLK hold895/X vssd1 vssd1 vccd1 vccd1 hold894/A sky130_fd_sc_hd__dfxtp_1
X_13532_ _17800_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13532_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_32_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16251_ _16264_/B _16251_/B vssd1 vssd1 vccd1 vccd1 _16269_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_152_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25449_ _25450_/CLK _25449_/D vssd1 vssd1 vccd1 vccd1 _25449_/Q sky130_fd_sc_hd__dfxtp_1
X_13463_ _13522_/A hold452/X vssd1 vssd1 vccd1 vccd1 hold453/A sky130_fd_sc_hd__nand2_1
X_15202_ _15956_/A hold927/X vssd1 vssd1 vccd1 vccd1 _15202_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_164_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16182_ _16182_/A _16182_/B vssd1 vssd1 vccd1 vccd1 _16184_/A sky130_fd_sc_hd__nand2_1
X_13394_ _13315_/X _13392_/X _13300_/X _13393_/X vssd1 vssd1 vccd1 vccd1 _13394_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15133_ _15133_/A vssd1 vssd1 vccd1 vccd1 _15144_/B sky130_fd_sc_hd__inv_2
XFILLER_0_23_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15064_ _15065_/B _15065_/A vssd1 vssd1 vccd1 vccd1 _15066_/A sky130_fd_sc_hd__or2_1
XFILLER_0_65_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19941_ _19936_/X _19940_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19941_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14015_ _25797_/Q vssd1 vssd1 vccd1 vccd1 _18102_/B sky130_fd_sc_hd__inv_2
X_19872_ _20790_/A _18867_/A _20795_/C vssd1 vssd1 vccd1 vccd1 _19948_/A sky130_fd_sc_hd__o21a_2
X_18823_ _18821_/Y _18822_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25685_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15966_ _16212_/A hold929/X vssd1 vssd1 vccd1 vccd1 _15966_/Y sky130_fd_sc_hd__nand2_1
X_18754_ _18754_/A _18754_/B _18754_/C vssd1 vssd1 vccd1 vccd1 _22465_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14917_ _14917_/A _14917_/B vssd1 vssd1 vccd1 vccd1 _14919_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17705_ _17705_/A _17705_/B _17705_/C vssd1 vssd1 vccd1 vccd1 _17738_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_175_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15897_ _15870_/Y _15895_/A _15896_/Y vssd1 vssd1 vccd1 vccd1 _15897_/X sky130_fd_sc_hd__a21o_1
X_18685_ _22391_/B _25632_/Q vssd1 vssd1 vccd1 vccd1 _18687_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14848_ _14864_/A _14848_/B vssd1 vssd1 vccd1 vccd1 _14848_/Y sky130_fd_sc_hd__nand2_1
X_17636_ _17634_/Y _17635_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _25642_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_188_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17567_ _17605_/A _17567_/B vssd1 vssd1 vccd1 vccd1 _17567_/Y sky130_fd_sc_hd__nand2_1
X_14779_ _15839_/A _25990_/Q vssd1 vssd1 vccd1 vccd1 _22036_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16518_ _16516_/X _16517_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 hold941/A sky130_fd_sc_hd__a21oi_1
X_19306_ _19322_/B _19393_/B vssd1 vssd1 vccd1 vccd1 _19308_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17498_ _17498_/A _17548_/A vssd1 vssd1 vccd1 vccd1 _17499_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16449_ _16447_/Y _16448_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 hold867/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19237_ _19235_/Y _21228_/A _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _19239_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19168_ _19166_/X _19167_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19168_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18119_ _18119_/A _18119_/B vssd1 vssd1 vccd1 vccd1 _18122_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19099_ _20247_/A _19097_/Y _20251_/C vssd1 vssd1 vccd1 vccd1 _19211_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_170_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21130_ _21132_/B _21132_/C vssd1 vssd1 vccd1 vccd1 _21131_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_112_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21061_ _21564_/B _21513_/C vssd1 vssd1 vccd1 vccd1 _21062_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20012_ _20014_/B _20014_/C vssd1 vssd1 vccd1 vccd1 _20013_/A sky130_fd_sc_hd__nand2_1
X_24820_ hold2561/X _26335_/Q _24835_/S vssd1 vssd1 vccd1 vccd1 _24820_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24751_ hold2742/X _26312_/Q _24817_/S vssd1 vssd1 vccd1 vccd1 _24751_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21963_ _21961_/X _21962_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _21963_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_146_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk clkbuf_leaf_95_clk/A vssd1 vssd1 vccd1 vccd1 _25913_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23702_ _25972_/Q hold2128/X _23754_/S vssd1 vssd1 vccd1 vccd1 _23702_/X sky130_fd_sc_hd__mux2_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20914_ _20916_/B _20916_/C vssd1 vssd1 vccd1 vccd1 _20915_/A sky130_fd_sc_hd__nand2_1
X_24682_ _24682_/A vssd1 vssd1 vccd1 vccd1 _26289_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21894_ _21892_/X _21893_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _21894_/Y sky130_fd_sc_hd__a21oi_2
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23633_ _23633_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23634_/A sky130_fd_sc_hd__and2_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20845_ _20845_/A _20845_/B vssd1 vssd1 vccd1 vccd1 _20846_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_178_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23564_ _24922_/S hold392/A _23563_/X vssd1 vssd1 vccd1 vccd1 _23564_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20776_ _20776_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _20776_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_153_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25303_ _26136_/CLK hold301/X vssd1 vssd1 vccd1 vccd1 hold299/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22515_ _22515_/A _22515_/B vssd1 vssd1 vccd1 vccd1 _22515_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_119_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26283_ _26283_/CLK _26283_/D vssd1 vssd1 vccd1 vccd1 _26283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23495_ _23491_/Y _23494_/Y _24858_/S vssd1 vssd1 vccd1 vccd1 _23495_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_135_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25234_ _25817_/CLK hold822/X vssd1 vssd1 vccd1 vccd1 hold821/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22446_ _22446_/A _22446_/B vssd1 vssd1 vccd1 vccd1 _22447_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25165_ _25748_/CLK hold403/X vssd1 vssd1 vccd1 vccd1 hold401/A sky130_fd_sc_hd__dfxtp_1
X_22377_ _22958_/B vssd1 vssd1 vccd1 vccd1 _22957_/B sky130_fd_sc_hd__inv_2
XFILLER_0_33_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24116_ _24116_/A vssd1 vssd1 vccd1 vccd1 _26105_/D sky130_fd_sc_hd__clkbuf_1
X_21328_ _21636_/A _21328_/B _21327_/X vssd1 vssd1 vccd1 vccd1 _21329_/B sky130_fd_sc_hd__or3b_2
X_25096_ _26308_/CLK _25096_/D vssd1 vssd1 vccd1 vccd1 _25096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24047_ _26083_/Q hold2326/X _24047_/S vssd1 vssd1 vccd1 vccd1 _24047_/X sky130_fd_sc_hd__mux2_1
X_21259_ _21259_/A _21259_/B vssd1 vssd1 vccd1 vccd1 _21260_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold480 hold480/A vssd1 vssd1 vccd1 vccd1 hold480/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 hold491/A vssd1 vssd1 vccd1 vccd1 hold491/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15820_ _15820_/A _15830_/A vssd1 vssd1 vccd1 vccd1 _15820_/Y sky130_fd_sc_hd__nand2_1
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25998_ _25998_/CLK _25998_/D vssd1 vssd1 vccd1 vccd1 _25998_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _15749_/X _15750_/Y _15464_/X vssd1 vssd1 vccd1 vccd1 _25471_/D sky130_fd_sc_hd__a21oi_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24949_ _24939_/X _24948_/X _24949_/S vssd1 vssd1 vccd1 vccd1 _24950_/A sky130_fd_sc_hd__mux2_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12963_ _26126_/Q _12907_/X _12962_/X vssd1 vssd1 vccd1 vccd1 _12963_/X sky130_fd_sc_hd__a21o_1
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1180 _16828_/Y vssd1 vssd1 vccd1 vccd1 _25557_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_84_clk clkbuf_leaf_95_clk/A vssd1 vssd1 vccd1 vccd1 _26046_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _14899_/B vssd1 vssd1 vccd1 vccd1 _14900_/A sky130_fd_sc_hd__inv_6
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1191 _25730_/Q vssd1 vssd1 vccd1 vccd1 _19410_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18470_ _18470_/A _18470_/B _18470_/C vssd1 vssd1 vccd1 vccd1 _22097_/A sky130_fd_sc_hd__nand3_2
X_15682_ _26037_/Q _25973_/Q _15773_/S vssd1 vssd1 vccd1 vccd1 _15683_/A sky130_fd_sc_hd__mux2_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _26113_/Q _12748_/X _12893_/X vssd1 vssd1 vccd1 vccd1 _12894_/X sky130_fd_sc_hd__a21o_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17421_ _19588_/A _17421_/B vssd1 vssd1 vccd1 vccd1 _17644_/B sky130_fd_sc_hd__xor2_4
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _14645_/A hold143/X vssd1 vssd1 vccd1 vccd1 hold144/A sky130_fd_sc_hd__nand2_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17352_ _17623_/A _17352_/B vssd1 vssd1 vccd1 vccd1 _17352_/X sky130_fd_sc_hd__xor2_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _14585_/A hold161/X vssd1 vssd1 vccd1 vccd1 hold162/A sky130_fd_sc_hd__nand2_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ hold958/X vssd1 vssd1 vccd1 vccd1 _16306_/B sky130_fd_sc_hd__inv_2
XFILLER_0_27_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13515_ hold769/X _13514_/Y _12558_/B vssd1 vssd1 vccd1 vccd1 hold770/A sky130_fd_sc_hd__a21oi_1
X_17283_ _17281_/X _17241_/X _17282_/X vssd1 vssd1 vccd1 vccd1 _17284_/A sky130_fd_sc_hd__a21o_1
X_14495_ _14525_/A hold110/X vssd1 vssd1 vccd1 vccd1 hold111/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19022_ _19186_/A _19802_/A vssd1 vssd1 vccd1 vccd1 _19022_/Y sky130_fd_sc_hd__nand2_1
X_16234_ _16235_/A _16401_/C hold972/X vssd1 vssd1 vccd1 vccd1 _16236_/A sky130_fd_sc_hd__a21oi_1
X_13446_ _19061_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13446_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16165_ _16676_/A _16165_/B vssd1 vssd1 vccd1 vccd1 _16168_/A sky130_fd_sc_hd__or2_1
X_13377_ _13377_/A vssd1 vssd1 vccd1 vccd1 _19729_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15116_ _22453_/B _15116_/B vssd1 vssd1 vccd1 vccd1 _22449_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_51_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16096_ _16096_/A _16096_/B vssd1 vssd1 vccd1 vccd1 _16103_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_121_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15047_ _15045_/X hold2289/X _14928_/X vssd1 vssd1 vccd1 vccd1 _15047_/Y sky130_fd_sc_hd__a21oi_1
X_19924_ _20087_/A _22718_/B _25645_/Q vssd1 vssd1 vccd1 vccd1 _20092_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_177_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19855_ _19854_/Y _19130_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19857_/A
+ sky130_fd_sc_hd__a211o_1
X_18806_ _20673_/B _19830_/A vssd1 vssd1 vccd1 vccd1 _18807_/B sky130_fd_sc_hd__nand2_1
X_19786_ _19785_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19787_/B
+ sky130_fd_sc_hd__a211o_1
X_16998_ _18529_/C vssd1 vssd1 vccd1 vccd1 _21716_/A sky130_fd_sc_hd__buf_8
X_18737_ _18940_/A _19003_/A vssd1 vssd1 vccd1 vccd1 _18738_/B sky130_fd_sc_hd__xnor2_1
X_15949_ _22001_/B _16691_/B vssd1 vssd1 vccd1 vccd1 _15951_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_183_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18668_ _25887_/Q _22369_/A vssd1 vssd1 vccd1 vccd1 _18676_/A sky130_fd_sc_hd__or2_2
XFILLER_0_148_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17619_ _17619_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _17619_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18599_ _21791_/A vssd1 vssd1 vccd1 vccd1 _18963_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20630_ _20630_/A _20630_/B vssd1 vssd1 vccd1 vccd1 _20632_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20561_ _23037_/B vssd1 vssd1 vccd1 vccd1 _22468_/B sky130_fd_sc_hd__inv_2
XFILLER_0_50_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22300_ _19687_/A _22299_/A _22299_/Y vssd1 vssd1 vccd1 vccd1 _22302_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23280_ _23280_/A vssd1 vssd1 vccd1 vccd1 _25918_/D sky130_fd_sc_hd__clkbuf_1
X_20492_ _20492_/A _20492_/B _21195_/C vssd1 vssd1 vccd1 vccd1 _20496_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_144_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22231_ _22229_/Y _22230_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _22231_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22162_ _22162_/A _22162_/B vssd1 vssd1 vccd1 vccd1 _22162_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_41_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21113_ _21597_/B _21548_/B vssd1 vssd1 vccd1 vccd1 _21114_/B sky130_fd_sc_hd__nand2_1
X_22093_ _22093_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _22093_/X sky130_fd_sc_hd__and2_1
XFILLER_0_160_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25921_ _25925_/CLK hold857/X vssd1 vssd1 vccd1 vccd1 hold855/A sky130_fd_sc_hd__dfxtp_1
X_21044_ _21044_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _21044_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_157_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25852_ _26207_/CLK _25852_/D vssd1 vssd1 vccd1 vccd1 _25852_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24803_ _24803_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24804_/A sky130_fd_sc_hd__and2_1
X_25783_ _25783_/CLK _25783_/D vssd1 vssd1 vccd1 vccd1 _25783_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_158_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22995_ _22995_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22995_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_66_clk _25472_/CLK vssd1 vssd1 vccd1 vccd1 _26060_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24734_ hold2476/X _26307_/Q _24740_/S vssd1 vssd1 vccd1 vccd1 _24734_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_96_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21946_ _21946_/A _25872_/Q vssd1 vssd1 vccd1 vccd1 _21946_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_119_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24665_ _24665_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24666_/A sky130_fd_sc_hd__and2_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21877_ _21877_/A _25870_/Q vssd1 vssd1 vccd1 vccd1 _21877_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23616_ hold2140/X _25945_/Q _23677_/S vssd1 vssd1 vccd1 vccd1 _23616_/X sky130_fd_sc_hd__mux2_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20828_ _20828_/A _22640_/B vssd1 vssd1 vccd1 vccd1 _20829_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24596_ _24596_/A vssd1 vssd1 vccd1 vccd1 _26261_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26335_ _26335_/CLK _26335_/D vssd1 vssd1 vccd1 vccd1 _26335_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23547_ _24942_/S hold470/A _23546_/X vssd1 vssd1 vccd1 vccd1 _23547_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_181_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20759_ _20758_/B _20759_/B _20759_/C vssd1 vssd1 vccd1 vccd1 _20760_/B sky130_fd_sc_hd__nand3b_1
X_13300_ _24560_/A vssd1 vssd1 vccd1 vccd1 _13300_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14280_ _14345_/A vssd1 vssd1 vccd1 vccd1 _14280_/X sky130_fd_sc_hd__buf_8
XFILLER_0_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26266_ _26267_/CLK _26266_/D vssd1 vssd1 vccd1 vccd1 _26266_/Q sky130_fd_sc_hd__dfxtp_2
X_23478_ _24956_/S hold197/A _23477_/X vssd1 vssd1 vccd1 vccd1 _23478_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_134_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25217_ _26303_/CLK hold505/X vssd1 vssd1 vccd1 vccd1 hold503/A sky130_fd_sc_hd__dfxtp_1
X_13231_ _18535_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13231_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22429_ _22429_/A _22900_/B vssd1 vssd1 vccd1 vccd1 _22429_/Y sky130_fd_sc_hd__nand2_1
X_26197_ _26198_/CLK _26197_/D vssd1 vssd1 vccd1 vccd1 _26197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25148_ _25727_/CLK hold466/X vssd1 vssd1 vccd1 vccd1 hold464/A sky130_fd_sc_hd__dfxtp_1
X_13162_ _18313_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13162_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25079_ _26164_/CLK _25079_/D vssd1 vssd1 vccd1 vccd1 _25079_/Q sky130_fd_sc_hd__dfxtp_1
X_13093_ _26279_/Q _25648_/Q vssd1 vssd1 vccd1 vccd1 _14497_/A sky130_fd_sc_hd__xor2_1
X_17970_ _21889_/A _25586_/Q vssd1 vssd1 vccd1 vccd1 _17971_/C sky130_fd_sc_hd__nand2_1
X_16921_ _16935_/A _16926_/B vssd1 vssd1 vccd1 vccd1 _16923_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19640_ _26250_/Q _19483_/X hold572/X vssd1 vssd1 vccd1 vccd1 _19640_/Y sky130_fd_sc_hd__a21oi_1
X_16852_ _16850_/Y _16851_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16852_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15803_ _15956_/A hold902/X vssd1 vssd1 vccd1 vccd1 _15803_/Y sky130_fd_sc_hd__nand2_1
X_16783_ _16781_/Y _15305_/A _16782_/Y vssd1 vssd1 vccd1 vccd1 _16783_/Y sky130_fd_sc_hd__o21ai_1
X_19571_ _26245_/Q hold791/X vssd1 vssd1 vccd1 vccd1 _19571_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13995_ _25794_/Q vssd1 vssd1 vccd1 vccd1 _17958_/B sky130_fd_sc_hd__inv_2
XFILLER_0_73_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15734_ _15956_/A hold883/X vssd1 vssd1 vccd1 vccd1 _15734_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18522_ _20132_/B _19630_/A vssd1 vssd1 vccd1 vccd1 _18523_/B sky130_fd_sc_hd__nand2_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ _26251_/Q _25620_/Q vssd1 vssd1 vccd1 vccd1 _14409_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15665_ _16926_/B vssd1 vssd1 vccd1 vccd1 _23063_/B sky130_fd_sc_hd__inv_2
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18453_ _18657_/A _18798_/A vssd1 vssd1 vccd1 vccd1 _18454_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12877_ _12726_/B _14367_/A _12752_/X _25607_/Q vssd1 vssd1 vccd1 vccd1 _12877_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ _17624_/A _17404_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17404_/X sky130_fd_sc_hd__and3_1
X_14616_ _14614_/Y hold75/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__a21oi_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18384_ _18446_/A _19624_/B _21716_/A vssd1 vssd1 vccd1 vccd1 _18385_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_96_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15596_ _26032_/Q _25968_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15597_/A sky130_fd_sc_hd__mux2_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _17335_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17335_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14547_ _14545_/Y hold129/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold130/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17266_ _25705_/Q _17266_/B vssd1 vssd1 vccd1 vccd1 _17622_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_114_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14478_ _14476_/Y hold69/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16217_ _16217_/A vssd1 vssd1 vccd1 vccd1 _16217_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_153_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19005_ _19026_/A _19005_/B _22786_/A vssd1 vssd1 vccd1 vccd1 _19005_/X sky130_fd_sc_hd__and3_1
X_13429_ _13220_/A _14669_/A _13242_/A _19844_/A vssd1 vssd1 vccd1 vccd1 _13429_/X
+ sky130_fd_sc_hd__a22o_1
X_17197_ _19802_/A _17197_/B vssd1 vssd1 vccd1 vccd1 _17585_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_12_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16148_ _16148_/A hold861/X vssd1 vssd1 vccd1 vccd1 _16149_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_12_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16079_ _22292_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _16081_/A sky130_fd_sc_hd__nand2_1
X_19907_ _19906_/Y _19130_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19909_/A
+ sky130_fd_sc_hd__a211o_1
Xhold2606 _26217_/Q vssd1 vssd1 vccd1 vccd1 hold2606/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2617 _26223_/Q vssd1 vssd1 vccd1 vccd1 hold2617/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2628 _26281_/Q vssd1 vssd1 vccd1 vccd1 hold2628/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2639 _26251_/Q vssd1 vssd1 vccd1 vccd1 hold2639/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1905 _25984_/Q vssd1 vssd1 vccd1 vccd1 _14723_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1916 _23249_/Y vssd1 vssd1 vccd1 vccd1 hold1916/X sky130_fd_sc_hd__dlygate4sd3_1
X_19838_ _19975_/A _19838_/B vssd1 vssd1 vccd1 vccd1 _19838_/Y sky130_fd_sc_hd__nand2_1
Xhold1927 _23635_/X vssd1 vssd1 vccd1 vccd1 _23636_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1938 _26210_/Q vssd1 vssd1 vccd1 vccd1 hold1938/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1949 _26162_/Q vssd1 vssd1 vccd1 vccd1 hold1949/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput1 io_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_2
X_19769_ _19767_/Y _19768_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19769_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_48_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _26032_/CLK sky130_fd_sc_hd__clkbuf_16
X_21800_ _21800_/A _25859_/Q vssd1 vssd1 vccd1 vccd1 _21800_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_91_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22780_ _15367_/B _22680_/X _14273_/X vssd1 vssd1 vccd1 vccd1 _22780_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21731_ _21731_/A _21731_/B vssd1 vssd1 vccd1 vccd1 _21731_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_91_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24450_ _24450_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24451_/A sky130_fd_sc_hd__and2_1
X_21662_ _21662_/A _21662_/B _21662_/C vssd1 vssd1 vccd1 vccd1 _21663_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_47_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23401_ hold245/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23401_/X sky130_fd_sc_hd__or2b_1
X_20613_ _20613_/A _21276_/C _20613_/C vssd1 vssd1 vccd1 vccd1 _20614_/B sky130_fd_sc_hd__nand3_1
X_24381_ _24381_/A vssd1 vssd1 vccd1 vccd1 _26191_/D sky130_fd_sc_hd__clkbuf_1
X_21593_ _21595_/A _21645_/B vssd1 vssd1 vccd1 vccd1 _21594_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26120_ _26121_/CLK _26120_/D vssd1 vssd1 vccd1 vccd1 _26120_/Q sky130_fd_sc_hd__dfxtp_1
X_23332_ _23332_/A vssd1 vssd1 vccd1 vccd1 _25928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20544_ _20660_/A _20544_/B vssd1 vssd1 vccd1 vccd1 _20544_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26051_ _26051_/CLK _26051_/D vssd1 vssd1 vccd1 vccd1 _26051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23263_ hold875/X _23264_/A vssd1 vssd1 vccd1 vccd1 _23263_/X sky130_fd_sc_hd__or2_1
XFILLER_0_171_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20475_ _20474_/B _20475_/B _20475_/C vssd1 vssd1 vccd1 vccd1 _20476_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_104_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25002_ _26249_/CLK hold79/X vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dfxtp_1
X_22214_ _22214_/A _22214_/B vssd1 vssd1 vccd1 vccd1 _22858_/B sky130_fd_sc_hd__nand2_2
X_23194_ _15808_/A _22421_/A _23188_/X _23189_/Y _23193_/X vssd1 vssd1 vccd1 vccd1
+ _23194_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22145_ _22145_/A _22145_/B vssd1 vssd1 vccd1 vccd1 _22145_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_112_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22076_ _25784_/Q _22076_/B vssd1 vssd1 vccd1 vccd1 _22076_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_22_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25904_ _26269_/CLK _25904_/D vssd1 vssd1 vccd1 vccd1 _25904_/Q sky130_fd_sc_hd__dfxtp_2
X_21027_ _21027_/A _21027_/B vssd1 vssd1 vccd1 vccd1 _21029_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25835_ _25835_/CLK _25835_/D vssd1 vssd1 vccd1 vccd1 _25835_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_96_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_clk _25184_/CLK vssd1 vssd1 vccd1 vccd1 _26269_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12800_ _26095_/Q _12748_/X _12799_/X vssd1 vssd1 vccd1 vccd1 _12800_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_97_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25766_ _25770_/CLK _25766_/D vssd1 vssd1 vccd1 vccd1 _25766_/Q sky130_fd_sc_hd__dfxtp_1
X_13780_ _13880_/A hold847/X vssd1 vssd1 vccd1 vccd1 _13780_/Y sky130_fd_sc_hd__nand2_1
X_22978_ _22978_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22978_/Y sky130_fd_sc_hd__nand2_1
X_12731_ _15795_/A vssd1 vssd1 vccd1 vccd1 _15543_/B sky130_fd_sc_hd__clkinv_8
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24717_ _24717_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24718_/A sky130_fd_sc_hd__and2_1
X_21929_ _21927_/X _21928_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _21929_/Y sky130_fd_sc_hd__a21oi_2
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25697_ _26324_/CLK _25697_/D vssd1 vssd1 vccd1 vccd1 _25697_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ _25455_/Q vssd1 vssd1 vccd1 vccd1 _15458_/B sky130_fd_sc_hd__inv_2
XFILLER_0_167_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12662_ _12662_/A _24836_/B _12662_/C vssd1 vssd1 vccd1 vccd1 _12662_/X sky130_fd_sc_hd__and3_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24648_ hold2725/X hold1945/X _24664_/S vssd1 vssd1 vccd1 vccd1 _24649_/A sky130_fd_sc_hd__mux2_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14401_ _14404_/A hold200/X vssd1 vssd1 vccd1 vccd1 hold201/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15381_ _16820_/B vssd1 vssd1 vccd1 vccd1 _22799_/B sky130_fd_sc_hd__inv_2
XFILLER_0_26_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12593_ _12593_/A vssd1 vssd1 vccd1 vccd1 _24971_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24579_ _24579_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24580_/A sky130_fd_sc_hd__and2_1
X_17120_ _17463_/A _17541_/A vssd1 vssd1 vccd1 vccd1 _17121_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14332_ _14344_/A hold335/X vssd1 vssd1 vccd1 vccd1 hold336/A sky130_fd_sc_hd__nand2_1
X_26318_ _26325_/CLK _26318_/D vssd1 vssd1 vccd1 vccd1 _26318_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17051_ _19138_/B _25841_/Q _25777_/Q vssd1 vssd1 vccd1 vccd1 _17052_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_135_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14263_ _26340_/Q _13518_/B _14170_/X _14262_/Y vssd1 vssd1 vccd1 vccd1 _14264_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26249_ _26249_/CLK _26249_/D vssd1 vssd1 vccd1 vccd1 _26249_/Q sky130_fd_sc_hd__dfxtp_2
X_16002_ _15987_/B _15999_/B _15986_/A vssd1 vssd1 vccd1 vccd1 _16002_/Y sky130_fd_sc_hd__o21ai_1
X_13214_ _13214_/A vssd1 vssd1 vccd1 vccd1 _19359_/A sky130_fd_sc_hd__buf_4
X_14194_ _14236_/A hold827/X vssd1 vssd1 vccd1 vccd1 _14194_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13145_ _13109_/X _13143_/X _13096_/X _13144_/X vssd1 vssd1 vccd1 vccd1 hold991/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ _18611_/A _17957_/B vssd1 vssd1 vccd1 vccd1 _17955_/A sky130_fd_sc_hd__nand2_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13076_ _13018_/X _13074_/X _13005_/X _13075_/X vssd1 vssd1 vccd1 vccd1 _13076_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16904_ _16904_/A _16904_/B vssd1 vssd1 vccd1 vccd1 _16904_/Y sky130_fd_sc_hd__nand2_1
X_17884_ _17884_/A vssd1 vssd1 vccd1 vccd1 _19032_/A sky130_fd_sc_hd__clkinv_4
X_19623_ _19615_/X _19622_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19623_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16835_ _16833_/Y _16834_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16835_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19554_ _19723_/A _19554_/B vssd1 vssd1 vccd1 vccd1 _19554_/Y sky130_fd_sc_hd__nand2_1
X_16766_ _16980_/A _16771_/B vssd1 vssd1 vccd1 vccd1 _16768_/B sky130_fd_sc_hd__nand2_1
X_13978_ _14061_/A _13978_/B vssd1 vssd1 vccd1 vccd1 _13978_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18505_ _18792_/A _18509_/B vssd1 vssd1 vccd1 vccd1 _18507_/A sky130_fd_sc_hd__nand2_1
X_15717_ _15715_/X _15716_/Y _15464_/X vssd1 vssd1 vccd1 vccd1 _25469_/D sky130_fd_sc_hd__a21oi_1
X_12929_ _12840_/X _12927_/X _12917_/X _12928_/X vssd1 vssd1 vccd1 vccd1 _12929_/X
+ sky130_fd_sc_hd__o211a_1
X_16697_ _16697_/A _16697_/B vssd1 vssd1 vccd1 vccd1 _16697_/Y sky130_fd_sc_hd__nand2_1
X_19485_ _26239_/Q hold841/X vssd1 vssd1 vccd1 vccd1 _19485_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_180_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18436_ _18434_/X _18269_/X _18435_/X vssd1 vssd1 vccd1 vccd1 _18437_/A sky130_fd_sc_hd__a21o_1
X_15648_ _26035_/Q _25971_/Q _15773_/S vssd1 vssd1 vccd1 vccd1 _15649_/A sky130_fd_sc_hd__mux2_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15579_ _15560_/A _15611_/A _15578_/X vssd1 vssd1 vccd1 vccd1 _15579_/X sky130_fd_sc_hd__a21bo_1
X_18367_ _18952_/A _18367_/B _18952_/C vssd1 vssd1 vccd1 vccd1 _18368_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17318_ _20088_/B _25901_/Q _25837_/Q vssd1 vssd1 vccd1 vccd1 _17319_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18298_ _19473_/A vssd1 vssd1 vccd1 vccd1 _21844_/B sky130_fd_sc_hd__inv_2
XFILLER_0_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17249_ _20909_/B _25862_/Q _25798_/Q vssd1 vssd1 vccd1 vccd1 _17250_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_25_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20260_ _20260_/A _21033_/C vssd1 vssd1 vccd1 vccd1 _20262_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20191_ _26281_/Q hold557/X vssd1 vssd1 vccd1 vccd1 _20191_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_122_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2403 _24029_/X vssd1 vssd1 vccd1 vccd1 _24030_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2414 _15294_/Y vssd1 vssd1 vccd1 vccd1 hold2414/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2425 _26071_/Q vssd1 vssd1 vccd1 vccd1 hold2425/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2436 _26173_/Q vssd1 vssd1 vccd1 vccd1 hold2436/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23950_ hold2180/X _26052_/Q _24001_/S vssd1 vssd1 vccd1 vccd1 _23950_/X sky130_fd_sc_hd__mux2_1
Xhold1702 _20584_/Y vssd1 vssd1 vccd1 vccd1 _25788_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2447 _25451_/Q vssd1 vssd1 vccd1 vccd1 _15380_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2458 _26076_/Q vssd1 vssd1 vccd1 vccd1 hold2458/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1713 _25583_/Q vssd1 vssd1 vccd1 vccd1 _17032_/B sky130_fd_sc_hd__clkbuf_2
Xhold2469 _26049_/Q vssd1 vssd1 vccd1 vccd1 hold2469/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1724 _25607_/Q vssd1 vssd1 vccd1 vccd1 _17356_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1735 _22873_/Y vssd1 vssd1 vccd1 vccd1 _25881_/D sky130_fd_sc_hd__dlygate4sd3_1
X_22901_ _22901_/A _22901_/B vssd1 vssd1 vccd1 vccd1 _22902_/A sky130_fd_sc_hd__nand2_1
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1746 _25603_/Q vssd1 vssd1 vccd1 vccd1 _17312_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23881_ _23881_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23882_/A sky130_fd_sc_hd__and2_1
Xhold1757 _17247_/Y vssd1 vssd1 vccd1 vccd1 _25598_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1768 _25589_/Q vssd1 vssd1 vccd1 vccd1 _17125_/B sky130_fd_sc_hd__buf_2
Xhold1779 _22613_/Y vssd1 vssd1 vccd1 vccd1 _25868_/D sky130_fd_sc_hd__dlygate4sd3_1
X_25620_ _26122_/CLK _25620_/D vssd1 vssd1 vccd1 vccd1 _25620_/Q sky130_fd_sc_hd__dfxtp_4
X_22832_ _22832_/A _22832_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22834_/A sky130_fd_sc_hd__or3_1
XFILLER_0_79_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25551_ _25877_/CLK _25551_/D vssd1 vssd1 vccd1 vccd1 _25551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22763_ _23188_/A _22763_/B vssd1 vssd1 vccd1 vccd1 _22763_/X sky130_fd_sc_hd__or2_1
XFILLER_0_17_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24502_ _24502_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24503_/A sky130_fd_sc_hd__and2_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21714_ _26340_/Q hold425/X vssd1 vssd1 vccd1 vccd1 _21714_/Y sky130_fd_sc_hd__nand2_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25482_ _25933_/CLK hold553/X vssd1 vssd1 vccd1 vccd1 hold551/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22694_ _22694_/A _22694_/B vssd1 vssd1 vccd1 vccd1 _22694_/Y sky130_fd_sc_hd__nand2_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24433_ hold1988/X hold1987/X _24433_/S vssd1 vssd1 vccd1 vccd1 _24434_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_75_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21645_ _21693_/B _21645_/B vssd1 vssd1 vccd1 vccd1 _21646_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_87_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24364_ _24364_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24365_/A sky130_fd_sc_hd__and2_1
XFILLER_0_133_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_50 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21576_ _21628_/B _21579_/A vssd1 vssd1 vccd1 vccd1 _21577_/B sky130_fd_sc_hd__nand2_1
XANTENNA_61 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26103_ _26103_/CLK _26103_/D vssd1 vssd1 vccd1 vccd1 _26103_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_72 _24940_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23315_ _23313_/X hold897/X _12702_/A vssd1 vssd1 vccd1 vccd1 hold898/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20527_ _20527_/A _20527_/B vssd1 vssd1 vccd1 vccd1 _21579_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_162_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24295_ _24295_/A vssd1 vssd1 vccd1 vccd1 _26163_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26034_ _26041_/CLK _26034_/D vssd1 vssd1 vccd1 vccd1 _26034_/Q sky130_fd_sc_hd__dfxtp_1
X_23246_ _23246_/A vssd1 vssd1 vccd1 vccd1 _25912_/D sky130_fd_sc_hd__inv_2
XFILLER_0_120_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20458_ _26288_/Q _20078_/X hold485/X vssd1 vssd1 vccd1 vccd1 _20461_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23177_ _23177_/A _23193_/B _23177_/C vssd1 vssd1 vccd1 vccd1 _23177_/X sky130_fd_sc_hd__and3_1
X_20389_ _20389_/A _22076_/B vssd1 vssd1 vccd1 vccd1 _20390_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22128_ _22128_/A _22808_/A vssd1 vssd1 vccd1 vccd1 _22139_/A sky130_fd_sc_hd__nand2_1
X_14950_ _14950_/A _14950_/B vssd1 vssd1 vccd1 vccd1 _14965_/A sky130_fd_sc_hd__nand2_1
X_22059_ _22057_/Y _22058_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _22059_/Y sky130_fd_sc_hd__a21oi_1
X_13901_ _20233_/B vssd1 vssd1 vccd1 vccd1 _18022_/B sky130_fd_sc_hd__inv_2
X_14881_ _14881_/A _14899_/B vssd1 vssd1 vccd1 vccd1 _14881_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_89_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16620_ _16620_/A _16629_/B _16629_/A vssd1 vssd1 vccd1 vccd1 _16620_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_138_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13832_ _13880_/A hold626/X vssd1 vssd1 vccd1 vccd1 hold627/A sky130_fd_sc_hd__nand2_1
X_25818_ _25835_/CLK _25818_/D vssd1 vssd1 vccd1 vccd1 _25818_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_159_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16551_ _16551_/A _16551_/B vssd1 vssd1 vccd1 vccd1 _16552_/B sky130_fd_sc_hd__nand2_1
X_25749_ _25750_/CLK _25749_/D vssd1 vssd1 vccd1 vccd1 _25749_/Q sky130_fd_sc_hd__dfxtp_1
X_13763_ _18632_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13763_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15502_ _15502_/A _15502_/B vssd1 vssd1 vccd1 vccd1 _15551_/B sky130_fd_sc_hd__nand2_1
X_12714_ _12714_/A _12714_/B hold2010/X vssd1 vssd1 vccd1 vccd1 _12718_/A sky130_fd_sc_hd__or3b_1
X_16482_ _16482_/A _16697_/B vssd1 vssd1 vccd1 vccd1 _16482_/Y sky130_fd_sc_hd__nand2_1
X_19270_ _26224_/Q _12537_/B hold458/X vssd1 vssd1 vccd1 vccd1 _19270_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13694_ _25746_/Q vssd1 vssd1 vccd1 vccd1 _18408_/B sky130_fd_sc_hd__inv_2
XFILLER_0_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15433_ _26023_/Q _25959_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15434_/A sky130_fd_sc_hd__mux2_1
X_18221_ _18221_/A _21019_/B _18221_/C vssd1 vssd1 vccd1 vccd1 _21002_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_183_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12645_ _12645_/A _12645_/B _12645_/C _12645_/D vssd1 vssd1 vccd1 vccd1 _12646_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_150_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15364_ _16813_/B vssd1 vssd1 vccd1 vccd1 _22782_/B sky130_fd_sc_hd__inv_2
XFILLER_0_124_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18152_ _17775_/A _17775_/C _18118_/B vssd1 vssd1 vccd1 vccd1 _18153_/A sky130_fd_sc_hd__a21boi_2
X_12576_ _12576_/A _24836_/B _12582_/A vssd1 vssd1 vccd1 vccd1 _12576_/X sky130_fd_sc_hd__and3_1
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17103_ _19216_/A _17103_/B vssd1 vssd1 vccd1 vccd1 _17456_/A sky130_fd_sc_hd__xor2_4
X_14315_ _14313_/Y hold258/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold259/A sky130_fd_sc_hd__a21oi_1
X_18083_ _18612_/A _19353_/B _18083_/C vssd1 vssd1 vccd1 vccd1 _18084_/C sky130_fd_sc_hd__nand3_1
X_15295_ _15293_/X hold2414/X _15090_/X vssd1 vssd1 vccd1 vccd1 _15295_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17034_ _25584_/Q vssd1 vssd1 vccd1 vccd1 _19115_/B sky130_fd_sc_hd__inv_2
X_14246_ _14264_/A _14246_/B vssd1 vssd1 vccd1 vccd1 _14246_/Y sky130_fd_sc_hd__nand2_1
Xhold309 hold309/A vssd1 vssd1 vccd1 vccd1 hold309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14177_ _25823_/Q vssd1 vssd1 vccd1 vccd1 _18674_/B sky130_fd_sc_hd__inv_2
XFILLER_0_81_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _18178_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13128_/X sky130_fd_sc_hd__or2_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ _18985_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _18985_/Y sky130_fd_sc_hd__nand2_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17936_ _22160_/B _25595_/Q vssd1 vssd1 vccd1 vccd1 _17938_/A sky130_fd_sc_hd__nand2_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _13018_/X _13057_/X _13005_/X _13058_/X vssd1 vssd1 vccd1 vccd1 _13059_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1009 _25083_/Q vssd1 vssd1 vccd1 vccd1 _18373_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17867_ _18252_/A _17867_/B vssd1 vssd1 vccd1 vccd1 _17867_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19606_ _19607_/B _19607_/A vssd1 vssd1 vccd1 vccd1 _19606_/X sky130_fd_sc_hd__or2_1
X_16818_ _16816_/X _16711_/X _16817_/Y _25877_/Q _14170_/X vssd1 vssd1 vccd1 vccd1
+ _16819_/A sky130_fd_sc_hd__a32o_1
X_17798_ _18528_/A _25720_/Q vssd1 vssd1 vccd1 vccd1 _17801_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19537_ _19537_/A _19537_/B vssd1 vssd1 vccd1 vccd1 _19537_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_177_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16749_ _16749_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16749_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19468_ _19465_/Y _19467_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19468_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18419_ _18417_/Y _18418_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25665_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_185_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19399_ _26233_/Q hold455/X vssd1 vssd1 vccd1 vccd1 _19399_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21430_ _21433_/A _21482_/A vssd1 vssd1 vccd1 vccd1 _21432_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_161_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21361_ _21361_/A _21361_/B vssd1 vssd1 vccd1 vccd1 _21362_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23100_ _23091_/Y _23099_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _23100_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_13_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20312_ _20312_/A _25846_/Q vssd1 vssd1 vccd1 vccd1 _20318_/A sky130_fd_sc_hd__nand2_1
X_24080_ hold1/X hold721/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24081_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_4_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold810 hold810/A vssd1 vssd1 vccd1 vccd1 hold810/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21292_ _21294_/B _21294_/C vssd1 vssd1 vccd1 vccd1 _21293_/A sky130_fd_sc_hd__nand2_1
Xhold821 hold821/A vssd1 vssd1 vccd1 vccd1 hold821/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 hold832/A vssd1 vssd1 vccd1 vccd1 hold832/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23031_ _23031_/A _23031_/B _23191_/C vssd1 vssd1 vccd1 vccd1 _23033_/A sky130_fd_sc_hd__or3_1
Xhold843 hold843/A vssd1 vssd1 vccd1 vccd1 hold843/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20243_ _20243_/A _20243_/B vssd1 vssd1 vccd1 vccd1 _20245_/A sky130_fd_sc_hd__nand2_1
Xhold854 hold854/A vssd1 vssd1 vccd1 vccd1 hold854/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 hold865/A vssd1 vssd1 vccd1 vccd1 hold865/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 hold876/A vssd1 vssd1 vccd1 vccd1 hold876/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 hold887/A vssd1 vssd1 vccd1 vccd1 hold887/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 hold898/A vssd1 vssd1 vccd1 vccd1 hold898/X sky130_fd_sc_hd__dlygate4sd3_1
X_20174_ _20174_/A _20174_/B vssd1 vssd1 vccd1 vccd1 _20175_/B sky130_fd_sc_hd__nand2_1
Xhold2200 _23773_/X vssd1 vssd1 vccd1 vccd1 _23774_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2211 _25931_/Q vssd1 vssd1 vccd1 vccd1 _23342_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2222 _26203_/Q vssd1 vssd1 vccd1 vccd1 hold2222/X sky130_fd_sc_hd__dlygate4sd3_1
X_24982_ _24983_/CLK _24982_/D vssd1 vssd1 vccd1 vccd1 _24982_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2233 _26120_/Q vssd1 vssd1 vccd1 vccd1 hold2233/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2244 _25982_/Q vssd1 vssd1 vccd1 vccd1 hold2244/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1510 _23194_/X vssd1 vssd1 vccd1 vccd1 _23195_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2255 _26092_/Q vssd1 vssd1 vccd1 vccd1 hold2255/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1521 _25616_/Q vssd1 vssd1 vccd1 vccd1 _17445_/B sky130_fd_sc_hd__dlygate4sd3_1
X_23933_ _23933_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23934_/A sky130_fd_sc_hd__and2_1
Xhold2266 _24360_/X vssd1 vssd1 vccd1 vccd1 _24361_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1532 _23086_/Y vssd1 vssd1 vccd1 vccd1 _25894_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2277 _26085_/Q vssd1 vssd1 vccd1 vccd1 hold2277/X sky130_fd_sc_hd__buf_1
Xhold2288 _25429_/Q vssd1 vssd1 vccd1 vccd1 _15042_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1543 _25809_/Q vssd1 vssd1 vccd1 vccd1 _21235_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2299 _25452_/Q vssd1 vssd1 vccd1 vccd1 _15394_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1554 _21429_/Y vssd1 vssd1 vccd1 vccd1 _25819_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1565 _20130_/Y vssd1 vssd1 vccd1 vccd1 _25776_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1576 _25898_/Q vssd1 vssd1 vccd1 vccd1 _23149_/B sky130_fd_sc_hd__buf_1
X_23864_ _23864_/A vssd1 vssd1 vccd1 vccd1 _26025_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1587 _21461_/Y vssd1 vssd1 vccd1 vccd1 _25821_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1598 _25584_/Q vssd1 vssd1 vccd1 vccd1 _17048_/B sky130_fd_sc_hd__clkbuf_2
X_25603_ _25604_/CLK _25603_/D vssd1 vssd1 vccd1 vccd1 _25603_/Q sky130_fd_sc_hd__dfxtp_4
X_22815_ _22815_/A _22815_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22817_/A sky130_fd_sc_hd__or3_1
XFILLER_0_79_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23795_ _23795_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23796_/A sky130_fd_sc_hd__and2_1
XFILLER_0_95_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25534_ _25534_/CLK hold949/X vssd1 vssd1 vccd1 vccd1 hold948/A sky130_fd_sc_hd__dfxtp_1
X_22746_ _22746_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22746_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_55_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xascon_wrapper_12 vssd1 vssd1 vccd1 vccd1 ascon_wrapper_12/HI io_oeb[9] sky130_fd_sc_hd__conb_1
XFILLER_0_164_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25465_ _26069_/CLK _25465_/D vssd1 vssd1 vccd1 vccd1 _25465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22677_ _22677_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _22677_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_165_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24416_ _24416_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24417_/A sky130_fd_sc_hd__and2_1
XFILLER_0_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21628_ _21676_/B _21628_/B vssd1 vssd1 vccd1 vccd1 _21630_/A sky130_fd_sc_hd__nand2_1
X_25396_ _26207_/CLK _25396_/D vssd1 vssd1 vccd1 vccd1 _25396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24347_ hold2334/X hold2016/X _24356_/S vssd1 vssd1 vccd1 vccd1 _24348_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21559_ _21562_/A _21612_/A vssd1 vssd1 vccd1 vccd1 _21561_/A sky130_fd_sc_hd__nand2_1
X_14100_ _14118_/A hold794/X vssd1 vssd1 vccd1 vccd1 _14100_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15080_ _15080_/A _15085_/B vssd1 vssd1 vccd1 vccd1 _15080_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_160_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24278_ _24278_/A vssd1 vssd1 vccd1 vccd1 _26158_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26017_ _26021_/CLK _26017_/D vssd1 vssd1 vccd1 vccd1 _26017_/Q sky130_fd_sc_hd__dfxtp_1
X_14031_ hold438/X _14030_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold439/A sky130_fd_sc_hd__a21oi_1
X_23229_ _23229_/A vssd1 vssd1 vccd1 vccd1 _25909_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18770_ _18793_/A _25764_/Q _18891_/C vssd1 vssd1 vccd1 vccd1 _18771_/C sky130_fd_sc_hd__nand3_1
X_15982_ hold771/X vssd1 vssd1 vccd1 vccd1 _15985_/B sky130_fd_sc_hd__inv_2
X_17721_ _17721_/A _17721_/B vssd1 vssd1 vccd1 vccd1 _17829_/A sky130_fd_sc_hd__nand2_1
X_14933_ _14925_/A _14925_/B _14923_/Y _14924_/A vssd1 vssd1 vccd1 vccd1 _14933_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17652_ _17652_/A _17652_/B vssd1 vssd1 vccd1 vccd1 _17652_/X sky130_fd_sc_hd__xor2_1
X_14864_ _14864_/A _14864_/B vssd1 vssd1 vccd1 vccd1 _14864_/Y sky130_fd_sc_hd__nand2_1
X_16603_ _16650_/A vssd1 vssd1 vccd1 vccd1 _16610_/B sky130_fd_sc_hd__inv_2
XFILLER_0_138_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13815_ _18793_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13815_/Y sky130_fd_sc_hd__nor2_1
X_14795_ _14900_/A _14795_/B vssd1 vssd1 vccd1 vccd1 _14795_/Y sky130_fd_sc_hd__nand2_1
X_17583_ _17605_/A _17583_/B vssd1 vssd1 vccd1 vccd1 _17583_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19322_ _19322_/A _19322_/B vssd1 vssd1 vccd1 vccd1 _19322_/Y sky130_fd_sc_hd__nand2_1
X_16534_ _16534_/A _16539_/B vssd1 vssd1 vccd1 vccd1 _16535_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_85_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13746_ _13823_/A _13746_/B vssd1 vssd1 vccd1 vccd1 _13746_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_168_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19253_ _19248_/X _18879_/X _19252_/X vssd1 vssd1 vccd1 vccd1 _19254_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16465_ _16466_/B _16466_/A vssd1 vssd1 vccd1 vccd1 _16492_/A sky130_fd_sc_hd__or2_1
X_13677_ _26246_/Q _13612_/X _13605_/X _13676_/Y vssd1 vssd1 vccd1 vccd1 _13678_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18204_ _20973_/B _21974_/A vssd1 vssd1 vccd1 vccd1 _20964_/A sky130_fd_sc_hd__nand2_2
X_15416_ _15416_/A vssd1 vssd1 vccd1 vccd1 _15425_/B sky130_fd_sc_hd__inv_2
X_12628_ _12628_/A _12645_/A vssd1 vssd1 vccd1 vccd1 _12628_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16396_ _16393_/A _16393_/B _16416_/B _16395_/Y vssd1 vssd1 vccd1 vccd1 _16396_/X
+ sky130_fd_sc_hd__a31o_1
X_19184_ _19182_/X _19183_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19184_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15347_ _15347_/A vssd1 vssd1 vccd1 vccd1 _15356_/B sky130_fd_sc_hd__inv_2
XFILLER_0_14_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18135_ _18446_/A _19467_/B _21716_/A vssd1 vssd1 vccd1 vccd1 _18136_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_170_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12559_ _12559_/A hold4/X vssd1 vssd1 vccd1 vccd1 _12564_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15278_ _15307_/B _15827_/A vssd1 vssd1 vccd1 vccd1 _15278_/X sky130_fd_sc_hd__or2_1
Xhold106 hold106/A vssd1 vssd1 vccd1 vccd1 hold106/X sky130_fd_sc_hd__dlygate4sd3_1
X_18066_ _25844_/Q vssd1 vssd1 vccd1 vccd1 _20251_/B sky130_fd_sc_hd__inv_2
XFILLER_0_151_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold117 hold117/A vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold128 hold128/A vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ hold567/X _14228_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold568/A sky130_fd_sc_hd__a21oi_1
X_17017_ _17012_/Y _17016_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _17017_/Y sky130_fd_sc_hd__a21oi_1
Xhold139 hold139/A vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18968_ _19026_/A _18968_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18968_/X sky130_fd_sc_hd__and3_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ _19138_/B _25649_/Q vssd1 vssd1 vccd1 vccd1 _17923_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18899_ _18899_/A _18899_/B vssd1 vssd1 vccd1 vccd1 _18899_/X sky130_fd_sc_hd__xor2_1
X_20930_ _21042_/A _20930_/B _20929_/X vssd1 vssd1 vccd1 vccd1 _20931_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20861_ _20863_/B _20863_/C vssd1 vssd1 vccd1 vccd1 _20862_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22600_ _22600_/A _22600_/B vssd1 vssd1 vccd1 vccd1 _22601_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_117_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23580_ _24870_/B _23532_/X _23579_/X vssd1 vssd1 vccd1 vccd1 _23581_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_159_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20792_ _20795_/A _20795_/C vssd1 vssd1 vccd1 vccd1 _20793_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22531_ _22531_/A _23001_/B _22531_/C vssd1 vssd1 vccd1 vccd1 _22531_/X sky130_fd_sc_hd__and3_1
XFILLER_0_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25250_ _26340_/CLK hold400/X vssd1 vssd1 vccd1 vccd1 hold398/A sky130_fd_sc_hd__dfxtp_1
X_22462_ _22462_/A _25891_/Q vssd1 vssd1 vccd1 vccd1 _22462_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24201_ _24201_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24202_/A sky130_fd_sc_hd__and2_1
XFILLER_0_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21413_ _21411_/Y _21412_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21413_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25181_ _25761_/CLK hold523/X vssd1 vssd1 vccd1 vccd1 hold521/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22393_ _22393_/A _22393_/B vssd1 vssd1 vccd1 vccd1 _22393_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_115_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24132_ _24132_/A vssd1 vssd1 vccd1 vccd1 _26110_/D sky130_fd_sc_hd__clkbuf_1
X_21344_ _21636_/A _21344_/B _21343_/X vssd1 vssd1 vccd1 vccd1 _21345_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_103_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24063_ _24063_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24064_/A sky130_fd_sc_hd__and2_1
XFILLER_0_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold640 hold640/A vssd1 vssd1 vccd1 vccd1 hold640/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21275_ _21694_/B _21643_/C vssd1 vssd1 vccd1 vccd1 _21276_/B sky130_fd_sc_hd__nand2_1
Xhold651 hold651/A vssd1 vssd1 vccd1 vccd1 hold651/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 hold662/A vssd1 vssd1 vccd1 vccd1 hold662/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23014_ _26073_/Q vssd1 vssd1 vccd1 vccd1 _23015_/A sky130_fd_sc_hd__inv_2
X_20226_ _20226_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20231_/A sky130_fd_sc_hd__nand2_1
Xhold673 hold673/A vssd1 vssd1 vccd1 vccd1 hold673/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold684 hold684/A vssd1 vssd1 vccd1 vccd1 hold684/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 hold695/A vssd1 vssd1 vccd1 vccd1 hold695/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_25_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20157_ _21042_/A _20157_/B _20156_/X vssd1 vssd1 vccd1 vccd1 _20158_/B sky130_fd_sc_hd__or3b_1
Xhold2030 _23375_/X vssd1 vssd1 vccd1 vccd1 _23377_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2041 _15360_/X vssd1 vssd1 vccd1 vccd1 hold2041/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2052 _23844_/X vssd1 vssd1 vccd1 vccd1 _23845_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2063 _25415_/Q vssd1 vssd1 vccd1 vccd1 _14923_/B sky130_fd_sc_hd__dlygate4sd3_1
X_24965_ _25418_/CLK _24965_/D vssd1 vssd1 vccd1 vccd1 _24965_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2074 _26001_/Q vssd1 vssd1 vccd1 vccd1 _14875_/B sky130_fd_sc_hd__buf_1
X_20088_ _20088_/A _20088_/B vssd1 vssd1 vccd1 vccd1 _20092_/A sky130_fd_sc_hd__nand2_1
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2085 _25966_/Q vssd1 vssd1 vccd1 vccd1 hold2085/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1340 _13059_/X vssd1 vssd1 vccd1 vccd1 _25061_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2096 _26087_/Q vssd1 vssd1 vccd1 vccd1 hold2096/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1351 _25733_/Q vssd1 vssd1 vccd1 vccd1 _19452_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23916_ _23916_/A vssd1 vssd1 vccd1 vccd1 _26042_/D sky130_fd_sc_hd__clkbuf_1
Xhold1362 _14769_/Y vssd1 vssd1 vccd1 vccd1 _25396_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24896_ _15761_/B _15780_/B _24945_/S vssd1 vssd1 vccd1 vccd1 _24896_/X sky130_fd_sc_hd__mux2_1
Xhold1373 _25394_/Q vssd1 vssd1 vccd1 vccd1 _14750_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1384 _15785_/Y vssd1 vssd1 vccd1 vccd1 _25473_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1395 _25769_/Q vssd1 vssd1 vccd1 vccd1 _19953_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23847_ hold2167/X hold1928/X _23907_/S vssd1 vssd1 vccd1 vccd1 _23848_/A sky130_fd_sc_hd__mux2_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _18002_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13600_/Y sky130_fd_sc_hd__nor2_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _14578_/Y hold360/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold361/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23778_ _23778_/A vssd1 vssd1 vccd1 vccd1 _25997_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13531_ _25720_/Q vssd1 vssd1 vccd1 vccd1 _17800_/B sky130_fd_sc_hd__inv_2
XFILLER_0_95_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25517_ _25537_/CLK hold967/X vssd1 vssd1 vccd1 vccd1 hold966/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22729_ _22729_/A _22729_/B vssd1 vssd1 vccd1 vccd1 _22730_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_138_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16250_ _16250_/A _16250_/B vssd1 vssd1 vccd1 vccd1 _16251_/B sky130_fd_sc_hd__nand2_1
X_25448_ _25511_/CLK hold976/X vssd1 vssd1 vccd1 vccd1 hold975/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13462_ _13522_/A _13460_/X _23629_/B _13461_/X vssd1 vssd1 vccd1 vccd1 _13462_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15201_ _15188_/X _15268_/B _15200_/Y vssd1 vssd1 vccd1 vccd1 _15201_/Y sky130_fd_sc_hd__o21ai_1
X_16181_ _16181_/A vssd1 vssd1 vccd1 vccd1 _16189_/A sky130_fd_sc_hd__inv_2
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25379_ _26205_/CLK hold394/X vssd1 vssd1 vccd1 vccd1 hold392/A sky130_fd_sc_hd__dfxtp_1
X_13393_ _18998_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13393_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15132_ _15129_/Y _15131_/Y _15090_/X vssd1 vssd1 vccd1 vccd1 hold932/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15063_ _15061_/X hold2453/X _14928_/X vssd1 vssd1 vccd1 vccd1 _15063_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19940_ _19938_/X _19939_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19940_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14014_ _14118_/A hold503/X vssd1 vssd1 vccd1 vccd1 hold504/A sky130_fd_sc_hd__nand2_1
XFILLER_0_103_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19871_ _20790_/A _22615_/B _25641_/Q vssd1 vssd1 vccd1 vccd1 _20795_/C sky130_fd_sc_hd__nand3_1
X_18822_ _18986_/A _19588_/A vssd1 vssd1 vccd1 vccd1 _18822_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18753_ _18955_/A _18753_/B _18894_/C vssd1 vssd1 vccd1 vccd1 _18754_/C sky130_fd_sc_hd__nand3_1
X_15965_ _16231_/A vssd1 vssd1 vccd1 vccd1 _16212_/A sky130_fd_sc_hd__clkbuf_8
X_17704_ _17704_/A vssd1 vssd1 vccd1 vccd1 _17705_/C sky130_fd_sc_hd__inv_2
X_14916_ _14916_/A _14916_/B vssd1 vssd1 vccd1 vccd1 _14917_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18684_ _19744_/A vssd1 vssd1 vccd1 vccd1 _22391_/B sky130_fd_sc_hd__inv_2
X_15896_ _15884_/C _15894_/B _15882_/A vssd1 vssd1 vccd1 vccd1 _15896_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17635_ _18252_/A _17635_/B vssd1 vssd1 vccd1 vccd1 _17635_/Y sky130_fd_sc_hd__nand2_1
X_14847_ _25854_/Q _14170_/A _15027_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14848_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17566_ _17566_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17566_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_81_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14778_ _14776_/Y _14777_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14778_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19305_ _20740_/A _19303_/Y _20745_/C vssd1 vssd1 vccd1 vccd1 _19393_/B sky130_fd_sc_hd__o21a_1
X_16517_ _16698_/A hold940/X vssd1 vssd1 vccd1 vccd1 _16517_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13729_ hold516/X _13728_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold517/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17497_ _17495_/Y _17496_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _25623_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19236_ _20986_/A vssd1 vssd1 vccd1 vccd1 _19236_/X sky130_fd_sc_hd__buf_12
X_16448_ _16473_/A hold866/X vssd1 vssd1 vccd1 vccd1 _16448_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_128_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19167_ _19167_/A _19972_/B vssd1 vssd1 vccd1 vccd1 _19167_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_82_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16379_ _16379_/A _16379_/B vssd1 vssd1 vccd1 vccd1 _16380_/A sky130_fd_sc_hd__and2_1
XFILLER_0_6_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18118_ _18118_/A _18118_/B vssd1 vssd1 vccd1 vccd1 _18119_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_182_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19098_ _20247_/A _21958_/A _25588_/Q vssd1 vssd1 vccd1 vccd1 _20251_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_83_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18049_ _18792_/A _25732_/Q vssd1 vssd1 vccd1 vccd1 _18053_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21060_ _21561_/C _21516_/B vssd1 vssd1 vccd1 vccd1 _21062_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20011_ _20011_/A _20011_/B vssd1 vssd1 vccd1 vccd1 _20014_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_39_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24750_ _24750_/A vssd1 vssd1 vccd1 vccd1 _26311_/D sky130_fd_sc_hd__clkbuf_1
X_21962_ _21962_/A _21962_/B _22994_/A vssd1 vssd1 vccd1 vccd1 _21962_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23701_ _23701_/A vssd1 vssd1 vccd1 vccd1 _25972_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20913_ _20913_/A _21909_/B _20913_/C vssd1 vssd1 vccd1 vccd1 _20916_/C sky130_fd_sc_hd__nand3_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24681_ _24681_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24682_/A sky130_fd_sc_hd__and2_1
X_21893_ _21893_/A _21893_/B _22960_/A vssd1 vssd1 vccd1 vccd1 _21893_/Y sky130_fd_sc_hd__nand3_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23632_ _24560_/A vssd1 vssd1 vccd1 vccd1 _23721_/B sky130_fd_sc_hd__buf_6
XFILLER_0_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20844_ _20844_/A _21387_/B _20844_/C vssd1 vssd1 vccd1 vccd1 _20845_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_138_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23563_ hold38/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23563_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20775_ _20775_/A _20775_/B vssd1 vssd1 vccd1 vccd1 _20776_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25302_ _26136_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__dfxtp_1
X_22514_ _18796_/A _25829_/Q _22512_/Y _22513_/Y vssd1 vssd1 vccd1 vccd1 _22515_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26282_ _26283_/CLK _26282_/D vssd1 vssd1 vccd1 vccd1 _26282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23494_ _24944_/S hold89/A _23493_/X vssd1 vssd1 vccd1 vccd1 _23494_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25233_ _25687_/CLK hold589/X vssd1 vssd1 vccd1 vccd1 hold587/A sky130_fd_sc_hd__dfxtp_1
X_22445_ _22859_/A _23008_/B vssd1 vssd1 vccd1 vccd1 _22446_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25164_ _25781_/CLK hold616/X vssd1 vssd1 vccd1 vccd1 hold614/A sky130_fd_sc_hd__dfxtp_1
X_22376_ _22376_/A _22376_/B vssd1 vssd1 vccd1 vccd1 _22958_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_32_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24115_ _24115_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24116_/A sky130_fd_sc_hd__and2_1
X_21327_ _21326_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21327_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_128_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25095_ _26308_/CLK _25095_/D vssd1 vssd1 vccd1 vccd1 _25095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_4__f_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _25184_/CLK sky130_fd_sc_hd__clkbuf_16
X_24046_ _24046_/A vssd1 vssd1 vccd1 vccd1 _26083_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21258_ _21636_/A _21258_/B _21257_/X vssd1 vssd1 vccd1 vccd1 _21259_/B sky130_fd_sc_hd__or3b_1
Xhold470 hold470/A vssd1 vssd1 vccd1 vccd1 hold470/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 hold481/A vssd1 vssd1 vccd1 vccd1 hold481/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 hold492/A vssd1 vssd1 vccd1 vccd1 hold492/X sky130_fd_sc_hd__dlygate4sd3_1
X_20209_ _20209_/A _20209_/B vssd1 vssd1 vccd1 vccd1 _21450_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_159_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21189_ _21189_/A _21189_/B vssd1 vssd1 vccd1 vccd1 _21191_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25997_ _25998_/CLK _25997_/D vssd1 vssd1 vccd1 vccd1 _25997_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _15750_/A _15750_/B vssd1 vssd1 vccd1 vccd1 _15750_/Y sky130_fd_sc_hd__nand2_1
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ _12891_/X _14419_/A _12909_/X _25623_/Q vssd1 vssd1 vccd1 vccd1 _12962_/X
+ sky130_fd_sc_hd__a22o_1
X_24948_ _24867_/S _24941_/Y _24943_/Y _24947_/X vssd1 vssd1 vccd1 vccd1 _24948_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_172_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1170 _13071_/X vssd1 vssd1 vccd1 vccd1 _25063_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ _14701_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14701_/Y sky130_fd_sc_hd__nand2_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1181 _25048_/Q vssd1 vssd1 vccd1 vccd1 _17529_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1192 _19411_/Y vssd1 vssd1 vccd1 vccd1 _25730_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15681_ _16933_/B vssd1 vssd1 vccd1 vccd1 _23079_/B sky130_fd_sc_hd__inv_2
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _12891_/X _14376_/A _12752_/X _25610_/Q vssd1 vssd1 vccd1 vccd1 _12893_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24879_ _24879_/A _24957_/S vssd1 vssd1 vccd1 vccd1 _24879_/Y sky130_fd_sc_hd__nand2_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _20011_/B _25877_/Q _25813_/Q vssd1 vssd1 vccd1 vccd1 _17421_/B sky130_fd_sc_hd__mux2_2
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _14632_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14632_/Y sky130_fd_sc_hd__nand2_1
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _17542_/A _17594_/A vssd1 vssd1 vccd1 vccd1 _17352_/B sky130_fd_sc_hd__xnor2_1
X_14563_ _14563_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14563_/Y sky130_fd_sc_hd__nand2_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _16300_/X _16301_/Y _16076_/X vssd1 vssd1 vccd1 vccd1 _25509_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13514_ _13583_/A _13514_/B vssd1 vssd1 vccd1 vccd1 _13514_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_137_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17282_ _17393_/A _17282_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17282_/X sky130_fd_sc_hd__and3_1
X_14494_ _14494_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14494_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_153_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19021_ _19021_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _19021_/Y sky130_fd_sc_hd__nand2_1
X_16233_ _16230_/X _16232_/Y _16076_/X vssd1 vssd1 vccd1 vccd1 _25504_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_181_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13445_ _26209_/Q _13426_/X _13444_/X vssd1 vssd1 vccd1 vccd1 _13445_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_64_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16164_ hold754/X vssd1 vssd1 vccd1 vccd1 _16168_/B sky130_fd_sc_hd__inv_2
XFILLER_0_153_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13376_ _13315_/X _13374_/X _13300_/X _13375_/X vssd1 vssd1 vccd1 vccd1 _13376_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15115_ _15115_/A _15810_/B vssd1 vssd1 vccd1 vccd1 _15116_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_23_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16095_ _16095_/A _16095_/B vssd1 vssd1 vccd1 vccd1 _16096_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_121_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15046_ _15046_/A _15051_/B vssd1 vssd1 vccd1 vccd1 _15046_/Y sky130_fd_sc_hd__nand2_1
X_19923_ _19923_/A _19980_/B _19923_/C vssd1 vssd1 vccd1 vccd1 _19923_/X sky130_fd_sc_hd__and3_1
XFILLER_0_167_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19854_ _26265_/Q hold733/X vssd1 vssd1 vccd1 vccd1 _19854_/Y sky130_fd_sc_hd__nand2_1
X_18805_ _22539_/B _25638_/Q vssd1 vssd1 vccd1 vccd1 _18807_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19785_ _26260_/Q hold671/X vssd1 vssd1 vccd1 vccd1 _19785_/Y sky130_fd_sc_hd__nand2_1
X_16997_ _17794_/A vssd1 vssd1 vccd1 vccd1 _18529_/C sky130_fd_sc_hd__buf_8
XFILLER_0_183_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18736_ _18736_/A _20517_/A vssd1 vssd1 vccd1 vccd1 _19003_/A sky130_fd_sc_hd__xor2_4
X_15948_ _16401_/C vssd1 vssd1 vccd1 vccd1 _16691_/B sky130_fd_sc_hd__buf_8
X_18667_ _18667_/A _18667_/B vssd1 vssd1 vccd1 vccd1 _22369_/A sky130_fd_sc_hd__nand2_1
X_15879_ _21830_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _15881_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_116_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17618_ _17616_/X _17528_/X _17617_/X vssd1 vssd1 vccd1 vccd1 _17619_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_116_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18598_ _18596_/X _18269_/X _18597_/X vssd1 vssd1 vccd1 vccd1 _18600_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_93_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17549_ _17549_/A _17549_/B vssd1 vssd1 vccd1 vccd1 _17549_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_86_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20560_ _20560_/A _25891_/Q vssd1 vssd1 vccd1 vccd1 _20566_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_117_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19219_ _19234_/A _19308_/B vssd1 vssd1 vccd1 vccd1 _19220_/B sky130_fd_sc_hd__xor2_1
X_20491_ _21562_/A _21279_/B vssd1 vssd1 vccd1 vccd1 _20492_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_15_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22230_ _22561_/A _22230_/B vssd1 vssd1 vccd1 vccd1 _22230_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_104_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22161_ _17947_/A _25787_/Q _22159_/Y _22160_/Y vssd1 vssd1 vccd1 vccd1 _22162_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21112_ _21594_/C vssd1 vssd1 vccd1 vccd1 _21597_/B sky130_fd_sc_hd__inv_2
X_22092_ _22090_/X _15839_/B _22091_/Y _14804_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _22093_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_125_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_207_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _25596_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25920_ _25925_/CLK _25920_/D vssd1 vssd1 vccd1 vccd1 _25920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21043_ _21043_/A _21043_/B vssd1 vssd1 vccd1 vccd1 _21044_/A sky130_fd_sc_hd__nand2_1
X_25851_ _26207_/CLK _25851_/D vssd1 vssd1 vccd1 vccd1 _25851_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_157_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24802_ hold2714/X hold2712/X _24817_/S vssd1 vssd1 vccd1 vccd1 _24803_/A sky130_fd_sc_hd__mux2_1
X_22994_ _22994_/A _22994_/B vssd1 vssd1 vccd1 vccd1 _22995_/A sky130_fd_sc_hd__xor2_1
Xclkbuf_4_12__f_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_82_clk/A
+ sky130_fd_sc_hd__clkbuf_16
X_25782_ _26286_/CLK _25782_/D vssd1 vssd1 vccd1 vccd1 _25782_/Q sky130_fd_sc_hd__dfxtp_2
X_21945_ _23152_/A vssd1 vssd1 vccd1 vccd1 _23151_/A sky130_fd_sc_hd__inv_2
X_24733_ _24733_/A vssd1 vssd1 vccd1 vccd1 _26306_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24664_ hold2718/X hold2372/X _24664_/S vssd1 vssd1 vccd1 vccd1 _24665_/A sky130_fd_sc_hd__mux2_1
X_21876_ _23120_/A vssd1 vssd1 vccd1 vccd1 _23119_/A sky130_fd_sc_hd__inv_2
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23615_ _23615_/A vssd1 vssd1 vccd1 vccd1 _25944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20827_ _21435_/B vssd1 vssd1 vccd1 vccd1 _21432_/C sky130_fd_sc_hd__inv_2
XFILLER_0_65_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24595_ _24595_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24596_/A sky130_fd_sc_hd__and2_1
XFILLER_0_181_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26334_ _26334_/CLK _26334_/D vssd1 vssd1 vccd1 vccd1 _26334_/Q sky130_fd_sc_hd__dfxtp_2
X_23546_ hold149/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23546_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_108_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20758_ _20758_/A _20758_/B vssd1 vssd1 vccd1 vccd1 _20760_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_80_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26265_ _26273_/CLK _26265_/D vssd1 vssd1 vccd1 vccd1 _26265_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23477_ hold59/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23477_/X sky130_fd_sc_hd__or2b_1
X_20689_ _20689_/A _21322_/B _20689_/C vssd1 vssd1 vccd1 vccd1 _20690_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_162_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25216_ _26303_/CLK hold580/X vssd1 vssd1 vccd1 vccd1 hold578/A sky130_fd_sc_hd__dfxtp_1
X_13230_ _26174_/Q _13065_/X _13229_/X vssd1 vssd1 vccd1 vccd1 _13230_/X sky130_fd_sc_hd__a21o_1
X_22428_ _22423_/B _22421_/X _22427_/X vssd1 vssd1 vccd1 vccd1 _22429_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_17_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26196_ _26198_/CLK _26196_/D vssd1 vssd1 vccd1 vccd1 _26196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25147_ _25727_/CLK hold788/X vssd1 vssd1 vccd1 vccd1 hold786/A sky130_fd_sc_hd__dfxtp_1
X_13161_ _26163_/Q _13065_/X _13160_/X vssd1 vssd1 vccd1 vccd1 _13161_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_62_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22359_ _22359_/A _23071_/A _22359_/C vssd1 vssd1 vccd1 vccd1 _22359_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_62_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25078_ _26289_/CLK _25078_/D vssd1 vssd1 vccd1 vccd1 _25078_/Q sky130_fd_sc_hd__dfxtp_1
X_13092_ _13018_/X _13090_/X _13005_/X _13091_/X vssd1 vssd1 vccd1 vccd1 _13092_/X
+ sky130_fd_sc_hd__o211a_1
X_16920_ _23047_/B _16773_/A _16916_/Y _16919_/Y _14345_/A vssd1 vssd1 vccd1 vccd1
+ _16920_/Y sky130_fd_sc_hd__a221oi_1
X_24029_ hold2402/X _26078_/Q _24047_/S vssd1 vssd1 vccd1 vccd1 _24029_/X sky130_fd_sc_hd__mux2_1
X_16851_ _16858_/A _16851_/B vssd1 vssd1 vccd1 vccd1 _16851_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_189_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15802_ _15789_/Y _15830_/B _15801_/Y vssd1 vssd1 vccd1 vccd1 _15802_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_176_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19570_ _26245_/Q _19483_/X hold791/X vssd1 vssd1 vccd1 vccd1 _19570_/Y sky130_fd_sc_hd__a21oi_1
X_16782_ _15302_/A _16781_/Y _15621_/A vssd1 vssd1 vccd1 vccd1 _16782_/Y sky130_fd_sc_hd__a21oi_1
X_13994_ _14000_/A hold623/X vssd1 vssd1 vccd1 vccd1 hold624/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18521_ _22179_/B _25624_/Q vssd1 vssd1 vccd1 vccd1 _18523_/A sky130_fd_sc_hd__nand2_1
X_15733_ _15720_/X _15764_/A _15732_/Y vssd1 vssd1 vccd1 vccd1 _15733_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _12930_/X _12943_/X _12917_/X _12944_/X vssd1 vssd1 vccd1 vccd1 _12945_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ _18452_/A _21290_/A vssd1 vssd1 vccd1 vccd1 _18798_/A sky130_fd_sc_hd__xor2_4
X_15664_ _25467_/Q vssd1 vssd1 vccd1 vccd1 _15673_/B sky130_fd_sc_hd__inv_2
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _26238_/Q _25607_/Q vssd1 vssd1 vccd1 vccd1 _14367_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_73_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17403_ _19082_/A vssd1 vssd1 vccd1 vccd1 _17624_/A sky130_fd_sc_hd__buf_6
XFILLER_0_28_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14615_ _14645_/A hold74/X vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__nand2_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _18445_/A _18387_/B vssd1 vssd1 vccd1 vccd1 _18385_/A sky130_fd_sc_hd__nand2_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _16900_/B vssd1 vssd1 vccd1 vccd1 _22999_/B sky130_fd_sc_hd__inv_2
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17334_ _17331_/X _17241_/X _17333_/X vssd1 vssd1 vccd1 vccd1 _17335_/A sky130_fd_sc_hd__a21o_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14546_ _14585_/A hold128/X vssd1 vssd1 vccd1 vccd1 hold129/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17265_ _20791_/B _25897_/Q _25833_/Q vssd1 vssd1 vccd1 vccd1 _17266_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_83_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14477_ _14525_/A hold68/X vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__nand2_1
XFILLER_0_114_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19004_ _19053_/A _19004_/B vssd1 vssd1 vccd1 vccd1 _19004_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16216_ _16216_/A _16271_/B vssd1 vssd1 vccd1 vccd1 _16227_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_141_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13428_ _26334_/Q _19844_/A vssd1 vssd1 vccd1 vccd1 _14669_/A sky130_fd_sc_hd__xor2_1
X_17196_ _20597_/B _25892_/Q _25828_/Q vssd1 vssd1 vccd1 vccd1 _17197_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_141_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16147_ hold861/X _16148_/A vssd1 vssd1 vccd1 vccd1 _16149_/A sky130_fd_sc_hd__or2_1
XFILLER_0_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13359_ _13359_/A vssd1 vssd1 vccd1 vccd1 _19687_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16078_ hold763/X vssd1 vssd1 vccd1 vccd1 _16081_/B sky130_fd_sc_hd__inv_2
X_15029_ _15029_/A _15034_/B vssd1 vssd1 vccd1 vccd1 _15030_/B sky130_fd_sc_hd__nor2_1
X_19906_ _26269_/Q hold803/X vssd1 vssd1 vccd1 vccd1 _19906_/Y sky130_fd_sc_hd__nand2_1
Xhold2607 _24461_/X vssd1 vssd1 vccd1 vccd1 _24462_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2618 _26337_/Q vssd1 vssd1 vccd1 vccd1 hold2618/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2629 _24658_/X vssd1 vssd1 vccd1 vccd1 _24659_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1906 _23739_/X vssd1 vssd1 vccd1 vccd1 _23740_/A sky130_fd_sc_hd__dlygate4sd3_1
X_19837_ _19829_/X _19836_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19837_/Y sky130_fd_sc_hd__o21ai_1
Xhold1917 _23250_/Y vssd1 vssd1 vccd1 vccd1 _25913_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1928 _26020_/Q vssd1 vssd1 vccd1 vccd1 hold1928/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1939 _24440_/X vssd1 vssd1 vccd1 vccd1 _24441_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput2 io_in[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19768_ _19975_/A _19768_/B vssd1 vssd1 vccd1 vccd1 _19768_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_155_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18719_ _19026_/A _18719_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18719_/X sky130_fd_sc_hd__and3_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19699_ _19698_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19700_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_151_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21730_ _17911_/A _25793_/Q _21728_/Y _21729_/Y vssd1 vssd1 vccd1 vccd1 _21731_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_176_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21661_ _21709_/B _21661_/B vssd1 vssd1 vccd1 vccd1 _21662_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_188_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23400_ _23397_/Y _23399_/Y _24858_/S vssd1 vssd1 vccd1 vccd1 _23400_/X sky130_fd_sc_hd__mux2_1
X_20612_ _21335_/C _21612_/A vssd1 vssd1 vccd1 vccd1 _20613_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_164_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24380_ _24380_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24381_/A sky130_fd_sc_hd__and2_1
X_21592_ _21644_/B _21596_/A vssd1 vssd1 vccd1 vccd1 _21594_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23331_ _23334_/A _23377_/B _23331_/C vssd1 vssd1 vccd1 vccd1 _23332_/A sky130_fd_sc_hd__and3_1
XFILLER_0_156_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20543_ _20543_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _20543_/Y sky130_fd_sc_hd__nand2_1
X_26050_ _26051_/CLK _26050_/D vssd1 vssd1 vccd1 vccd1 _26050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23262_ _23262_/A vssd1 vssd1 vccd1 vccd1 _25914_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20474_ _20474_/A _20474_/B vssd1 vssd1 vccd1 vccd1 _20476_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_131_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25001_ _25865_/CLK _25001_/D vssd1 vssd1 vccd1 vccd1 _25001_/Q sky130_fd_sc_hd__dfxtp_1
X_22213_ _22213_/A _22872_/B vssd1 vssd1 vccd1 vccd1 _22214_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_104_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23193_ _23193_/A _23193_/B _23193_/C vssd1 vssd1 vccd1 vccd1 _23193_/X sky130_fd_sc_hd__and3_1
XFILLER_0_42_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22144_ _22653_/A _22144_/B vssd1 vssd1 vccd1 vccd1 _22144_/X sky130_fd_sc_hd__or2_1
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22075_ _22075_/A _25848_/Q vssd1 vssd1 vccd1 vccd1 _22075_/Y sky130_fd_sc_hd__nand2_1
X_25903_ _26269_/CLK _25903_/D vssd1 vssd1 vccd1 vccd1 _25903_/Q sky130_fd_sc_hd__dfxtp_2
X_21026_ _21028_/B _21028_/C vssd1 vssd1 vccd1 vccd1 _21027_/A sky130_fd_sc_hd__nand2_1
X_25834_ _25865_/CLK _25834_/D vssd1 vssd1 vccd1 vccd1 _25834_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_57_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22977_ _22977_/A _22977_/B vssd1 vssd1 vccd1 vccd1 _22978_/A sky130_fd_sc_hd__xor2_1
X_25765_ _25765_/CLK _25765_/D vssd1 vssd1 vccd1 vccd1 _25765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _13518_/B _26085_/Q vssd1 vssd1 vccd1 vccd1 _12730_/Y sky130_fd_sc_hd__nand2_1
X_24716_ hold2667/X hold2594/X _24740_/S vssd1 vssd1 vccd1 vccd1 _24717_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_179_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21928_ _21928_/A _21928_/B _22977_/A vssd1 vssd1 vccd1 vccd1 _21928_/Y sky130_fd_sc_hd__nand3_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25696_ _26324_/CLK _25696_/D vssd1 vssd1 vccd1 vccd1 _25696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12664_/A _12661_/B _24983_/Q vssd1 vssd1 vccd1 vccd1 _12662_/C sky130_fd_sc_hd__or3b_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21859_ _21859_/A _21859_/B _22943_/A vssd1 vssd1 vccd1 vccd1 _21859_/Y sky130_fd_sc_hd__nand3_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24647_ _24647_/A vssd1 vssd1 vccd1 vccd1 _26278_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _14400_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14400_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_132_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15380_ _15380_/A vssd1 vssd1 vccd1 vccd1 _15387_/B sky130_fd_sc_hd__inv_2
X_12592_ _12646_/A _24836_/B _12592_/C vssd1 vssd1 vccd1 vccd1 _12593_/A sky130_fd_sc_hd__and3_1
XFILLER_0_148_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24578_ hold2708/X hold2707/X _24587_/S vssd1 vssd1 vccd1 vccd1 _24579_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_107_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14331_ _14331_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14331_/Y sky130_fd_sc_hd__nand2_1
X_26317_ _26317_/CLK _26317_/D vssd1 vssd1 vccd1 vccd1 _26317_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_107_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23529_ _23526_/Y _23528_/Y _24858_/S vssd1 vssd1 vccd1 vccd1 _23529_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_80_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14262_ _18956_/B _14262_/B vssd1 vssd1 vccd1 vccd1 _14262_/Y sky130_fd_sc_hd__nor2_1
X_17050_ _25585_/Q vssd1 vssd1 vccd1 vccd1 _19138_/B sky130_fd_sc_hd__inv_2
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26248_ _26248_/CLK _26248_/D vssd1 vssd1 vccd1 vccd1 _26248_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_123_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16001_ _16054_/C _16054_/B vssd1 vssd1 vccd1 vccd1 _16001_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_33_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13213_ _13207_/X _13211_/X _13192_/X _13212_/X vssd1 vssd1 vccd1 vccd1 _13213_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14193_ hold423/X _14192_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold424/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26179_ _26181_/CLK _26179_/D vssd1 vssd1 vccd1 vccd1 _26179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13144_ hold990/X _13320_/B vssd1 vssd1 vccd1 vccd1 _13144_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17952_ _25858_/Q _21763_/A vssd1 vssd1 vccd1 vccd1 _17960_/A sky130_fd_sc_hd__or2_2
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13075_ _17646_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13075_/X sky130_fd_sc_hd__or2_1
X_16903_ _16904_/B _16904_/A vssd1 vssd1 vccd1 vccd1 _16903_/X sky130_fd_sc_hd__or2_1
X_17883_ _17883_/A _19114_/A vssd1 vssd1 vccd1 vccd1 _17884_/A sky130_fd_sc_hd__xor2_2
X_19622_ _19620_/X _19621_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19622_/Y sky130_fd_sc_hd__a21oi_1
X_16834_ _16858_/A _16834_/B vssd1 vssd1 vccd1 vccd1 _16834_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19553_ _19545_/X _19552_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19553_/Y sky130_fd_sc_hd__o21ai_1
X_16765_ _16763_/Y _16764_/Y _16594_/X vssd1 vssd1 vccd1 vccd1 _16765_/Y sky130_fd_sc_hd__a21oi_1
X_13977_ _26294_/Q _13801_/X _13793_/X _13976_/Y vssd1 vssd1 vccd1 vccd1 _13978_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18504_ _25879_/Q _22148_/A vssd1 vssd1 vccd1 vccd1 _18512_/A sky130_fd_sc_hd__or2_2
X_15716_ _15716_/A _15718_/B vssd1 vssd1 vccd1 vccd1 _15716_/Y sky130_fd_sc_hd__nand2_1
X_12928_ _17442_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12928_/X sky130_fd_sc_hd__or2_1
X_19484_ _26239_/Q _19483_/X hold841/X vssd1 vssd1 vccd1 vccd1 _19484_/Y sky130_fd_sc_hd__a21oi_1
X_16696_ _16696_/A _16696_/B vssd1 vssd1 vccd1 vccd1 _16697_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_158_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18435_ _18535_/A _18435_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18435_/X sky130_fd_sc_hd__and3_1
X_15647_ _15647_/A vssd1 vssd1 vccd1 vccd1 _23047_/B sky130_fd_sc_hd__inv_2
XFILLER_0_69_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _17309_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12859_/X sky130_fd_sc_hd__or2_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18366_ _18951_/A _25744_/Q vssd1 vssd1 vccd1 vccd1 _18368_/A sky130_fd_sc_hd__nand2_1
X_15578_ _15547_/A _15577_/A _15572_/A vssd1 vssd1 vccd1 vccd1 _15578_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_150_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17317_ _25645_/Q vssd1 vssd1 vccd1 vccd1 _20088_/B sky130_fd_sc_hd__inv_2
XFILLER_0_126_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14529_ _14529_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14529_/Y sky130_fd_sc_hd__nand2_1
X_18297_ _18295_/Y _18296_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25659_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17248_ _25606_/Q vssd1 vssd1 vccd1 vccd1 _20909_/B sky130_fd_sc_hd__inv_2
XFILLER_0_113_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17179_ _25601_/Q vssd1 vssd1 vccd1 vccd1 _20741_/B sky130_fd_sc_hd__inv_2
XFILLER_0_24_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20190_ _26281_/Q _20078_/X hold557/X vssd1 vssd1 vccd1 vccd1 _20194_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2404 _26177_/Q vssd1 vssd1 vccd1 vccd1 hold2404/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2415 _15295_/Y vssd1 vssd1 vccd1 vccd1 _25445_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2426 _24011_/X vssd1 vssd1 vccd1 vccd1 _24012_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2437 _26068_/Q vssd1 vssd1 vccd1 vccd1 hold2437/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2448 _25665_/Q vssd1 vssd1 vccd1 vccd1 _13188_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1703 _25835_/Q vssd1 vssd1 vccd1 vccd1 _21687_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2459 _25454_/Q vssd1 vssd1 vccd1 vccd1 _15439_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1714 _17033_/Y vssd1 vssd1 vccd1 vccd1 _25583_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1725 _25861_/Q vssd1 vssd1 vccd1 vccd1 _22432_/B sky130_fd_sc_hd__dlygate4sd3_1
X_22900_ _22900_/A _22900_/B vssd1 vssd1 vccd1 vccd1 _22901_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23880_ hold2075/X _26031_/Q _23907_/S vssd1 vssd1 vccd1 vccd1 _23880_/X sky130_fd_sc_hd__mux2_1
Xhold1736 _25786_/Q vssd1 vssd1 vccd1 vccd1 _20504_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1747 _25597_/Q vssd1 vssd1 vccd1 vccd1 _17230_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1758 _25654_/Q vssd1 vssd1 vccd1 vccd1 _18181_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1769 _25873_/Q vssd1 vssd1 vccd1 vccd1 _22740_/B sky130_fd_sc_hd__buf_1
X_22831_ _26062_/Q vssd1 vssd1 vccd1 vccd1 _22832_/A sky130_fd_sc_hd__inv_2
XFILLER_0_17_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25550_ _25877_/CLK _25550_/D vssd1 vssd1 vccd1 vccd1 _25550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22762_ _22762_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22762_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21713_ _26340_/Q _19130_/X hold425/X vssd1 vssd1 vccd1 vccd1 _21716_/B sky130_fd_sc_hd__a21oi_1
X_24501_ hold2559/X _26231_/Q _24510_/S vssd1 vssd1 vccd1 vccd1 _24501_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_177_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25481_ _25483_/CLK hold859/X vssd1 vssd1 vccd1 vccd1 hold858/A sky130_fd_sc_hd__dfxtp_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22693_ _18938_/A _25836_/Q _22691_/Y _22692_/Y vssd1 vssd1 vccd1 vccd1 _22694_/B
+ sky130_fd_sc_hd__a31o_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24432_ _24432_/A vssd1 vssd1 vccd1 vccd1 _26208_/D sky130_fd_sc_hd__clkbuf_1
X_21644_ _21692_/B _21644_/B vssd1 vssd1 vccd1 vccd1 _21646_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24363_ hold2322/X hold2241/X _24433_/S vssd1 vssd1 vccd1 vccd1 _24364_/A sky130_fd_sc_hd__mux2_1
XANTENNA_40 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21575_ _21578_/A _21629_/B vssd1 vssd1 vccd1 vccd1 _21577_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_151_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_51 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23314_ _23314_/A hold896/X vssd1 vssd1 vccd1 vccd1 hold897/A sky130_fd_sc_hd__nand2_1
XFILLER_0_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26102_ _26103_/CLK _26102_/D vssd1 vssd1 vccd1 vccd1 _26102_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_62 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20526_ _20526_/A _20526_/B _20526_/C vssd1 vssd1 vccd1 vccd1 _20527_/B sky130_fd_sc_hd__nand3_1
XANTENNA_73 _17549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_24294_ _24294_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24295_/A sky130_fd_sc_hd__and2_1
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23245_ _23245_/A _23245_/B _23249_/A vssd1 vssd1 vccd1 vccd1 _23246_/A sky130_fd_sc_hd__or3_1
XFILLER_0_160_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26033_ _26041_/CLK _26033_/D vssd1 vssd1 vccd1 vccd1 _26033_/Q sky130_fd_sc_hd__dfxtp_1
X_20457_ _20457_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20462_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23176_ _23175_/A _22999_/C _23175_/B vssd1 vssd1 vccd1 vccd1 _23177_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20388_ _20386_/Y _20387_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _20388_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22127_ _22807_/B vssd1 vssd1 vccd1 vccd1 _22808_/A sky130_fd_sc_hd__inv_2
XFILLER_0_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22058_ _22058_/A _22058_/B vssd1 vssd1 vccd1 vccd1 _22058_/Y sky130_fd_sc_hd__nand2_1
X_13900_ _14000_/A hold611/X vssd1 vssd1 vccd1 vccd1 hold612/A sky130_fd_sc_hd__nand2_1
X_21009_ _21483_/B _21529_/C vssd1 vssd1 vccd1 vccd1 _21010_/C sky130_fd_sc_hd__nand2_1
X_14880_ _25858_/Q _13466_/A _14879_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14881_/A
+ sky130_fd_sc_hd__a22o_1
X_25817_ _25817_/CLK _25817_/D vssd1 vssd1 vccd1 vccd1 _25817_/Q sky130_fd_sc_hd__dfxtp_2
X_13831_ hold660/X _13830_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold661/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16550_ _16550_/A vssd1 vssd1 vccd1 vccd1 _16564_/B sky130_fd_sc_hd__inv_2
XFILLER_0_98_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25748_ _25748_/CLK _25748_/D vssd1 vssd1 vccd1 vccd1 _25748_/Q sky130_fd_sc_hd__dfxtp_1
X_13762_ _14120_/A vssd1 vssd1 vccd1 vccd1 _13876_/B sky130_fd_sc_hd__buf_6
XFILLER_0_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15501_ hold2672/X _15500_/Y _15464_/X vssd1 vssd1 vccd1 vccd1 _15501_/Y sky130_fd_sc_hd__a21oi_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12713_ _12713_/A _12713_/B _12713_/C _12713_/D vssd1 vssd1 vccd1 vccd1 _12714_/B
+ sky130_fd_sc_hd__or4_1
X_16481_ _16485_/A _16481_/B vssd1 vssd1 vccd1 vccd1 _16482_/A sky130_fd_sc_hd__xor2_1
X_25679_ _26313_/CLK _25679_/D vssd1 vssd1 vccd1 vccd1 _25679_/Q sky130_fd_sc_hd__dfxtp_1
X_13693_ _13760_/A hold665/X vssd1 vssd1 vccd1 vccd1 hold666/A sky130_fd_sc_hd__nand2_1
XFILLER_0_127_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18220_ _18446_/A _25737_/Q _18952_/C vssd1 vssd1 vccd1 vccd1 _18221_/C sky130_fd_sc_hd__nand3_1
X_15432_ _16837_/B vssd1 vssd1 vccd1 vccd1 _22848_/B sky130_fd_sc_hd__inv_2
X_12644_ _12644_/A _12644_/B _12644_/C vssd1 vssd1 vccd1 vccd1 _12645_/D sky130_fd_sc_hd__or3_1
XFILLER_0_183_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18151_ _25846_/Q _18151_/B _18150_/Y vssd1 vssd1 vccd1 vccd1 _18161_/A sky130_fd_sc_hd__or3b_2
XFILLER_0_65_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15363_ _15363_/A vssd1 vssd1 vccd1 vccd1 _15373_/B sky130_fd_sc_hd__inv_2
X_12575_ _12575_/A _12575_/B vssd1 vssd1 vccd1 vccd1 _12582_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17102_ _20507_/B _25851_/Q _25787_/Q vssd1 vssd1 vccd1 vccd1 _17103_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_108_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14314_ _14344_/A hold257/X vssd1 vssd1 vccd1 vccd1 hold258/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18082_ _18611_/A _18086_/B vssd1 vssd1 vccd1 vccd1 _18084_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15294_ _15294_/A _15307_/A vssd1 vssd1 vccd1 vccd1 _15294_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_123_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17033_ _17031_/Y _17032_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _17033_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14245_ _26337_/Q _13518_/B _14170_/X _14244_/Y vssd1 vssd1 vccd1 vccd1 _14246_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14176_ _14236_/A hold698/X vssd1 vssd1 vccd1 vccd1 hold699/A sky130_fd_sc_hd__nand2_1
XFILLER_0_22_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13127_ _26157_/Q _13065_/X _13126_/X vssd1 vssd1 vccd1 vccd1 _13127_/X sky130_fd_sc_hd__a21o_1
X_18984_ _18982_/X _18879_/X _18983_/X vssd1 vssd1 vccd1 vccd1 _18985_/A sky130_fd_sc_hd__a21o_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17935_ _19216_/A vssd1 vssd1 vccd1 vccd1 _22160_/B sky130_fd_sc_hd__inv_2
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _17624_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13058_/X sky130_fd_sc_hd__or2_1
XFILLER_0_178_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17866_ _17866_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _17866_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_178_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16817_ _16817_/A _16817_/B vssd1 vssd1 vccd1 vccd1 _16817_/Y sky130_fd_sc_hd__nand2_1
X_19605_ _19621_/B _19692_/B vssd1 vssd1 vccd1 vccd1 _19607_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17797_ _18098_/A vssd1 vssd1 vccd1 vccd1 _18528_/A sky130_fd_sc_hd__buf_12
XFILLER_0_178_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19536_ _19537_/B _19537_/A vssd1 vssd1 vccd1 vccd1 _19536_/X sky130_fd_sc_hd__or2_1
XFILLER_0_88_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16748_ _16746_/X _16711_/X _16747_/Y _25867_/Q _14170_/X vssd1 vssd1 vccd1 vccd1
+ _16749_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_177_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19467_ _19723_/A _19467_/B vssd1 vssd1 vccd1 vccd1 _19467_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16679_ _16695_/B _16679_/B vssd1 vssd1 vccd1 vccd1 _16685_/B sky130_fd_sc_hd__and2_1
XFILLER_0_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18418_ _18641_/A _19303_/A vssd1 vssd1 vccd1 vccd1 _18418_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_146_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19398_ _26233_/Q _12537_/B hold455/X vssd1 vssd1 vccd1 vccd1 _19398_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18349_ _21164_/C _21915_/A vssd1 vssd1 vccd1 vccd1 _21156_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_173_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21360_ _21636_/A _21360_/B _21359_/X vssd1 vssd1 vccd1 vccd1 _21361_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_185_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20311_ _20314_/A _20314_/C vssd1 vssd1 vccd1 vccd1 _20312_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold800 hold800/A vssd1 vssd1 vccd1 vccd1 hold800/X sky130_fd_sc_hd__dlygate4sd3_1
X_21291_ _21291_/A _21291_/B vssd1 vssd1 vccd1 vccd1 _21294_/B sky130_fd_sc_hd__nand2_1
Xhold811 hold811/A vssd1 vssd1 vccd1 vccd1 hold811/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23030_ _26074_/Q vssd1 vssd1 vccd1 vccd1 _23031_/A sky130_fd_sc_hd__inv_2
Xhold822 hold822/A vssd1 vssd1 vccd1 vccd1 hold822/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 hold833/A vssd1 vssd1 vccd1 vccd1 hold833/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20242_ _20244_/B vssd1 vssd1 vccd1 vccd1 _20243_/B sky130_fd_sc_hd__inv_2
Xhold844 hold844/A vssd1 vssd1 vccd1 vccd1 hold844/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 hold855/A vssd1 vssd1 vccd1 vccd1 hold855/X sky130_fd_sc_hd__buf_1
Xhold866 hold866/A vssd1 vssd1 vccd1 vccd1 hold866/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold877 hold877/A vssd1 vssd1 vccd1 vccd1 hold877/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 hold888/A vssd1 vssd1 vccd1 vccd1 hold888/X sky130_fd_sc_hd__dlygate4sd3_1
X_20173_ _21434_/A vssd1 vssd1 vccd1 vccd1 _21433_/A sky130_fd_sc_hd__inv_2
Xhold899 hold899/A vssd1 vssd1 vccd1 vccd1 hold899/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_0_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2201 _26155_/Q vssd1 vssd1 vccd1 vccd1 hold2201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2212 _26000_/Q vssd1 vssd1 vccd1 vccd1 _14866_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2223 _24418_/X vssd1 vssd1 vccd1 vccd1 _24419_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24981_ _24983_/CLK _24981_/D vssd1 vssd1 vccd1 vccd1 _24981_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2234 _26138_/Q vssd1 vssd1 vccd1 vccd1 hold2234/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1500 _23118_/Y vssd1 vssd1 vccd1 vccd1 _25896_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2245 _26149_/Q vssd1 vssd1 vccd1 vccd1 hold2245/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2256 _26004_/Q vssd1 vssd1 vccd1 vccd1 hold2256/X sky130_fd_sc_hd__buf_1
Xhold1511 _25775_/Q vssd1 vssd1 vccd1 vccd1 _20085_/B sky130_fd_sc_hd__buf_1
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23932_ hold2456/X hold2126/X _24001_/S vssd1 vssd1 vccd1 vccd1 _23933_/A sky130_fd_sc_hd__mux2_1
Xhold2267 _26098_/Q vssd1 vssd1 vccd1 vccd1 hold2267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 _17446_/Y vssd1 vssd1 vccd1 vccd1 _25616_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1533 _25116_/Q vssd1 vssd1 vccd1 vccd1 _18990_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2278 _25702_/Q vssd1 vssd1 vccd1 vccd1 _13420_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1544 _21236_/Y vssd1 vssd1 vccd1 vccd1 _25809_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2289 _15046_/Y vssd1 vssd1 vccd1 vccd1 hold2289/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1555 _25823_/Q vssd1 vssd1 vccd1 vccd1 _21492_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1566 _25816_/Q vssd1 vssd1 vccd1 vccd1 _21380_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23863_ _23863_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23864_/A sky130_fd_sc_hd__and2_1
Xhold1577 _23150_/Y vssd1 vssd1 vccd1 vccd1 _25898_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1588 _25822_/Q vssd1 vssd1 vccd1 vccd1 _21476_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1599 _17049_/Y vssd1 vssd1 vccd1 vccd1 _25584_/D sky130_fd_sc_hd__dlygate4sd3_1
X_25602_ _25604_/CLK _25602_/D vssd1 vssd1 vccd1 vccd1 _25602_/Q sky130_fd_sc_hd__dfxtp_2
X_22814_ _26061_/Q vssd1 vssd1 vccd1 vccd1 _22815_/A sky130_fd_sc_hd__inv_2
X_23794_ _14884_/B _14893_/B _23831_/S vssd1 vssd1 vccd1 vccd1 _23795_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_79_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25533_ _25533_/CLK hold888/X vssd1 vssd1 vccd1 vccd1 hold887/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22745_ _22745_/A _22745_/B vssd1 vssd1 vccd1 vccd1 _22746_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_181_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xascon_wrapper_13 vssd1 vssd1 vccd1 vccd1 ascon_wrapper_13/HI io_oeb[10] sky130_fd_sc_hd__conb_1
XFILLER_0_109_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25464_ _25532_/CLK hold947/X vssd1 vssd1 vccd1 vccd1 hold946/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22676_ _22676_/A _22676_/B vssd1 vssd1 vccd1 vccd1 _22677_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_164_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24415_ hold1989/X _26203_/Q _24433_/S vssd1 vssd1 vccd1 vccd1 _24415_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21627_ _21627_/A _21627_/B _21627_/C vssd1 vssd1 vccd1 vccd1 _21631_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_35_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25395_ _26208_/CLK _25395_/D vssd1 vssd1 vccd1 vccd1 _25395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21558_ _21556_/Y _21557_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21558_/Y sky130_fd_sc_hd__a21oi_1
X_24346_ _24346_/A vssd1 vssd1 vccd1 vccd1 _26180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20509_ _20509_/A _25851_/Q vssd1 vssd1 vccd1 vccd1 _20514_/B sky130_fd_sc_hd__nand2_1
X_24277_ _24277_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24278_/A sky130_fd_sc_hd__and2_1
XFILLER_0_106_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21489_ _21636_/A _21489_/B _21488_/X vssd1 vssd1 vccd1 vccd1 _21490_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_160_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14030_ _14061_/A _14030_/B vssd1 vssd1 vccd1 vccd1 _14030_/Y sky130_fd_sc_hd__nand2_1
X_23228_ _23231_/A _24836_/B _23228_/C vssd1 vssd1 vccd1 vccd1 _23229_/A sky130_fd_sc_hd__and3_1
X_26016_ _26021_/CLK _26016_/D vssd1 vssd1 vccd1 vccd1 _26016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23159_ _23159_/A _23159_/B _23191_/C vssd1 vssd1 vccd1 vccd1 _23161_/A sky130_fd_sc_hd__or3_1
XFILLER_0_30_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15981_ _15979_/Y hold810/X _15805_/X vssd1 vssd1 vccd1 vccd1 hold811/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17720_ _17725_/A _17764_/B _17725_/C vssd1 vssd1 vccd1 vccd1 _17724_/B sky130_fd_sc_hd__nand3_1
X_14932_ _14932_/A _14932_/B vssd1 vssd1 vccd1 vccd1 _14947_/A sky130_fd_sc_hd__nand2_1
X_17651_ _17651_/A _17651_/B vssd1 vssd1 vccd1 vccd1 _17652_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14863_ _25856_/Q _14170_/A _15049_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14864_/B
+ sky130_fd_sc_hd__a22o_1
X_16602_ _16602_/A _16602_/B vssd1 vssd1 vccd1 vccd1 _16650_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_159_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13814_ _25765_/Q vssd1 vssd1 vccd1 vccd1 _18793_/B sky130_fd_sc_hd__inv_2
X_17582_ _17582_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17582_/Y sky130_fd_sc_hd__nand2_1
X_14794_ _14794_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14794_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_98_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19321_ _19322_/B _19322_/A vssd1 vssd1 vccd1 vccd1 _19321_/X sky130_fd_sc_hd__or2_1
XFILLER_0_187_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16533_ _16539_/B _16534_/A vssd1 vssd1 vccd1 vccd1 _16533_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_58_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13745_ _26257_/Q _13612_/X _13605_/X _13744_/Y vssd1 vssd1 vccd1 vccd1 _13746_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19252_ _19252_/A _19994_/B _19252_/C vssd1 vssd1 vccd1 vccd1 _19252_/X sky130_fd_sc_hd__and3_1
X_16464_ _16676_/A _16464_/B vssd1 vssd1 vccd1 vccd1 _16466_/A sky130_fd_sc_hd__or2_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13676_ _18347_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13676_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_155_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18203_ _18203_/A _18203_/B _18203_/C vssd1 vssd1 vccd1 vccd1 _21974_/A sky130_fd_sc_hd__nand3_2
X_15415_ _15413_/X _15414_/Y _15090_/X vssd1 vssd1 vccd1 vccd1 _25452_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12627_ _12629_/B vssd1 vssd1 vccd1 vccd1 _12645_/A sky130_fd_sc_hd__inv_2
X_19183_ _19183_/A _19983_/B vssd1 vssd1 vccd1 vccd1 _19183_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_66_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16395_ _16404_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16395_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_5_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18134_ _18445_/A _18138_/B vssd1 vssd1 vccd1 vccd1 _18136_/A sky130_fd_sc_hd__nand2_1
X_15346_ _15344_/Y _15345_/Y _15090_/X vssd1 vssd1 vccd1 vccd1 hold976/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12558_ hold4/X _12558_/B vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__nor2_1
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18065_ _21958_/A _25588_/Q vssd1 vssd1 vccd1 vccd1 _18067_/B sky130_fd_sc_hd__nand2_1
X_15277_ _15277_/A _15277_/B vssd1 vssd1 vccd1 vccd1 _15827_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_124_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12489_ input7/X vssd1 vssd1 vccd1 vccd1 _24745_/A sky130_fd_sc_hd__inv_6
XFILLER_0_124_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold107 hold107/A vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold118 hold118/A vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 hold129/A vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__dlygate4sd3_1
X_17016_ _17272_/A _17016_/B vssd1 vssd1 vccd1 vccd1 _17016_/Y sky130_fd_sc_hd__nand2_1
X_14228_ _14264_/A _14228_/B vssd1 vssd1 vccd1 vccd1 _14228_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ _18613_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14159_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18967_ _19018_/A _18967_/B vssd1 vssd1 vccd1 vccd1 _18967_/X sky130_fd_sc_hd__xor2_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17918_ _17916_/Y _17917_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _17918_/Y sky130_fd_sc_hd__a21oi_1
X_18898_ _19010_/A _19059_/B vssd1 vssd1 vccd1 vccd1 _18899_/B sky130_fd_sc_hd__xnor2_1
X_17849_ _17849_/A _20701_/A vssd1 vssd1 vccd1 vccd1 _18392_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_179_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20860_ _20860_/A _21840_/B _20860_/C vssd1 vssd1 vccd1 vccd1 _20863_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_178_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19519_ _21183_/A _21947_/B _25616_/Q vssd1 vssd1 vccd1 vccd1 _21187_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_92_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20791_ _20791_/A _20791_/B vssd1 vssd1 vccd1 vccd1 _20795_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22530_ _22529_/A _22454_/X _22529_/B vssd1 vssd1 vccd1 vccd1 _22531_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22461_ _22459_/X _22460_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22461_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24200_ hold2110/X hold1930/X _24203_/S vssd1 vssd1 vccd1 vccd1 _24201_/A sky130_fd_sc_hd__mux2_1
X_21412_ _21573_/A _21412_/B vssd1 vssd1 vccd1 vccd1 _21412_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_146_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25180_ _25773_/CLK hold848/X vssd1 vssd1 vccd1 vccd1 hold847/A sky130_fd_sc_hd__dfxtp_1
X_22392_ _18696_/A _25824_/Q _22390_/Y _22391_/Y vssd1 vssd1 vccd1 vccd1 _22393_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24131_ _24131_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24132_/A sky130_fd_sc_hd__and2_1
XFILLER_0_142_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21343_ _21342_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21343_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_103_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24062_ hold2096/X _26088_/Q _24126_/S vssd1 vssd1 vccd1 vccd1 _24062_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold630 hold630/A vssd1 vssd1 vccd1 vccd1 hold630/X sky130_fd_sc_hd__dlygate4sd3_1
X_21274_ _21691_/C vssd1 vssd1 vccd1 vccd1 _21694_/B sky130_fd_sc_hd__inv_2
XFILLER_0_25_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold641 hold641/A vssd1 vssd1 vccd1 vccd1 hold641/X sky130_fd_sc_hd__dlygate4sd3_1
X_23013_ _15619_/B _22893_/A _22829_/X vssd1 vssd1 vccd1 vccd1 _23013_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold652 hold652/A vssd1 vssd1 vccd1 vccd1 hold652/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold663 hold663/A vssd1 vssd1 vccd1 vccd1 hold663/X sky130_fd_sc_hd__dlygate4sd3_1
X_20225_ _20225_/A _20225_/B vssd1 vssd1 vccd1 vccd1 _20226_/A sky130_fd_sc_hd__nand2_1
Xhold674 hold674/A vssd1 vssd1 vccd1 vccd1 hold674/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 hold685/A vssd1 vssd1 vccd1 vccd1 hold685/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 hold696/A vssd1 vssd1 vccd1 vccd1 hold696/X sky130_fd_sc_hd__dlygate4sd3_1
X_20156_ _20155_/Y _21228_/A _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20156_/X
+ sky130_fd_sc_hd__a211o_1
Xhold2020 _25930_/Q vssd1 vssd1 vccd1 vccd1 _23336_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2031 _23377_/X vssd1 vssd1 vccd1 vccd1 _23378_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2042 _15362_/Y vssd1 vssd1 vccd1 vccd1 _25449_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2053 _26065_/Q vssd1 vssd1 vccd1 vccd1 hold2053/X sky130_fd_sc_hd__dlygate4sd3_1
X_24964_ _25418_/CLK hold5/X vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfxtp_1
X_20087_ _20087_/A _22718_/B vssd1 vssd1 vccd1 vccd1 _20088_/A sky130_fd_sc_hd__nand2_1
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2064 _14933_/Y vssd1 vssd1 vccd1 vccd1 _14948_/A sky130_fd_sc_hd__buf_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1330 _14901_/Y vssd1 vssd1 vccd1 vccd1 _25411_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2075 _26030_/Q vssd1 vssd1 vccd1 vccd1 hold2075/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2086 _25954_/Q vssd1 vssd1 vccd1 vccd1 hold2086/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1341 _25571_/Q vssd1 vssd1 vccd1 vccd1 _15647_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23915_ _23915_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23916_/A sky130_fd_sc_hd__and2_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2097 _24062_/X vssd1 vssd1 vccd1 vccd1 _24063_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1352 _19453_/Y vssd1 vssd1 vccd1 vccd1 _25733_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1363 _25772_/Q vssd1 vssd1 vccd1 vccd1 _19987_/B sky130_fd_sc_hd__dlygate4sd3_1
X_24895_ _24893_/X _24894_/X _24957_/S vssd1 vssd1 vccd1 vccd1 _24895_/X sky130_fd_sc_hd__mux2_1
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1374 _14751_/Y vssd1 vssd1 vccd1 vccd1 _25394_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1385 _25723_/Q vssd1 vssd1 vccd1 vccd1 _19311_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1396 _19954_/Y vssd1 vssd1 vccd1 vccd1 _25769_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23846_ _23846_/A vssd1 vssd1 vccd1 vccd1 _26019_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23777_ _23777_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23778_/A sky130_fd_sc_hd__and2_1
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20989_ _20989_/A _20989_/B vssd1 vssd1 vccd1 vccd1 _20990_/A sky130_fd_sc_hd__nand2_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25516_ _25537_/CLK hold520/X vssd1 vssd1 vccd1 vccd1 hold518/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13530_ _13642_/A hold509/X vssd1 vssd1 vccd1 vccd1 hold510/A sky130_fd_sc_hd__nand2_1
X_22728_ _22728_/A _22728_/B vssd1 vssd1 vccd1 vccd1 _22729_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25447_ _25511_/CLK _25447_/D vssd1 vssd1 vccd1 vccd1 _25447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13461_ _19082_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13461_/X sky130_fd_sc_hd__or2_1
X_22659_ _16771_/B _22421_/X _22653_/X _22654_/Y _22658_/X vssd1 vssd1 vccd1 vccd1
+ _22660_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15200_ _15188_/X _15268_/B _16698_/A vssd1 vssd1 vccd1 vccd1 _15200_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16180_ _16180_/A _16180_/B vssd1 vssd1 vccd1 vccd1 _16181_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_129_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25378_ _25378_/CLK hold43/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dfxtp_1
X_13392_ _26200_/Q _13239_/X _13391_/X vssd1 vssd1 vccd1 vccd1 _13392_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15131_ _15956_/A hold931/X vssd1 vssd1 vccd1 vccd1 _15131_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24329_ hold2400/X hold1891/X _24356_/S vssd1 vssd1 vccd1 vccd1 _24330_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_62_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15062_ _15062_/A _15067_/B vssd1 vssd1 vccd1 vccd1 _15062_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14013_ hold579/X _14012_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold580/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19870_ _19870_/A _19980_/B _19870_/C vssd1 vssd1 vccd1 vccd1 _19870_/X sky130_fd_sc_hd__and3_1
X_18821_ _18821_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18821_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_156_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18752_ _18954_/A _25763_/Q vssd1 vssd1 vccd1 vccd1 _18754_/A sky130_fd_sc_hd__nand2_1
X_15964_ _15962_/X _15963_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _15964_/X sky130_fd_sc_hd__a21o_1
X_17703_ _17703_/A _17704_/A vssd1 vssd1 vccd1 vccd1 _17709_/A sky130_fd_sc_hd__nand2_1
X_14915_ _14915_/A vssd1 vssd1 vccd1 vccd1 _14919_/B sky130_fd_sc_hd__inv_2
XFILLER_0_76_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18683_ _18681_/Y _18682_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25678_/D sky130_fd_sc_hd__a21oi_1
X_15895_ _15895_/A _15895_/B vssd1 vssd1 vccd1 vccd1 _15942_/B sky130_fd_sc_hd__and2_1
XFILLER_0_37_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17634_ _17634_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _17634_/Y sky130_fd_sc_hd__nand2_1
X_14846_ _14846_/A vssd1 vssd1 vccd1 vccd1 _15027_/A sky130_fd_sc_hd__inv_2
XFILLER_0_77_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17565_ _17563_/X _17528_/X _17564_/X vssd1 vssd1 vccd1 vccd1 _17566_/A sky130_fd_sc_hd__a21o_1
X_14777_ _14900_/A _14777_/B vssd1 vssd1 vccd1 vccd1 _14777_/Y sky130_fd_sc_hd__nand2_1
X_19304_ _20740_/A _21729_/B _25601_/Q vssd1 vssd1 vccd1 vccd1 _20745_/C sky130_fd_sc_hd__nand3_1
X_16516_ _16514_/X _16515_/Y _16231_/A vssd1 vssd1 vccd1 vccd1 _16516_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_129_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13728_ _13823_/A _13728_/B vssd1 vssd1 vccd1 vccd1 _13728_/Y sky130_fd_sc_hd__nand2_1
X_17496_ _17605_/A _17496_/B vssd1 vssd1 vccd1 vccd1 _17496_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19235_ _26221_/Q hold843/X vssd1 vssd1 vccd1 vccd1 _19235_/Y sky130_fd_sc_hd__nand2_1
X_16447_ _16447_/A _16686_/B _16447_/C vssd1 vssd1 vccd1 vccd1 _16447_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13659_ _26243_/Q _13612_/X _13605_/X _13658_/Y vssd1 vssd1 vccd1 vccd1 _13660_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19166_ _19972_/B _19167_/A vssd1 vssd1 vccd1 vccd1 _19166_/X sky130_fd_sc_hd__or2_1
X_16378_ _16378_/A _16378_/B vssd1 vssd1 vccd1 vccd1 _16379_/A sky130_fd_sc_hd__and2_1
XFILLER_0_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18117_ _25845_/Q _18117_/B _18117_/C vssd1 vssd1 vccd1 vccd1 _18127_/A sky130_fd_sc_hd__nor3_2
X_15329_ _15321_/B _15306_/A _15321_/A vssd1 vssd1 vccd1 vccd1 _15329_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_42_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19097_ _25652_/Q _20248_/B vssd1 vssd1 vccd1 vccd1 _19097_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_170_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18048_ _18098_/A vssd1 vssd1 vccd1 vccd1 _18792_/A sky130_fd_sc_hd__buf_12
XFILLER_0_111_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20010_ _20010_/A _22095_/B vssd1 vssd1 vccd1 vccd1 _20011_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19999_ _19999_/A _22665_/B vssd1 vssd1 vccd1 vccd1 _20000_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_158_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21961_ _21962_/A _21962_/B _22994_/A vssd1 vssd1 vccd1 vccd1 _21961_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23700_ _23700_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23701_/A sky130_fd_sc_hd__and2_1
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20912_ _25862_/Q vssd1 vssd1 vccd1 vccd1 _21909_/B sky130_fd_sc_hd__inv_2
X_21892_ _21893_/A _21893_/B _22960_/A vssd1 vssd1 vccd1 vccd1 _21892_/X sky130_fd_sc_hd__a21o_1
X_24680_ hold2675/X hold2495/X _24740_/S vssd1 vssd1 vccd1 vccd1 _24681_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23631_ hold1947/X hold1926/X _23677_/S vssd1 vssd1 vccd1 vccd1 _23633_/A sky130_fd_sc_hd__mux2_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20843_ _21435_/B _21709_/B vssd1 vssd1 vccd1 vccd1 _20844_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_178_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23562_ _24922_/S hold167/A _23561_/X vssd1 vssd1 vccd1 vccd1 _23562_/Y sky130_fd_sc_hd__o21ai_1
X_20774_ _21042_/A _20774_/B _20773_/X vssd1 vssd1 vccd1 vccd1 _20775_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_92_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25301_ _26136_/CLK hold139/X vssd1 vssd1 vccd1 vccd1 hold137/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22513_ _25829_/Q _22513_/B vssd1 vssd1 vccd1 vccd1 _22513_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23493_ hold125/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23493_/X sky130_fd_sc_hd__or2b_1
X_26281_ _26281_/CLK _26281_/D vssd1 vssd1 vccd1 vccd1 _26281_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_162_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_170_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _25729_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_107_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22444_ _23007_/A _22858_/B vssd1 vssd1 vccd1 vccd1 _22446_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25232_ _25687_/CLK hold529/X vssd1 vssd1 vccd1 vccd1 hold527/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22375_ _22375_/A _22375_/B vssd1 vssd1 vccd1 vccd1 _22376_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25163_ _25743_/CLK hold547/X vssd1 vssd1 vccd1 vccd1 hold545/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24114_ hold2382/X _26105_/Q _24126_/S vssd1 vssd1 vccd1 vccd1 _24114_/X sky130_fd_sc_hd__mux2_1
X_21326_ _26316_/Q hold587/A vssd1 vssd1 vccd1 vccd1 _21326_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25094_ _26308_/CLK _25094_/D vssd1 vssd1 vccd1 vccd1 _25094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24045_ _24045_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24046_/A sky130_fd_sc_hd__and2_1
Xhold460 hold460/A vssd1 vssd1 vccd1 vccd1 hold460/X sky130_fd_sc_hd__dlygate4sd3_1
X_21257_ _21256_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21257_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_102_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold471 hold471/A vssd1 vssd1 vccd1 vccd1 hold471/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 hold482/A vssd1 vssd1 vccd1 vccd1 hold482/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 hold493/A vssd1 vssd1 vccd1 vccd1 hold493/X sky130_fd_sc_hd__dlygate4sd3_1
X_20208_ _20208_/A _20208_/B _20208_/C vssd1 vssd1 vccd1 vccd1 _20209_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_159_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21188_ _21190_/B _21190_/C vssd1 vssd1 vccd1 vccd1 _21189_/A sky130_fd_sc_hd__nand2_1
X_20139_ _20139_/A _20139_/B _20139_/C vssd1 vssd1 vccd1 vccd1 _20148_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_95_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25996_ _25998_/CLK _25996_/D vssd1 vssd1 vccd1 vccd1 _25996_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24947_ _24946_/A _24944_/X _24958_/B _24946_/Y vssd1 vssd1 vccd1 vccd1 _24947_/X
+ sky130_fd_sc_hd__a211o_1
X_12961_ _26254_/Q _25623_/Q vssd1 vssd1 vccd1 vccd1 _14419_/A sky130_fd_sc_hd__xor2_2
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1160 _12885_/X vssd1 vssd1 vccd1 vccd1 _25028_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _14899_/B vssd1 vssd1 vccd1 vccd1 _14864_/A sky130_fd_sc_hd__clkbuf_8
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1171 _25059_/Q vssd1 vssd1 vccd1 vccd1 _17609_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1182 _12991_/X vssd1 vssd1 vccd1 vccd1 _25048_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15680_ _15680_/A vssd1 vssd1 vccd1 vccd1 _15690_/B sky130_fd_sc_hd__inv_2
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24878_ _15971_/B _15985_/B _24942_/S vssd1 vssd1 vccd1 vccd1 _24879_/A sky130_fd_sc_hd__mux2_1
X_12892_ _26241_/Q _25610_/Q vssd1 vssd1 vccd1 vccd1 _14376_/A sky130_fd_sc_hd__xor2_1
Xhold1193 _25805_/Q vssd1 vssd1 vccd1 vccd1 _21844_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _14629_/Y hold261/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold262/A sky130_fd_sc_hd__a21oi_1
X_23829_ _23829_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23830_/A sky130_fd_sc_hd__and2_1
XFILLER_0_135_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17350_ _19488_/A _17350_/B vssd1 vssd1 vccd1 vccd1 _17594_/A sky130_fd_sc_hd__xor2_4
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _14560_/Y hold213/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold214/A sky130_fd_sc_hd__a21oi_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _16473_/A hold863/X vssd1 vssd1 vccd1 vccd1 _16301_/Y sky130_fd_sc_hd__nand2_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _26220_/Q _13426_/X _13468_/X _13512_/Y vssd1 vssd1 vccd1 vccd1 _13514_/B
+ sky130_fd_sc_hd__a22o_1
X_17281_ _17499_/A _17281_/B vssd1 vssd1 vccd1 vccd1 _17281_/X sky130_fd_sc_hd__xor2_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_161_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _26299_/CLK sky130_fd_sc_hd__clkbuf_16
X_14493_ _14491_/Y hold297/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold298/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_181_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19020_ _19018_/Y _18879_/X _19019_/X vssd1 vssd1 vccd1 vccd1 _19021_/A sky130_fd_sc_hd__a21o_1
X_16232_ _16473_/A hold957/X vssd1 vssd1 vccd1 vccd1 _16232_/Y sky130_fd_sc_hd__nand2_1
X_13444_ _13220_/A _14678_/A _13242_/A _25706_/Q vssd1 vssd1 vccd1 vccd1 _13444_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16163_ _16109_/A _16158_/A _16162_/Y vssd1 vssd1 vccd1 vccd1 _16171_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_180_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13375_ _18976_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13375_/X sky130_fd_sc_hd__or2_1
XFILLER_0_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15114_ _26005_/Q _25941_/Q _15773_/S vssd1 vssd1 vccd1 vccd1 _15115_/A sky130_fd_sc_hd__mux2_1
X_16094_ _16095_/B _16095_/A vssd1 vssd1 vccd1 vccd1 _16096_/A sky130_fd_sc_hd__or2_2
XFILLER_0_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15045_ _15051_/B _15046_/A vssd1 vssd1 vccd1 vccd1 _15045_/X sky130_fd_sc_hd__or2_1
X_19922_ _26270_/Q _19134_/X hold659/X vssd1 vssd1 vccd1 vccd1 _19923_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19853_ _19851_/Y _19852_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19853_/Y sky130_fd_sc_hd__a21oi_1
X_18804_ _19830_/A vssd1 vssd1 vccd1 vccd1 _22539_/B sky130_fd_sc_hd__inv_2
X_19784_ _26260_/Q _19134_/X hold671/X vssd1 vssd1 vccd1 vccd1 _19784_/Y sky130_fd_sc_hd__a21oi_1
X_16996_ _17688_/A _17683_/B _16996_/C vssd1 vssd1 vccd1 vccd1 _17794_/A sky130_fd_sc_hd__nand3_4
XFILLER_0_78_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15947_ hold880/X vssd1 vssd1 vccd1 vccd1 _15951_/B sky130_fd_sc_hd__inv_2
X_18735_ _20526_/B _22438_/A vssd1 vssd1 vccd1 vccd1 _20517_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_162_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18666_ _20401_/B _19729_/A vssd1 vssd1 vccd1 vccd1 _18667_/B sky130_fd_sc_hd__nand2_1
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15878_ hold461/X vssd1 vssd1 vccd1 vccd1 _15881_/B sky130_fd_sc_hd__inv_2
XFILLER_0_116_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14829_ _25852_/Q _13466_/A _14828_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14830_/A
+ sky130_fd_sc_hd__a22o_1
X_17617_ _17624_/A _17617_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _17617_/X sky130_fd_sc_hd__and3_1
XFILLER_0_58_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18597_ _19026_/A _18597_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18597_/X sky130_fd_sc_hd__and3_1
XFILLER_0_175_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17548_ _17548_/A _17600_/A vssd1 vssd1 vccd1 vccd1 _17549_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17479_ _17624_/A _17479_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17479_/X sky130_fd_sc_hd__and3_1
XFILLER_0_46_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_152_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _26301_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19218_ _20506_/A _19216_/Y _20511_/C vssd1 vssd1 vccd1 vccd1 _19308_/B sky130_fd_sc_hd__o21a_4
XFILLER_0_132_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20490_ _21563_/A vssd1 vssd1 vccd1 vccd1 _21562_/A sky130_fd_sc_hd__inv_2
XFILLER_0_85_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19149_ _22902_/B vssd1 vssd1 vccd1 vccd1 _19149_/X sky130_fd_sc_hd__buf_8
XFILLER_0_143_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22160_ _25787_/Q _22160_/B vssd1 vssd1 vccd1 vccd1 _22160_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_140_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21111_ _21545_/C _21594_/C vssd1 vssd1 vccd1 vccd1 _21114_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22091_ _22091_/A _22145_/B vssd1 vssd1 vccd1 vccd1 _22091_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21042_ _21042_/A _21042_/B _21041_/X vssd1 vssd1 vccd1 vccd1 _21043_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_160_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25850_ _26336_/CLK _25850_/D vssd1 vssd1 vccd1 vccd1 _25850_/Q sky130_fd_sc_hd__dfxtp_4
X_24801_ _24801_/A vssd1 vssd1 vccd1 vccd1 _26328_/D sky130_fd_sc_hd__clkbuf_1
X_25781_ _25781_/CLK _25781_/D vssd1 vssd1 vccd1 vccd1 _25781_/Q sky130_fd_sc_hd__dfxtp_2
X_22993_ _22993_/A _22993_/B vssd1 vssd1 vccd1 vccd1 _22994_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_119_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24732_ _24732_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24733_/A sky130_fd_sc_hd__and2_1
X_21944_ _21944_/A _21944_/B vssd1 vssd1 vccd1 vccd1 _23152_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_97_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24663_ _24663_/A vssd1 vssd1 vccd1 vccd1 _26283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_173_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21875_ _21875_/A _21875_/B vssd1 vssd1 vccd1 vccd1 _23120_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_96_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23614_ _23614_/A _23629_/B vssd1 vssd1 vccd1 vccd1 _23615_/A sky130_fd_sc_hd__and2_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20826_ _20826_/A _20826_/B vssd1 vssd1 vccd1 vccd1 _21435_/B sky130_fd_sc_hd__nand2_4
X_24594_ hold2739/X hold2738/X _24664_/S vssd1 vssd1 vccd1 vccd1 _24595_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26333_ _26334_/CLK _26333_/D vssd1 vssd1 vccd1 vccd1 _26333_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_49_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23545_ _24942_/S hold314/A _23544_/X vssd1 vssd1 vccd1 vccd1 _23545_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_181_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_143_clk clkbuf_4_11__f_clk/X vssd1 vssd1 vccd1 vccd1 _25812_/CLK sky130_fd_sc_hd__clkbuf_16
X_20757_ _20759_/B _20759_/C vssd1 vssd1 vccd1 vccd1 _20758_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_119_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26264_ _26264_/CLK _26264_/D vssd1 vssd1 vccd1 vccd1 _26264_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_18_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20688_ _21371_/B _21645_/B vssd1 vssd1 vccd1 vccd1 _20689_/C sky130_fd_sc_hd__nand2_1
X_23476_ _24956_/S hold311/A _23475_/X vssd1 vssd1 vccd1 vccd1 _23476_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25215_ _25797_/CLK hold556/X vssd1 vssd1 vccd1 vccd1 hold554/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22427_ _23001_/B _22423_/Y _22424_/X _22425_/X _22426_/Y vssd1 vssd1 vccd1 vccd1
+ _22427_/X sky130_fd_sc_hd__a32o_1
X_26195_ _26198_/CLK _26195_/D vssd1 vssd1 vccd1 vccd1 _26195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25146_ _25727_/CLK hold850/X vssd1 vssd1 vccd1 vccd1 hold849/A sky130_fd_sc_hd__dfxtp_1
X_13160_ _13049_/X _14536_/A _13067_/X _19230_/A vssd1 vssd1 vccd1 vccd1 _13160_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22358_ _22359_/A _22359_/C _23071_/A vssd1 vssd1 vccd1 vccd1 _22358_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13091_ _17864_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13091_/X sky130_fd_sc_hd__or2_1
X_21309_ _26315_/Q _21228_/X hold527/X vssd1 vssd1 vccd1 vccd1 _21312_/B sky130_fd_sc_hd__a21oi_1
X_22289_ _22265_/X _22288_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _22289_/Y sky130_fd_sc_hd__o21ai_1
X_25077_ _26164_/CLK hold991/X vssd1 vssd1 vccd1 vccd1 hold990/A sky130_fd_sc_hd__dfxtp_1
X_24028_ _24028_/A vssd1 vssd1 vccd1 vccd1 _26077_/D sky130_fd_sc_hd__clkbuf_1
Xhold290 hold290/A vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__dlygate4sd3_1
X_16850_ _16850_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16850_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15801_ _15789_/Y _15830_/B _15233_/X vssd1 vssd1 vccd1 vccd1 _15801_/Y sky130_fd_sc_hd__a21oi_1
X_16781_ _16980_/A _16781_/B vssd1 vssd1 vccd1 vccd1 _16781_/Y sky130_fd_sc_hd__nand2_1
X_25979_ _26042_/CLK _25979_/D vssd1 vssd1 vccd1 vccd1 _25979_/Q sky130_fd_sc_hd__dfxtp_1
X_13993_ hold657/X _13992_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold658/A sky130_fd_sc_hd__a21oi_1
X_18520_ _19630_/A vssd1 vssd1 vccd1 vccd1 _22179_/B sky130_fd_sc_hd__inv_2
X_15732_ _15720_/X _15764_/A _15233_/X vssd1 vssd1 vccd1 vccd1 _15732_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ _17464_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12944_/X sky130_fd_sc_hd__or2_1
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18451_ _21296_/B _22067_/A vssd1 vssd1 vccd1 vccd1 _21290_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_185_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15663_ _15661_/X _15662_/Y _15464_/X vssd1 vssd1 vccd1 vccd1 _25466_/D sky130_fd_sc_hd__a21oi_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _12840_/X _12873_/X _12827_/X _12874_/X vssd1 vssd1 vccd1 vccd1 _12875_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _17402_/A _17402_/B vssd1 vssd1 vccd1 vccd1 _17402_/X sky130_fd_sc_hd__xor2_1
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14614_ _14614_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14614_/Y sky130_fd_sc_hd__nand2_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _25873_/Q _21980_/A vssd1 vssd1 vccd1 vccd1 _18390_/A sky130_fd_sc_hd__or2_2
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _15592_/Y _15593_/Y _15464_/X vssd1 vssd1 vccd1 vccd1 hold909/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _17393_/A hold983/X _17572_/C vssd1 vssd1 vccd1 vccd1 _17333_/X sky130_fd_sc_hd__and3_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14545_ _14545_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14545_/Y sky130_fd_sc_hd__nand2_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_134_clk clkbuf_leaf_82_clk/A vssd1 vssd1 vccd1 vccd1 _25709_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17264_ _25641_/Q vssd1 vssd1 vccd1 vccd1 _20791_/B sky130_fd_sc_hd__inv_2
XFILLER_0_181_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14476_ _14476_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14476_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19003_ _19003_/A _19073_/B vssd1 vssd1 vccd1 vccd1 _19004_/B sky130_fd_sc_hd__xnor2_1
X_16215_ _16215_/A _16217_/A vssd1 vssd1 vccd1 vccd1 _16271_/B sky130_fd_sc_hd__and2_1
XFILLER_0_126_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13427_ _13427_/A vssd1 vssd1 vccd1 vccd1 _19844_/A sky130_fd_sc_hd__buf_6
XFILLER_0_52_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17195_ _25636_/Q vssd1 vssd1 vccd1 vccd1 _20597_/B sky130_fd_sc_hd__inv_2
XFILLER_0_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16146_ _16676_/A _16146_/B vssd1 vssd1 vccd1 vccd1 _16148_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_106_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ _13315_/X _13356_/X _13300_/X _13357_/X vssd1 vssd1 vccd1 vccd1 _13358_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16077_ _16074_/X hold549/X _16076_/X vssd1 vssd1 vccd1 vccd1 hold550/A sky130_fd_sc_hd__a21oi_1
X_13289_ _13289_/A vssd1 vssd1 vccd1 vccd1 _19532_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15028_ _15028_/A _15028_/B vssd1 vssd1 vccd1 vccd1 _15051_/A sky130_fd_sc_hd__nand2_1
X_19905_ _19903_/Y _19904_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19905_/Y sky130_fd_sc_hd__a21oi_1
Xhold2608 _26269_/Q vssd1 vssd1 vccd1 vccd1 hold2608/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2619 _24829_/X vssd1 vssd1 vccd1 vccd1 _24830_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19836_ _19834_/X _19835_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19836_/Y sky130_fd_sc_hd__a21oi_1
Xhold1907 _26023_/Q vssd1 vssd1 vccd1 vccd1 hold1907/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1918 _26324_/Q vssd1 vssd1 vccd1 vccd1 hold1918/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1929 _23850_/X vssd1 vssd1 vccd1 vccd1 _23851_/A sky130_fd_sc_hd__dlygate4sd3_1
X_19767_ _19757_/X _19765_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19767_/Y sky130_fd_sc_hd__o21ai_1
X_16979_ _23197_/B _13468_/X _16774_/Y vssd1 vssd1 vccd1 vccd1 _16979_/Y sky130_fd_sc_hd__a21oi_1
Xinput3 io_in[2] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
X_18718_ _18718_/A _18718_/B vssd1 vssd1 vccd1 vccd1 _18718_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_116_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19698_ _26254_/Q hold515/X vssd1 vssd1 vccd1 vccd1 _19698_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_91_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18649_ _18952_/A _25758_/Q _18891_/C vssd1 vssd1 vccd1 vccd1 _18650_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21660_ _21708_/B _21660_/B vssd1 vssd1 vccd1 vccd1 _21662_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20611_ _21338_/B _21611_/A vssd1 vssd1 vccd1 vccd1 _20613_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_129_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21591_ _21588_/Y _21590_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21591_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_125_clk clkbuf_4_11__f_clk/X vssd1 vssd1 vccd1 vccd1 _25689_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_117_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23330_ _23330_/A _23330_/B vssd1 vssd1 vccd1 vccd1 _23331_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_62_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20542_ _23199_/A vssd1 vssd1 vccd1 vccd1 _21125_/B sky130_fd_sc_hd__buf_6
XFILLER_0_149_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23261_ _23264_/A _23377_/B _23261_/C vssd1 vssd1 vccd1 vccd1 _23262_/A sky130_fd_sc_hd__and3_1
XFILLER_0_15_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20473_ _20475_/B _20475_/C vssd1 vssd1 vccd1 vccd1 _20474_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_172_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25000_ _26004_/CLK _25000_/D vssd1 vssd1 vccd1 vccd1 output8/A sky130_fd_sc_hd__dfxtp_4
XFILLER_0_131_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22212_ _25881_/Q _22213_/A vssd1 vssd1 vccd1 vccd1 _22214_/A sky130_fd_sc_hd__or2_1
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23192_ _23191_/A _22999_/C _23191_/B vssd1 vssd1 vccd1 vccd1 _23193_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22143_ _22141_/Y _22142_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _22143_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22074_ _22575_/A _22774_/B vssd1 vssd1 vccd1 vccd1 _22084_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_22_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25902_ _26269_/CLK _25902_/D vssd1 vssd1 vccd1 vccd1 _25902_/Q sky130_fd_sc_hd__dfxtp_2
X_21025_ _25866_/Q _21025_/B _21025_/C vssd1 vssd1 vccd1 vccd1 _21028_/C sky130_fd_sc_hd__nand3b_1
X_25833_ _25838_/CLK _25833_/D vssd1 vssd1 vccd1 vccd1 _25833_/Q sky130_fd_sc_hd__dfxtp_4
X_25764_ _25765_/CLK _25764_/D vssd1 vssd1 vccd1 vccd1 _25764_/Q sky130_fd_sc_hd__dfxtp_1
X_22976_ _22976_/A _22976_/B vssd1 vssd1 vccd1 vccd1 _22977_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24715_ _24715_/A vssd1 vssd1 vccd1 vccd1 _26300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21927_ _21928_/A _21928_/B _22977_/A vssd1 vssd1 vccd1 vccd1 _21927_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_167_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25695_ _26324_/CLK _25695_/D vssd1 vssd1 vccd1 vccd1 _25695_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12664_/B _12664_/A vssd1 vssd1 vccd1 vccd1 _12660_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_139_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24646_ _24646_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24647_/A sky130_fd_sc_hd__and2_1
X_21858_ _21859_/A _21859_/B _22943_/A vssd1 vssd1 vccd1 vccd1 _21858_/X sky130_fd_sc_hd__a21o_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20809_ _26297_/Q _20731_/X hold623/X vssd1 vssd1 vccd1 vccd1 _20812_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12591_ _12591_/A _23923_/A vssd1 vssd1 vccd1 vccd1 _12592_/C sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_116_clk clkbuf_4_14__f_clk/X vssd1 vssd1 vccd1 vccd1 _25418_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24577_ _24577_/A vssd1 vssd1 vccd1 vccd1 _26255_/D sky130_fd_sc_hd__clkbuf_1
X_21789_ _21789_/A vssd1 vssd1 vccd1 vccd1 _21789_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_182_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14330_ _14328_/Y hold207/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold208/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26316_ _26317_/CLK _26316_/D vssd1 vssd1 vccd1 vccd1 _26316_/Q sky130_fd_sc_hd__dfxtp_1
X_23528_ _24944_/S hold176/A _23527_/X vssd1 vssd1 vccd1 vccd1 _23528_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14261_ _25837_/Q vssd1 vssd1 vccd1 vccd1 _18956_/B sky130_fd_sc_hd__inv_2
X_26247_ _26248_/CLK _26247_/D vssd1 vssd1 vccd1 vccd1 _26247_/Q sky130_fd_sc_hd__dfxtp_2
X_23459_ hold17/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23459_/X sky130_fd_sc_hd__or2b_1
X_16000_ _16000_/A _16000_/B vssd1 vssd1 vccd1 vccd1 _16054_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_150_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13212_ _18475_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13212_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14192_ _14264_/A _14192_/B vssd1 vssd1 vccd1 vccd1 _14192_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_33_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26178_ _26181_/CLK _26178_/D vssd1 vssd1 vccd1 vccd1 _26178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25129_ _25249_/CLK _25129_/D vssd1 vssd1 vccd1 vccd1 _25129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13143_ _26160_/Q _13065_/X _13142_/X vssd1 vssd1 vccd1 vccd1 _13143_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_103_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17951_ _17951_/A _17951_/B vssd1 vssd1 vccd1 vccd1 _21763_/A sky130_fd_sc_hd__nand2_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _26147_/Q _13065_/X _13073_/X vssd1 vssd1 vccd1 vccd1 _13074_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_104_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16902_ _16935_/A _25569_/Q vssd1 vssd1 vccd1 vccd1 _16904_/B sky130_fd_sc_hd__nand2_1
X_17882_ _20111_/A _17882_/B vssd1 vssd1 vccd1 vccd1 _19114_/A sky130_fd_sc_hd__nand2_2
X_19621_ _19621_/A _19621_/B vssd1 vssd1 vccd1 vccd1 _19621_/Y sky130_fd_sc_hd__nand2_1
X_16833_ _16833_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16833_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_40_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16764_ _16858_/A _16764_/B vssd1 vssd1 vccd1 vccd1 _16764_/Y sky130_fd_sc_hd__nand2_1
X_19552_ _19550_/X _19551_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19552_/Y sky130_fd_sc_hd__a21oi_1
X_13976_ _17814_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13976_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_189_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15715_ _15718_/B _15716_/A vssd1 vssd1 vccd1 vccd1 _15715_/X sky130_fd_sc_hd__or2_1
X_18503_ _18503_/A _18503_/B vssd1 vssd1 vccd1 vccd1 _22148_/A sky130_fd_sc_hd__nand2_1
X_12927_ _26119_/Q _12907_/X _12926_/X vssd1 vssd1 vccd1 vccd1 _12927_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_186_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16695_ _16695_/A _16695_/B _16695_/C vssd1 vssd1 vccd1 vccd1 _16696_/B sky130_fd_sc_hd__nand3_1
X_19483_ _19483_/A vssd1 vssd1 vccd1 vccd1 _19483_/X sky130_fd_sc_hd__clkbuf_8
X_15646_ hold2489/X _15645_/Y _15464_/X vssd1 vssd1 vccd1 vccd1 _15646_/Y sky130_fd_sc_hd__a21oi_1
X_18434_ _18434_/A _18434_/B vssd1 vssd1 vccd1 vccd1 _18434_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_158_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12858_ _26106_/Q _12748_/X _12857_/X vssd1 vssd1 vccd1 vccd1 _12858_/X sky130_fd_sc_hd__a21o_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18365_ _18365_/A _21208_/B _18365_/C vssd1 vssd1 vccd1 vccd1 _21189_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_185_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15577_ _15577_/A _15577_/B vssd1 vssd1 vccd1 vccd1 _15611_/A sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_107_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _24983_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12789_ _12726_/B _14313_/A _12752_/X _25590_/Q vssd1 vssd1 vccd1 vccd1 _12789_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17316_ _19444_/A _17316_/B vssd1 vssd1 vccd1 vccd1 _17571_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_185_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14528_ _14588_/A vssd1 vssd1 vccd1 vccd1 _14584_/B sky130_fd_sc_hd__buf_4
X_18296_ _18641_/A _19216_/A vssd1 vssd1 vccd1 vccd1 _18296_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17247_ _17245_/Y _17246_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _17247_/Y sky130_fd_sc_hd__a21oi_1
X_14459_ _14465_/A hold224/X vssd1 vssd1 vccd1 vccd1 hold225/A sky130_fd_sc_hd__nand2_1
XFILLER_0_141_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17178_ _17176_/Y _17177_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _17178_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16129_ _16212_/A hold644/X vssd1 vssd1 vccd1 vccd1 hold645/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2405 _24338_/X vssd1 vssd1 vccd1 vccd1 _24339_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2416 _25668_/Q vssd1 vssd1 vccd1 vccd1 _13208_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2427 _24968_/Q vssd1 vssd1 vccd1 vccd1 _12575_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2438 _23998_/X vssd1 vssd1 vccd1 vccd1 _23999_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2449 _26069_/Q vssd1 vssd1 vccd1 vccd1 hold2449/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1704 _21688_/Y vssd1 vssd1 vccd1 vccd1 _25835_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1715 _25795_/Q vssd1 vssd1 vccd1 vccd1 _20853_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1726 _22434_/Y vssd1 vssd1 vccd1 vccd1 _25861_/D sky130_fd_sc_hd__dlygate4sd3_1
X_19819_ _19835_/B _19901_/B vssd1 vssd1 vccd1 vccd1 _19821_/A sky130_fd_sc_hd__xnor2_1
Xhold1737 _20505_/Y vssd1 vssd1 vccd1 vccd1 _25786_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1748 _17231_/Y vssd1 vssd1 vccd1 vccd1 _25597_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1759 _25826_/Q vssd1 vssd1 vccd1 vccd1 _21541_/B sky130_fd_sc_hd__dlygate4sd3_1
X_22830_ _15420_/B _22680_/X _22829_/X vssd1 vssd1 vccd1 vccd1 _22830_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22761_ _22909_/A _22761_/B vssd1 vssd1 vccd1 vccd1 _22762_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24500_ _24500_/A vssd1 vssd1 vccd1 vccd1 _26230_/D sky130_fd_sc_hd__clkbuf_1
X_21712_ _21712_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _21717_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_176_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25480_ _25495_/CLK hold655/X vssd1 vssd1 vccd1 vccd1 hold653/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22692_ _25836_/Q _22692_/B vssd1 vssd1 vccd1 vccd1 _22692_/Y sky130_fd_sc_hd__nor2_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24431_ _24431_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24432_/A sky130_fd_sc_hd__and2_1
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21643_ _21643_/A _21643_/B _21643_/C vssd1 vssd1 vccd1 vccd1 _21647_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_35_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24362_ _24362_/A vssd1 vssd1 vccd1 vccd1 _26185_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21574_ _21572_/Y _21573_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21574_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_30 _19031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_52 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26101_ _26103_/CLK _26101_/D vssd1 vssd1 vccd1 vccd1 _26101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23313_ hold896/X _23314_/A vssd1 vssd1 vccd1 vccd1 _23313_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_63 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20525_ _20525_/A _20525_/B vssd1 vssd1 vccd1 vccd1 _20527_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24293_ hold1949/X _26163_/Q _24356_/S vssd1 vssd1 vccd1 vccd1 _24293_/X sky130_fd_sc_hd__mux2_1
XANTENNA_74 _18899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26032_ _26032_/CLK _26032_/D vssd1 vssd1 vccd1 vccd1 _26032_/Q sky130_fd_sc_hd__dfxtp_1
X_23244_ _24950_/B _23244_/B vssd1 vssd1 vccd1 vccd1 _23249_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_160_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20456_ _20456_/A _20456_/B vssd1 vssd1 vccd1 vccd1 _20457_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_132_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23175_ _23175_/A _23175_/B _23191_/C vssd1 vssd1 vccd1 vccd1 _23177_/A sky130_fd_sc_hd__or3_1
XFILLER_0_127_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20387_ _20660_/A _20387_/B vssd1 vssd1 vccd1 vccd1 _20387_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22126_ _22126_/A _22126_/B vssd1 vssd1 vccd1 vccd1 _22807_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_101_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22057_ _22038_/X _22056_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _22057_/Y sky130_fd_sc_hd__o21ai_1
X_21008_ _21480_/C _21532_/B vssd1 vssd1 vccd1 vccd1 _21010_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_173_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25816_ _25835_/CLK _25816_/D vssd1 vssd1 vccd1 vccd1 _25816_/Q sky130_fd_sc_hd__dfxtp_2
X_13830_ _13941_/A _13830_/B vssd1 vssd1 vccd1 vccd1 _13830_/Y sky130_fd_sc_hd__nand2_1
X_25747_ _25752_/CLK _25747_/D vssd1 vssd1 vccd1 vccd1 _25747_/Q sky130_fd_sc_hd__dfxtp_1
X_13761_ _25757_/Q vssd1 vssd1 vccd1 vccd1 _18632_/B sky130_fd_sc_hd__inv_2
XFILLER_0_134_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22959_ _22959_/A _22959_/B vssd1 vssd1 vccd1 vccd1 _22960_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15500_ _15500_/A _15500_/B vssd1 vssd1 vccd1 vccd1 _15500_/Y sky130_fd_sc_hd__nand2_1
X_12712_ _12712_/A _12712_/B vssd1 vssd1 vccd1 vccd1 _12713_/D sky130_fd_sc_hd__nand2_1
X_16480_ _16480_/A _16492_/A vssd1 vssd1 vccd1 vccd1 _16481_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_167_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25678_ _25678_/CLK _25678_/D vssd1 vssd1 vccd1 vccd1 _25678_/Q sky130_fd_sc_hd__dfxtp_1
X_13692_ hold402/X _13691_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold403/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15431_ _15429_/X hold2300/X _15090_/X vssd1 vssd1 vccd1 vccd1 _15431_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12643_ hold868/X _12643_/B vssd1 vssd1 vccd1 vccd1 _12644_/C sky130_fd_sc_hd__nand2_1
X_24629_ _24629_/A vssd1 vssd1 vccd1 vccd1 _26272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18150_ _20310_/B _25654_/Q vssd1 vssd1 vccd1 vccd1 _18150_/Y sky130_fd_sc_hd__nand2_1
X_15362_ hold2041/X _15361_/Y _15090_/X vssd1 vssd1 vccd1 vccd1 _15362_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12574_ _12574_/A _23596_/B vssd1 vssd1 vccd1 vccd1 _12574_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_38_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17101_ _25595_/Q vssd1 vssd1 vccd1 vccd1 _20507_/B sky130_fd_sc_hd__inv_2
XFILLER_0_109_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14313_ _14313_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14313_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18081_ _25854_/Q _22247_/A vssd1 vssd1 vccd1 vccd1 _18089_/A sky130_fd_sc_hd__or2_2
X_15293_ _15307_/A _15294_/A vssd1 vssd1 vccd1 vccd1 _15293_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17032_ _17272_/A _17032_/B vssd1 vssd1 vccd1 vccd1 _17032_/Y sky130_fd_sc_hd__nand2_1
X_14244_ _18895_/B _14262_/B vssd1 vssd1 vccd1 vccd1 _14244_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_68_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14175_ hold441/X _14174_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold442/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13126_ _13049_/X _14515_/A _13067_/X _25654_/Q vssd1 vssd1 vccd1 vccd1 _13126_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ _19026_/A _18983_/B _22786_/A vssd1 vssd1 vccd1 vccd1 _18983_/X sky130_fd_sc_hd__and3_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ _17934_/A vssd1 vssd1 vccd1 vccd1 _19039_/A sky130_fd_sc_hd__clkinv_4
X_13057_ _26144_/Q _12907_/X _13056_/X vssd1 vssd1 vccd1 vccd1 _13057_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17865_ _17863_/Y _17528_/X _17864_/X vssd1 vssd1 vccd1 vccd1 _17866_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_75_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19604_ _20054_/A _19602_/Y _20058_/C vssd1 vssd1 vccd1 vccd1 _19692_/B sky130_fd_sc_hd__o21a_2
X_16816_ _16817_/B _16817_/A vssd1 vssd1 vccd1 vccd1 _16816_/X sky130_fd_sc_hd__or2_1
X_17796_ _17796_/A _20426_/B _17796_/C vssd1 vssd1 vccd1 vccd1 _20396_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19535_ _19551_/B _19621_/B vssd1 vssd1 vccd1 vccd1 _19537_/A sky130_fd_sc_hd__xnor2_1
X_16747_ _16747_/A _16747_/B vssd1 vssd1 vccd1 vccd1 _16747_/Y sky130_fd_sc_hd__nand2_1
X_13959_ _26291_/Q _13801_/X _13793_/X _13958_/Y vssd1 vssd1 vccd1 vccd1 _13960_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16678_ _16678_/A _16678_/B vssd1 vssd1 vccd1 vccd1 _16679_/B sky130_fd_sc_hd__nand2_1
X_19466_ _22586_/A vssd1 vssd1 vccd1 vccd1 _19723_/A sky130_fd_sc_hd__buf_6
XFILLER_0_159_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18417_ _18417_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18417_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15629_ _15956_/A hold946/X vssd1 vssd1 vccd1 vccd1 _15629_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_146_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19397_ _19395_/Y _19396_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19397_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18348_ _18348_/A _18348_/B _18348_/C vssd1 vssd1 vccd1 vccd1 _21915_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_185_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18279_ _18279_/A _18279_/B vssd1 vssd1 vccd1 vccd1 _21809_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_140_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20310_ _20310_/A _20310_/B vssd1 vssd1 vccd1 vccd1 _20314_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_115_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21290_ _21290_/A _22065_/B vssd1 vssd1 vccd1 vccd1 _21291_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_142_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold801 hold801/A vssd1 vssd1 vccd1 vccd1 hold801/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold812 hold812/A vssd1 vssd1 vccd1 vccd1 hold812/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 hold823/A vssd1 vssd1 vccd1 vccd1 hold823/X sky130_fd_sc_hd__buf_1
XFILLER_0_4_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20241_ _20244_/A _20244_/C vssd1 vssd1 vccd1 vccd1 _20243_/A sky130_fd_sc_hd__nand2_1
Xhold834 hold834/A vssd1 vssd1 vccd1 vccd1 hold834/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold845 hold845/A vssd1 vssd1 vccd1 vccd1 hold845/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 hold856/A vssd1 vssd1 vccd1 vccd1 hold856/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 hold867/A vssd1 vssd1 vccd1 vccd1 hold867/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 hold878/A vssd1 vssd1 vccd1 vccd1 hold878/X sky130_fd_sc_hd__buf_1
XFILLER_0_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20172_ _20172_/A _20172_/B vssd1 vssd1 vccd1 vccd1 _21434_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold889 hold889/A vssd1 vssd1 vccd1 vccd1 hold889/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2202 _25928_/Q vssd1 vssd1 vccd1 vccd1 _23327_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24980_ _24983_/CLK _24980_/D vssd1 vssd1 vccd1 vccd1 _24980_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2213 _25987_/Q vssd1 vssd1 vccd1 vccd1 _14752_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2224 _25961_/Q vssd1 vssd1 vccd1 vccd1 hold2224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2235 _26153_/Q vssd1 vssd1 vccd1 vccd1 hold2235/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2246 _25423_/Q vssd1 vssd1 vccd1 vccd1 _14989_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1501 _25891_/Q vssd1 vssd1 vccd1 vccd1 _23037_/B sky130_fd_sc_hd__buf_1
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23931_ _23931_/A vssd1 vssd1 vccd1 vccd1 _26045_/D sky130_fd_sc_hd__clkbuf_1
Xhold1512 _20086_/Y vssd1 vssd1 vccd1 vccd1 _25775_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2257 _26109_/Q vssd1 vssd1 vccd1 vccd1 hold2257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1523 _25900_/Q vssd1 vssd1 vccd1 vccd1 _23181_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2268 _26137_/Q vssd1 vssd1 vccd1 vccd1 hold2268/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 _13388_/X vssd1 vssd1 vccd1 vccd1 _25116_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2279 _26108_/Q vssd1 vssd1 vccd1 vccd1 hold2279/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1545 _25115_/Q vssd1 vssd1 vccd1 vccd1 _18983_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1556 _21494_/Y vssd1 vssd1 vccd1 vccd1 _25823_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23862_ hold2343/X hold2193/X _23907_/S vssd1 vssd1 vccd1 vccd1 _23863_/A sky130_fd_sc_hd__mux2_1
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1567 _21381_/Y vssd1 vssd1 vccd1 vccd1 _25816_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1578 _25888_/Q vssd1 vssd1 vccd1 vccd1 _22988_/B sky130_fd_sc_hd__buf_1
X_25601_ _26231_/CLK _25601_/D vssd1 vssd1 vccd1 vccd1 _25601_/Q sky130_fd_sc_hd__dfxtp_2
Xhold1589 _21477_/Y vssd1 vssd1 vccd1 vccd1 _25822_/D sky130_fd_sc_hd__dlygate4sd3_1
X_22813_ _15398_/B _22680_/X _14273_/X vssd1 vssd1 vccd1 vccd1 _22813_/Y sky130_fd_sc_hd__a21oi_1
X_23793_ _23793_/A vssd1 vssd1 vccd1 vccd1 _26002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25532_ _25532_/CLK hold872/X vssd1 vssd1 vccd1 vccd1 hold871/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22744_ _22744_/A _22744_/B vssd1 vssd1 vccd1 vccd1 _22745_/B sky130_fd_sc_hd__nand2_1
X_25463_ _26009_/CLK _25463_/D vssd1 vssd1 vccd1 vccd1 _25463_/Q sky130_fd_sc_hd__dfxtp_1
Xascon_wrapper_14 vssd1 vssd1 vccd1 vccd1 io_oeb[0] ascon_wrapper_14/LO sky130_fd_sc_hd__conb_1
XFILLER_0_181_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22675_ _22675_/A _22675_/B vssd1 vssd1 vccd1 vccd1 _22676_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24414_ _24414_/A vssd1 vssd1 vccd1 vccd1 _26202_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21626_ _21628_/B _21677_/B vssd1 vssd1 vccd1 vccd1 _21627_/B sky130_fd_sc_hd__nand2_1
X_25394_ _25991_/CLK _25394_/D vssd1 vssd1 vccd1 vccd1 _25394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24345_ _24345_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24346_/A sky130_fd_sc_hd__and2_1
X_21557_ _21573_/A _21557_/B vssd1 vssd1 vccd1 vccd1 _21557_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_133_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20508_ _20511_/A _20511_/C vssd1 vssd1 vccd1 vccd1 _20509_/A sky130_fd_sc_hd__nand2_1
X_24276_ hold1985/X _26158_/Q _24279_/S vssd1 vssd1 vccd1 vccd1 _24276_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_105_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21488_ _21487_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21488_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26015_ _26021_/CLK _26015_/D vssd1 vssd1 vccd1 vccd1 _26015_/Q sky130_fd_sc_hd__dfxtp_1
X_23227_ _23227_/A _24946_/A vssd1 vssd1 vccd1 vccd1 _23228_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_120_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20439_ _20439_/A _20439_/B vssd1 vssd1 vccd1 vccd1 _20443_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_120_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23158_ _26082_/Q vssd1 vssd1 vccd1 vccd1 _23159_/A sky130_fd_sc_hd__inv_2
X_22109_ _22110_/A _22110_/C _23074_/A vssd1 vssd1 vccd1 vccd1 _22109_/X sky130_fd_sc_hd__a21o_1
X_15980_ _16212_/A hold809/X vssd1 vssd1 vccd1 vccd1 hold810/A sky130_fd_sc_hd__nand2_1
X_23089_ _23089_/A _23089_/B vssd1 vssd1 vccd1 vccd1 _23090_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14931_ _14931_/A _14931_/B vssd1 vssd1 vccd1 vccd1 _14932_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_175_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14862_ _14862_/A vssd1 vssd1 vccd1 vccd1 _15049_/A sky130_fd_sc_hd__inv_2
X_17650_ _17648_/Y _17649_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _25644_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16601_ _16554_/B _16598_/A _16600_/X vssd1 vssd1 vccd1 vccd1 _16602_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_138_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13813_ _13880_/A hold677/X vssd1 vssd1 vccd1 vccd1 hold678/A sky130_fd_sc_hd__nand2_1
XFILLER_0_188_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17581_ _17578_/X _17528_/X _17580_/X vssd1 vssd1 vccd1 vccd1 _17582_/A sky130_fd_sc_hd__a21o_1
X_14793_ _25848_/Q _13466_/A _14792_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14794_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16532_ _16676_/A _16532_/B vssd1 vssd1 vccd1 vccd1 _16534_/A sky130_fd_sc_hd__nor2_1
X_19320_ _19336_/B _19407_/B vssd1 vssd1 vccd1 vccd1 _19322_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13744_ _18571_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13744_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16463_ hold970/X vssd1 vssd1 vccd1 vccd1 _16466_/B sky130_fd_sc_hd__inv_2
XFILLER_0_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19251_ _26222_/Q _19483_/A hold533/X vssd1 vssd1 vccd1 vccd1 _19252_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_167_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13675_ _25743_/Q vssd1 vssd1 vccd1 vccd1 _18347_/B sky130_fd_sc_hd__inv_2
XFILLER_0_39_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15414_ _15414_/A _15443_/A vssd1 vssd1 vccd1 vccd1 _15414_/Y sky130_fd_sc_hd__nand2_1
X_18202_ _18612_/A _18202_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18203_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_155_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12626_ _12626_/A vssd1 vssd1 vccd1 vccd1 _24978_/D sky130_fd_sc_hd__clkbuf_1
X_19182_ _19983_/B _19183_/A vssd1 vssd1 vccd1 vccd1 _19182_/X sky130_fd_sc_hd__or2_1
X_16394_ _16394_/A _16394_/B vssd1 vssd1 vccd1 vccd1 _16404_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_171_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18133_ _25862_/Q _21903_/A vssd1 vssd1 vccd1 vccd1 _18141_/A sky130_fd_sc_hd__or2_2
X_15345_ _15956_/A hold975/X vssd1 vssd1 vccd1 vccd1 _15345_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_170_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12557_ _17674_/A _12549_/X hold1840/X _12551_/Y _12556_/X vssd1 vssd1 vccd1 vccd1
+ _12557_/X sky130_fd_sc_hd__o2111a_1
XFILLER_0_182_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18064_ _25652_/Q vssd1 vssd1 vccd1 vccd1 _21958_/A sky130_fd_sc_hd__inv_2
X_15276_ _15111_/Y _15271_/X _15275_/Y vssd1 vssd1 vccd1 vccd1 _15277_/B sky130_fd_sc_hd__a21oi_1
X_12488_ _15839_/A _12496_/A vssd1 vssd1 vccd1 vccd1 _14270_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_184_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 hold108/A vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__dlygate4sd3_1
X_17015_ _19199_/A vssd1 vssd1 vccd1 vccd1 _17272_/A sky130_fd_sc_hd__clkbuf_8
X_14227_ _26334_/Q _13518_/B _14170_/X _14226_/Y vssd1 vssd1 vccd1 vccd1 _14228_/B
+ sky130_fd_sc_hd__a22o_1
Xhold119 hold119/A vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14158_ _25820_/Q vssd1 vssd1 vccd1 vccd1 _18613_/B sky130_fd_sc_hd__inv_2
XFILLER_0_81_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _14260_/A vssd1 vssd1 vccd1 vccd1 _13109_/X sky130_fd_sc_hd__buf_6
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ _25809_/Q vssd1 vssd1 vccd1 vccd1 _18388_/B sky130_fd_sc_hd__inv_2
X_18966_ _18966_/A _19038_/B vssd1 vssd1 vccd1 vccd1 _18967_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ _18252_/A _17917_/B vssd1 vssd1 vccd1 vccd1 _17917_/Y sky130_fd_sc_hd__nand2_1
X_18897_ _18897_/A _20828_/A vssd1 vssd1 vccd1 vccd1 _19059_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17848_ _20707_/B _22310_/A vssd1 vssd1 vccd1 vccd1 _20701_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_179_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17779_ _17779_/A _17779_/B vssd1 vssd1 vccd1 vccd1 _17780_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19518_ _19518_/A _21184_/B vssd1 vssd1 vccd1 vccd1 _19518_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_77_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20790_ _20790_/A _22615_/B vssd1 vssd1 vccd1 vccd1 _20791_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19449_ _19449_/A _19449_/B vssd1 vssd1 vccd1 vccd1 _19449_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22460_ _22561_/A _22460_/B vssd1 vssd1 vccd1 vccd1 _22460_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21411_ _21411_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21411_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22391_ _25824_/Q _22391_/B vssd1 vssd1 vccd1 vccd1 _22391_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_60_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24130_ hold2257/X hold2252/X _24203_/S vssd1 vssd1 vccd1 vccd1 _24131_/A sky130_fd_sc_hd__mux2_1
X_21342_ _26317_/Q hold821/X vssd1 vssd1 vccd1 vccd1 _21342_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_114_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24061_ _24061_/A vssd1 vssd1 vccd1 vccd1 _26087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold620 hold620/A vssd1 vssd1 vccd1 vccd1 hold620/X sky130_fd_sc_hd__dlygate4sd3_1
X_21273_ _21646_/B _21691_/C vssd1 vssd1 vccd1 vccd1 _21276_/A sky130_fd_sc_hd__nand2_1
Xhold631 hold631/A vssd1 vssd1 vccd1 vccd1 hold631/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold642 hold642/A vssd1 vssd1 vccd1 vccd1 hold642/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 hold653/A vssd1 vssd1 vccd1 vccd1 hold653/X sky130_fd_sc_hd__dlygate4sd3_1
X_23012_ _23188_/A _23012_/B vssd1 vssd1 vccd1 vccd1 _23012_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20224_ _20224_/A _20224_/B _21010_/B vssd1 vssd1 vccd1 vccd1 _20225_/B sky130_fd_sc_hd__nand3_1
Xhold664 hold664/A vssd1 vssd1 vccd1 vccd1 hold664/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 hold675/A vssd1 vssd1 vccd1 vccd1 hold675/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold686 hold686/A vssd1 vssd1 vccd1 vccd1 hold686/X sky130_fd_sc_hd__buf_1
Xhold697 hold697/A vssd1 vssd1 vccd1 vccd1 hold697/X sky130_fd_sc_hd__dlygate4sd3_1
X_20155_ _26280_/Q hold851/X vssd1 vssd1 vccd1 vccd1 _20155_/Y sky130_fd_sc_hd__nand2_1
Xhold2010 _24994_/Q vssd1 vssd1 vccd1 vccd1 hold2010/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2021 _23338_/X vssd1 vssd1 vccd1 vccd1 _23339_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold2032 _26011_/Q vssd1 vssd1 vccd1 vccd1 hold2032/X sky130_fd_sc_hd__dlygate4sd3_1
X_24963_ _24909_/X _23593_/X _24910_/X _24961_/X hold1982/X vssd1 vssd1 vccd1 vccd1
+ _24963_/X sky130_fd_sc_hd__a41o_1
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2043 _26026_/Q vssd1 vssd1 vccd1 vccd1 hold2043/X sky130_fd_sc_hd__dlygate4sd3_1
X_20086_ _20084_/Y _20085_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _20086_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2054 _23992_/X vssd1 vssd1 vccd1 vccd1 _23993_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_96_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _25999_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold2065 _14935_/Y vssd1 vssd1 vccd1 vccd1 hold2065/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1320 hold2758/X vssd1 vssd1 vccd1 vccd1 _23021_/B sky130_fd_sc_hd__clkbuf_2
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1331 _25578_/Q vssd1 vssd1 vccd1 vccd1 _16970_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2076 _23880_/X vssd1 vssd1 vccd1 vccd1 _23881_/A sky130_fd_sc_hd__dlygate4sd3_1
X_23914_ hold1934/X _26042_/Q _23920_/S vssd1 vssd1 vccd1 vccd1 _23914_/X sky130_fd_sc_hd__mux2_1
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2087 _25993_/Q vssd1 vssd1 vccd1 vccd1 _14806_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1342 _23050_/X vssd1 vssd1 vccd1 vccd1 _23051_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2098 _25936_/Q vssd1 vssd1 vccd1 vccd1 _23363_/A sky130_fd_sc_hd__dlygate4sd3_1
X_24894_ _15730_/A _15745_/A _24945_/S vssd1 vssd1 vccd1 vccd1 _24894_/X sky130_fd_sc_hd__mux2_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1353 _25754_/Q vssd1 vssd1 vccd1 vccd1 _19752_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1364 _19988_/Y vssd1 vssd1 vccd1 vccd1 _25772_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1375 _25779_/Q vssd1 vssd1 vccd1 vccd1 _20233_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1386 _19312_/Y vssd1 vssd1 vccd1 vccd1 _25723_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23845_ _23845_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23846_/A sky130_fd_sc_hd__and2_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1397 _25774_/Q vssd1 vssd1 vccd1 vccd1 _20041_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23776_ hold2216/X _25997_/Q _23831_/S vssd1 vssd1 vccd1 vccd1 _23776_/X sky130_fd_sc_hd__mux2_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20988_ _21042_/A _20988_/B _20987_/X vssd1 vssd1 vccd1 vccd1 _20989_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25515_ _25515_/CLK hold915/X vssd1 vssd1 vccd1 vccd1 hold914/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22727_ _23039_/A _23184_/B vssd1 vssd1 vccd1 vccd1 _22728_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25446_ _26052_/CLK _25446_/D vssd1 vssd1 vccd1 vccd1 _25446_/Q sky130_fd_sc_hd__dfxtp_1
X_13460_ _26212_/Q _13426_/X _13459_/X vssd1 vssd1 vccd1 vccd1 _13460_/X sky130_fd_sc_hd__a21o_1
X_22658_ _22658_/A _23001_/B _22658_/C vssd1 vssd1 vccd1 vccd1 _22658_/X sky130_fd_sc_hd__and3_1
XFILLER_0_125_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21609_ _21611_/A _21661_/B vssd1 vssd1 vccd1 vccd1 _21610_/B sky130_fd_sc_hd__nand2_1
X_25377_ _25418_/CLK hold169/X vssd1 vssd1 vccd1 vccd1 hold167/A sky130_fd_sc_hd__dfxtp_1
X_13391_ _13220_/X _14651_/A _13242_/X _19758_/A vssd1 vssd1 vccd1 vccd1 _13391_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22589_ _22589_/A _25896_/Q vssd1 vssd1 vccd1 vccd1 _22589_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_20_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _26154_/CLK sky130_fd_sc_hd__clkbuf_16
X_15130_ _16231_/A vssd1 vssd1 vccd1 vccd1 _15956_/A sky130_fd_sc_hd__buf_8
XFILLER_0_90_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24328_ _24328_/A vssd1 vssd1 vccd1 vccd1 _26174_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15061_ _15067_/B _15062_/A vssd1 vssd1 vccd1 vccd1 _15061_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24259_ _24259_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24260_/A sky130_fd_sc_hd__and2_1
XFILLER_0_121_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14012_ _14061_/A _14012_/B vssd1 vssd1 vccd1 vccd1 _14012_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_142_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18820_ _18818_/X _18269_/X _18819_/X vssd1 vssd1 vccd1 vccd1 _18821_/A sky130_fd_sc_hd__a21o_1
X_18751_ _18751_/A _25827_/Q _18751_/C vssd1 vssd1 vccd1 vccd1 _20566_/B sky130_fd_sc_hd__nand3_2
X_15963_ _15963_/A _16000_/A vssd1 vssd1 vccd1 vccd1 _15963_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_65_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_87_clk clkbuf_leaf_95_clk/A vssd1 vssd1 vccd1 vccd1 _26051_/CLK sky130_fd_sc_hd__clkbuf_16
X_17702_ _23208_/B _17752_/B _17719_/B vssd1 vssd1 vccd1 vccd1 _17704_/A sky130_fd_sc_hd__o21a_1
X_14914_ _14914_/A _14925_/B vssd1 vssd1 vccd1 vccd1 _14915_/A sky130_fd_sc_hd__nand2_1
X_15894_ _15894_/A _15894_/B vssd1 vssd1 vccd1 vccd1 _15895_/A sky130_fd_sc_hd__nor2_1
X_18682_ _18986_/A _19488_/A vssd1 vssd1 vccd1 vccd1 _18682_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_76_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17633_ _17630_/X _17528_/X _17632_/X vssd1 vssd1 vccd1 vccd1 _17634_/A sky130_fd_sc_hd__a21o_1
X_14845_ _22232_/B _15543_/B vssd1 vssd1 vccd1 vccd1 _14846_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14776_ _14776_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14776_/Y sky130_fd_sc_hd__nand2_1
X_17564_ _17624_/A _17564_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17564_/X sky130_fd_sc_hd__and3_1
XFILLER_0_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19303_ _19303_/A _20741_/B vssd1 vssd1 vccd1 vccd1 _19303_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16515_ _16515_/A _16524_/B vssd1 vssd1 vccd1 vccd1 _16515_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13727_ _26254_/Q _13612_/X _13605_/X _13726_/Y vssd1 vssd1 vccd1 vccd1 _13728_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17495_ _17495_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17495_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19234_ _19234_/A _19234_/B vssd1 vssd1 vccd1 vccd1 _19234_/X sky130_fd_sc_hd__xor2_1
X_16446_ _16462_/A _16461_/A vssd1 vssd1 vccd1 vccd1 _16447_/C sky130_fd_sc_hd__nand2_1
X_13658_ _18287_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13658_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_186_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _12610_/A _24974_/Q hold868/X vssd1 vssd1 vccd1 vccd1 hold869/A sky130_fd_sc_hd__a21oi_1
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16377_ _16375_/X _16376_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 hold915/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19165_ _19983_/B _19248_/A vssd1 vssd1 vccd1 vccd1 _19167_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13589_ _26232_/Q _13426_/X _13468_/X _13588_/Y vssd1 vssd1 vccd1 vccd1 _13590_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk _25184_/CLK vssd1 vssd1 vccd1 vccd1 _26267_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15328_ _15328_/A vssd1 vssd1 vccd1 vccd1 _15407_/B sky130_fd_sc_hd__inv_2
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18116_ _25653_/Q _20285_/B vssd1 vssd1 vccd1 vccd1 _18117_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_81_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19096_ _19092_/Y _17828_/B _19095_/Y vssd1 vssd1 vccd1 vccd1 _19950_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_112_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15259_ _15795_/A _16282_/B vssd1 vssd1 vccd1 vccd1 _15262_/A sky130_fd_sc_hd__nor2_1
X_18047_ _18047_/A _20880_/B _18047_/C vssd1 vssd1 vccd1 vccd1 _20862_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19998_ _19996_/Y _19997_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _19998_/Y sky130_fd_sc_hd__a21oi_1
X_18949_ _18949_/A _18949_/B vssd1 vssd1 vccd1 vccd1 _22717_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_78_clk clkbuf_leaf_82_clk/A vssd1 vssd1 vccd1 vccd1 _25865_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_146_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21960_ _21960_/A _21960_/B vssd1 vssd1 vccd1 vccd1 _22994_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_94_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20911_ _20911_/A _25862_/Q vssd1 vssd1 vccd1 vccd1 _20916_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21891_ _21891_/A _21891_/B vssd1 vssd1 vccd1 vccd1 _22960_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23630_ _23630_/A vssd1 vssd1 vccd1 vccd1 _25949_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20842_ _21432_/C _21708_/B vssd1 vssd1 vccd1 vccd1 _20844_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_166_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23561_ hold41/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23561_/X sky130_fd_sc_hd__or2b_1
X_20773_ _20772_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20773_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25300_ _25716_/CLK hold310/X vssd1 vssd1 vccd1 vccd1 hold308/A sky130_fd_sc_hd__dfxtp_1
X_22512_ _22512_/A _25893_/Q vssd1 vssd1 vccd1 vccd1 _22512_/Y sky130_fd_sc_hd__nand2_1
X_26280_ _26281_/CLK _26280_/D vssd1 vssd1 vccd1 vccd1 _26280_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_76_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23492_ _24860_/S vssd1 vssd1 vccd1 vccd1 _24944_/S sky130_fd_sc_hd__buf_12
XFILLER_0_135_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25231_ _25687_/CLK hold795/X vssd1 vssd1 vccd1 vccd1 hold794/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22443_ _23008_/B vssd1 vssd1 vccd1 vccd1 _23007_/A sky130_fd_sc_hd__inv_2
XFILLER_0_73_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25162_ _25743_/CLK hold793/X vssd1 vssd1 vccd1 vccd1 hold791/A sky130_fd_sc_hd__dfxtp_1
X_22374_ _22375_/B _22375_/A vssd1 vssd1 vccd1 vccd1 _22376_/A sky130_fd_sc_hd__or2_1
XFILLER_0_115_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24113_ _24113_/A vssd1 vssd1 vccd1 vccd1 _26104_/D sky130_fd_sc_hd__clkbuf_1
X_21325_ _26316_/Q _21228_/X hold587/X vssd1 vssd1 vccd1 vccd1 _21328_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25093_ _26305_/CLK _25093_/D vssd1 vssd1 vccd1 vccd1 _25093_/Q sky130_fd_sc_hd__dfxtp_1
X_24044_ _26082_/Q hold2534/X _24047_/S vssd1 vssd1 vccd1 vccd1 _24044_/X sky130_fd_sc_hd__mux2_1
X_21256_ _26313_/Q hold539/X vssd1 vssd1 vccd1 vccd1 _21256_/Y sky130_fd_sc_hd__nand2_1
Xhold450 hold450/A vssd1 vssd1 vccd1 vccd1 hold450/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 hold461/A vssd1 vssd1 vccd1 vccd1 hold461/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold472 hold472/A vssd1 vssd1 vccd1 vccd1 hold472/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold483 hold483/A vssd1 vssd1 vccd1 vccd1 hold483/X sky130_fd_sc_hd__dlygate4sd3_1
X_20207_ _20207_/A _20207_/B vssd1 vssd1 vccd1 vccd1 _20209_/A sky130_fd_sc_hd__nand2_1
Xhold494 hold494/A vssd1 vssd1 vccd1 vccd1 hold494/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21187_ _25872_/Q _21187_/B _21187_/C vssd1 vssd1 vccd1 vccd1 _21190_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_102_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20138_ _20138_/A _20138_/B vssd1 vssd1 vccd1 vccd1 _20148_/A sky130_fd_sc_hd__nand2_1
X_25995_ _25998_/CLK _25995_/D vssd1 vssd1 vccd1 vccd1 _25995_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_69_clk _25472_/CLK vssd1 vssd1 vccd1 vccd1 _26065_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24946_ _24946_/A _24946_/B vssd1 vssd1 vccd1 vccd1 _24946_/Y sky130_fd_sc_hd__nor2_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ _12930_/X _12958_/X _12917_/X _12959_/X vssd1 vssd1 vccd1 vccd1 _12960_/X
+ sky130_fd_sc_hd__o211a_1
X_20069_ _20069_/A _20069_/B vssd1 vssd1 vccd1 vccd1 _20070_/B sky130_fd_sc_hd__xor2_2
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 _13163_/X vssd1 vssd1 vccd1 vccd1 _25080_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1161 _25549_/Q vssd1 vssd1 vccd1 vccd1 _16771_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1172 _13048_/X vssd1 vssd1 vccd1 vccd1 _25059_/D sky130_fd_sc_hd__dlygate4sd3_1
X_24877_ _24957_/S _24877_/B vssd1 vssd1 vccd1 vccd1 _24877_/X sky130_fd_sc_hd__or2_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1183 _25072_/Q vssd1 vssd1 vccd1 vccd1 _18107_/B sky130_fd_sc_hd__dlygate4sd3_1
X_12891_ _13220_/A vssd1 vssd1 vccd1 vccd1 _12891_/X sky130_fd_sc_hd__clkbuf_16
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 _21127_/Y vssd1 vssd1 vccd1 vccd1 _25805_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _14645_/A hold260/X vssd1 vssd1 vccd1 vccd1 hold261/A sky130_fd_sc_hd__nand2_1
X_23828_ hold2165/X hold1900/X _23831_/S vssd1 vssd1 vccd1 vccd1 _23829_/A sky130_fd_sc_hd__mux2_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _14585_/A hold212/X vssd1 vssd1 vccd1 vccd1 hold213/A sky130_fd_sc_hd__nand2_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23759_ _23759_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23760_/A sky130_fd_sc_hd__and2_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _16298_/X _16299_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _16300_/X sky130_fd_sc_hd__a21o_1
X_13512_ _18122_/B _13518_/B vssd1 vssd1 vccd1 vccd1 _13512_/Y sky130_fd_sc_hd__nor2_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17280_ _17549_/A _17629_/A vssd1 vssd1 vccd1 vccd1 _17281_/B sky130_fd_sc_hd__xnor2_2
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _14525_/A hold296/X vssd1 vssd1 vccd1 vccd1 hold297/A sky130_fd_sc_hd__nand2_1
XFILLER_0_166_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16231_ _16231_/A vssd1 vssd1 vccd1 vccd1 _16473_/A sky130_fd_sc_hd__clkbuf_8
X_25429_ _26001_/CLK _25429_/D vssd1 vssd1 vccd1 vccd1 _25429_/Q sky130_fd_sc_hd__dfxtp_1
X_13443_ _26337_/Q _25706_/Q vssd1 vssd1 vccd1 vccd1 _14678_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_181_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16162_ _16150_/B _16156_/B _16149_/B _16161_/Y vssd1 vssd1 vccd1 vccd1 _16162_/Y
+ sky130_fd_sc_hd__o211ai_1
X_13374_ _26197_/Q _13239_/X _13373_/X vssd1 vssd1 vccd1 vccd1 _13374_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15113_ _16715_/B vssd1 vssd1 vccd1 vccd1 _22453_/B sky130_fd_sc_hd__inv_2
XFILLER_0_180_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16093_ _22322_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _16095_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15044_ _15270_/A _15028_/A _15028_/B vssd1 vssd1 vccd1 vccd1 _15046_/A sky130_fd_sc_hd__a21bo_1
X_19921_ _19920_/Y _19130_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19923_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19852_ _19975_/A _19852_/B vssd1 vssd1 vccd1 vccd1 _19852_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18803_ _18801_/Y _18802_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25684_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19783_ _19781_/Y _19782_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19783_/Y sky130_fd_sc_hd__a21oi_1
X_16995_ _25905_/Q _25904_/Q vssd1 vssd1 vccd1 vccd1 _17683_/B sky130_fd_sc_hd__nor2_1
X_18734_ _18734_/A _18734_/B _18734_/C vssd1 vssd1 vccd1 vccd1 _22438_/A sky130_fd_sc_hd__nand3_2
X_15946_ _16274_/A _16273_/B _15945_/X vssd1 vssd1 vccd1 vccd1 _15953_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_clk _26093_/CLK vssd1 vssd1 vccd1 vccd1 _26130_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_183_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18665_ _22370_/B _25631_/Q vssd1 vssd1 vccd1 vccd1 _18667_/A sky130_fd_sc_hd__nand2_1
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15877_ _15875_/Y hold775/X _15805_/X vssd1 vssd1 vccd1 vccd1 hold776/A sky130_fd_sc_hd__a21oi_1
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17616_ _17616_/A _17616_/B vssd1 vssd1 vccd1 vccd1 _17616_/X sky130_fd_sc_hd__xor2_1
X_14828_ _25852_/Q _12527_/A _15013_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14828_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18596_ _18596_/A _18596_/B vssd1 vssd1 vccd1 vccd1 _18596_/X sky130_fd_sc_hd__xor2_1
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17547_ _17545_/Y _17546_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _17547_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14759_ _14900_/A _14759_/B vssd1 vssd1 vccd1 vccd1 _14759_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17478_ _17478_/A _17478_/B vssd1 vssd1 vccd1 vccd1 _17478_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_129_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19217_ _20506_/A _22160_/B _25595_/Q vssd1 vssd1 vccd1 vccd1 _20511_/C sky130_fd_sc_hd__nand3_1
X_16429_ _16441_/B _16430_/A vssd1 vssd1 vccd1 vccd1 _16429_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19148_ _23199_/A vssd1 vssd1 vccd1 vccd1 _22902_/B sky130_fd_sc_hd__buf_8
XFILLER_0_131_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19079_ _19077_/Y _19078_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25708_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_160_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21110_ _21110_/A _21110_/B vssd1 vssd1 vccd1 vccd1 _21594_/C sky130_fd_sc_hd__nand2_2
X_22090_ _22653_/A _22090_/B vssd1 vssd1 vccd1 vccd1 _22090_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21041_ _21040_/Y _20192_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21041_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24800_ _24800_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24801_/A sky130_fd_sc_hd__and2_1
X_25780_ _26281_/CLK _25780_/D vssd1 vssd1 vccd1 vccd1 _25780_/Q sky130_fd_sc_hd__dfxtp_2
X_22992_ _23138_/A _22992_/B vssd1 vssd1 vccd1 vccd1 _22993_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_179_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24731_ hold1959/X _26306_/Q _24740_/S vssd1 vssd1 vccd1 vccd1 _24731_/X sky130_fd_sc_hd__mux2_1
X_21943_ _21943_/A _21943_/B vssd1 vssd1 vccd1 vccd1 _21944_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_55_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24662_ _24662_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24663_/A sky130_fd_sc_hd__and2_1
XFILLER_0_96_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21874_ _21874_/A _21874_/B vssd1 vssd1 vccd1 vccd1 _21875_/B sky130_fd_sc_hd__nand2_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23613_ hold2023/X _25944_/Q _23677_/S vssd1 vssd1 vccd1 vccd1 _23613_/X sky130_fd_sc_hd__mux2_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20825_ _20824_/B _20825_/B _20825_/C vssd1 vssd1 vccd1 vccd1 _20826_/B sky130_fd_sc_hd__nand3b_1
X_24593_ _24593_/A vssd1 vssd1 vccd1 vccd1 _26260_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26332_ _26334_/CLK _26332_/D vssd1 vssd1 vccd1 vccd1 _26332_/Q sky130_fd_sc_hd__dfxtp_2
X_23544_ hold233/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23544_/X sky130_fd_sc_hd__or2b_1
X_20756_ _20756_/A _22595_/B _20756_/C vssd1 vssd1 vccd1 vccd1 _20759_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_65_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26263_ _26263_/CLK _26263_/D vssd1 vssd1 vccd1 vccd1 _26263_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23475_ hold80/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23475_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20687_ _21368_/C _21644_/B vssd1 vssd1 vccd1 vccd1 _20689_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25214_ _26289_/CLK hold625/X vssd1 vssd1 vccd1 vccd1 hold623/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22426_ _15095_/B _22893_/A _22829_/A vssd1 vssd1 vccd1 vccd1 _22426_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26194_ _26198_/CLK _26194_/D vssd1 vssd1 vccd1 vccd1 _26194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25145_ _25727_/CLK hold562/X vssd1 vssd1 vccd1 vccd1 hold560/A sky130_fd_sc_hd__dfxtp_1
X_22357_ _22791_/B _22941_/B vssd1 vssd1 vccd1 vccd1 _22359_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_66_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21308_ _21308_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21313_/A sky130_fd_sc_hd__nand2_1
X_25076_ _25797_/CLK _25076_/D vssd1 vssd1 vccd1 vccd1 _25076_/Q sky130_fd_sc_hd__dfxtp_1
X_13090_ _26150_/Q _13065_/X _13089_/X vssd1 vssd1 vccd1 vccd1 _13090_/X sky130_fd_sc_hd__a21o_1
X_22288_ _22286_/X _22287_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _22288_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24027_ _24027_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24028_/A sky130_fd_sc_hd__and2_1
XFILLER_0_130_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold280 hold280/A vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
X_21239_ _21241_/B _21241_/C vssd1 vssd1 vccd1 vccd1 _21240_/A sky130_fd_sc_hd__nand2_1
Xhold291 hold291/A vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15800_ _15800_/A _15800_/B vssd1 vssd1 vccd1 vccd1 _15830_/B sky130_fd_sc_hd__nor2_1
X_16780_ _25872_/Q _13468_/X _16774_/Y vssd1 vssd1 vccd1 vccd1 _16780_/Y sky130_fd_sc_hd__a21oi_1
X_13992_ _14061_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13992_/Y sky130_fd_sc_hd__nand2_1
X_25978_ _26041_/CLK _25978_/D vssd1 vssd1 vccd1 vccd1 _25978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15731_ _15731_/A _15731_/B vssd1 vssd1 vccd1 vccd1 _15764_/A sky130_fd_sc_hd__nor2_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ _26122_/Q _12907_/X _12942_/X vssd1 vssd1 vccd1 vccd1 _12943_/X sky130_fd_sc_hd__a21o_1
X_24929_ _24919_/X _24928_/X _24949_/S vssd1 vssd1 vccd1 vccd1 _24930_/A sky130_fd_sc_hd__mux2_2
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ _18450_/A _18450_/B _18450_/C vssd1 vssd1 vccd1 vccd1 _22067_/A sky130_fd_sc_hd__nand3_2
X_15662_ _15662_/A _15692_/A vssd1 vssd1 vccd1 vccd1 _15662_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_158_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ _17343_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12874_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _17578_/A _17629_/B vssd1 vssd1 vccd1 vccd1 _17402_/B sky130_fd_sc_hd__xnor2_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14613_ _14611_/Y hold357/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold358/A sky130_fd_sc_hd__a21oi_1
X_15593_ _15956_/A hold908/X vssd1 vssd1 vccd1 vccd1 _15593_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_29_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18381_ _18381_/A _18381_/B vssd1 vssd1 vccd1 vccd1 _21980_/A sky130_fd_sc_hd__nand2_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14544_ _14542_/Y hold267/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold268/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17332_ _22786_/A vssd1 vssd1 vccd1 vccd1 _17572_/C sky130_fd_sc_hd__buf_8
XFILLER_0_154_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17263_ _19388_/A _17263_/B vssd1 vssd1 vccd1 vccd1 _17542_/A sky130_fd_sc_hd__xor2_4
X_14475_ _14473_/Y hold195/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold196/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19002_ _19000_/Y _19001_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25697_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16214_ _16214_/A _16214_/B vssd1 vssd1 vccd1 vccd1 _16217_/A sky130_fd_sc_hd__nor2_1
X_13426_ _14262_/B vssd1 vssd1 vccd1 vccd1 _13426_/X sky130_fd_sc_hd__buf_12
XFILLER_0_180_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17194_ _19317_/A _17194_/B vssd1 vssd1 vccd1 vccd1 _17506_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_181_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16145_ _16143_/X _16144_/Y _16076_/X vssd1 vssd1 vccd1 vccd1 hold965/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13357_ _18941_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13357_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16076_ _17568_/A vssd1 vssd1 vccd1 vccd1 _16076_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13288_ _13207_/X _13286_/X _13192_/X _13287_/X vssd1 vssd1 vccd1 vccd1 _13288_/X
+ sky130_fd_sc_hd__o211a_1
X_15027_ _15027_/A _15027_/B vssd1 vssd1 vccd1 vccd1 _15028_/B sky130_fd_sc_hd__nand2_1
X_19904_ _19975_/A _19904_/B vssd1 vssd1 vccd1 vccd1 _19904_/Y sky130_fd_sc_hd__nand2_1
Xhold2609 _24621_/X vssd1 vssd1 vccd1 vccd1 _24622_/A sky130_fd_sc_hd__dlygate4sd3_1
X_19835_ _19835_/A _19835_/B vssd1 vssd1 vccd1 vccd1 _19835_/Y sky130_fd_sc_hd__nand2_1
Xhold1908 _23859_/X vssd1 vssd1 vccd1 vccd1 _23860_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1919 _24790_/X vssd1 vssd1 vccd1 vccd1 _24791_/A sky130_fd_sc_hd__dlygate4sd3_1
X_19766_ _22902_/B vssd1 vssd1 vccd1 vccd1 _19766_/X sky130_fd_sc_hd__buf_6
X_16978_ _16976_/Y _16977_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _16978_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput4 io_in[3] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_2
X_18717_ _18919_/A _18996_/A vssd1 vssd1 vccd1 vccd1 _18718_/B sky130_fd_sc_hd__xnor2_1
X_15929_ hold443/X vssd1 vssd1 vccd1 vccd1 _15932_/B sky130_fd_sc_hd__inv_2
XFILLER_0_189_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19697_ _26254_/Q _19483_/X hold515/X vssd1 vssd1 vccd1 vccd1 _19697_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18648_ _18951_/A _18652_/B vssd1 vssd1 vccd1 vccd1 _18650_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_189_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18579_ _18579_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18579_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20610_ _20610_/A _20610_/B _21279_/B vssd1 vssd1 vccd1 vccd1 _20614_/A sky130_fd_sc_hd__nand3_1
X_21590_ _22058_/A _21590_/B vssd1 vssd1 vccd1 vccd1 _21590_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20541_ _20541_/A _20541_/B vssd1 vssd1 vccd1 vccd1 _20543_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_117_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23260_ _23267_/B _23484_/B vssd1 vssd1 vccd1 vccd1 _23261_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_85_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20472_ _20472_/A _22136_/B _20472_/C vssd1 vssd1 vccd1 vccd1 _20475_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_43_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22211_ _19644_/A _22210_/A _22210_/Y vssd1 vssd1 vccd1 vccd1 _22213_/A sky130_fd_sc_hd__o21ai_1
X_23191_ _23191_/A _23191_/B _23191_/C vssd1 vssd1 vccd1 vccd1 _23193_/A sky130_fd_sc_hd__or3_1
XFILLER_0_131_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22142_ _22561_/A _22142_/B vssd1 vssd1 vccd1 vccd1 _22142_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_112_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22073_ _22073_/A _22775_/A vssd1 vssd1 vccd1 vccd1 _22084_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_22_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25901_ _25901_/CLK _25901_/D vssd1 vssd1 vccd1 vccd1 _25901_/Q sky130_fd_sc_hd__dfxtp_1
X_21024_ _21024_/A _25866_/Q vssd1 vssd1 vccd1 vccd1 _21028_/B sky130_fd_sc_hd__nand2_1
X_25832_ _25835_/CLK _25832_/D vssd1 vssd1 vccd1 vccd1 _25832_/Q sky130_fd_sc_hd__dfxtp_2
X_22975_ _23122_/A _22975_/B vssd1 vssd1 vccd1 vccd1 _22976_/B sky130_fd_sc_hd__nand2_1
X_25763_ _25765_/CLK _25763_/D vssd1 vssd1 vccd1 vccd1 _25763_/Q sky130_fd_sc_hd__dfxtp_1
X_24714_ _24714_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24715_/A sky130_fd_sc_hd__and2_1
X_21926_ _21926_/A _21926_/B vssd1 vssd1 vccd1 vccd1 _22977_/A sky130_fd_sc_hd__xor2_4
X_25694_ _26324_/CLK _25694_/D vssd1 vssd1 vccd1 vccd1 _25694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24645_ hold2661/X _26278_/Q _24664_/S vssd1 vssd1 vccd1 vccd1 _24645_/X sky130_fd_sc_hd__mux2_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21857_ _21857_/A _21857_/B vssd1 vssd1 vccd1 vccd1 _22943_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_139_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20808_ _20808_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _20813_/A sky130_fd_sc_hd__nand2_1
X_12590_ _23923_/A _12591_/A vssd1 vssd1 vccd1 vccd1 _12646_/A sky130_fd_sc_hd__or2_1
XFILLER_0_65_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24576_ _24576_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24577_/A sky130_fd_sc_hd__and2_1
X_21788_ _21788_/A _21788_/B _22909_/A vssd1 vssd1 vccd1 vccd1 _21788_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_65_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23527_ hold35/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23527_/X sky130_fd_sc_hd__or2b_1
X_26315_ _26317_/CLK _26315_/D vssd1 vssd1 vccd1 vccd1 _26315_/Q sky130_fd_sc_hd__dfxtp_2
X_20739_ _20737_/Y _20738_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _20739_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14260_ _14260_/A hold425/X vssd1 vssd1 vccd1 vccd1 hold426/A sky130_fd_sc_hd__nand2_1
X_26246_ _26248_/CLK _26246_/D vssd1 vssd1 vccd1 vccd1 _26246_/Q sky130_fd_sc_hd__dfxtp_2
X_23458_ _25912_/Q _24870_/B vssd1 vssd1 vccd1 vccd1 _24959_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_34_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13211_ _26171_/Q _13065_/X _13210_/X vssd1 vssd1 vccd1 vccd1 _13211_/X sky130_fd_sc_hd__a21o_1
X_22409_ _18716_/A _25825_/Q _22407_/Y _22408_/Y vssd1 vssd1 vccd1 vccd1 _22410_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26177_ _26181_/CLK _26177_/D vssd1 vssd1 vccd1 vccd1 _26177_/Q sky130_fd_sc_hd__dfxtp_1
X_14191_ _26328_/Q _13518_/B _14170_/X _14190_/Y vssd1 vssd1 vccd1 vccd1 _14192_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23389_ hold11/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23389_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_104_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25128_ _26335_/CLK _25128_/D vssd1 vssd1 vccd1 vccd1 _25128_/Q sky130_fd_sc_hd__dfxtp_1
X_13142_ _13049_/X _14524_/A _13067_/X _25657_/Q vssd1 vssd1 vccd1 vccd1 _13142_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17950_ _20780_/B _19317_/A vssd1 vssd1 vccd1 vccd1 _17951_/B sky130_fd_sc_hd__nand2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25059_ _26146_/CLK _25059_/D vssd1 vssd1 vccd1 vccd1 _25059_/Q sky130_fd_sc_hd__dfxtp_1
X_13073_ _13049_/X _14485_/A _13067_/X _25644_/Q vssd1 vssd1 vccd1 vccd1 _13073_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16901_ _16899_/Y _16900_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16901_/Y sky130_fd_sc_hd__a21oi_1
X_17881_ _17881_/A _17881_/B vssd1 vssd1 vccd1 vccd1 _17882_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_139_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19620_ _19621_/B _19621_/A vssd1 vssd1 vccd1 vccd1 _19620_/X sky130_fd_sc_hd__or2_1
X_16832_ _16830_/X _16711_/X _16831_/Y _25879_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16833_/A sky130_fd_sc_hd__a32o_1
X_19551_ _19551_/A _19551_/B vssd1 vssd1 vccd1 vccd1 _19551_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_189_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16763_ _16763_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16763_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13975_ _25791_/Q vssd1 vssd1 vccd1 vccd1 _17814_/B sky130_fd_sc_hd__inv_2
X_18502_ _20099_/B _19616_/A vssd1 vssd1 vccd1 vccd1 _18503_/B sky130_fd_sc_hd__nand2_1
X_15714_ _15701_/A _15691_/B _15689_/A vssd1 vssd1 vccd1 vccd1 _15716_/A sky130_fd_sc_hd__a21o_1
X_12926_ _12891_/X _14394_/A _12909_/X _25616_/Q vssd1 vssd1 vccd1 vccd1 _12926_/X
+ sky130_fd_sc_hd__a22o_1
X_19482_ _19480_/Y _19481_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19482_/Y sky130_fd_sc_hd__a21oi_1
X_16694_ _16694_/A _16694_/B vssd1 vssd1 vccd1 vccd1 _16696_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_158_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18433_ _18637_/A _18778_/A vssd1 vssd1 vccd1 vccd1 _18434_/B sky130_fd_sc_hd__xnor2_1
X_15645_ _15645_/A _15645_/B vssd1 vssd1 vccd1 vccd1 _15645_/Y sky130_fd_sc_hd__nand2_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12857_ _12726_/B _14355_/A _12752_/X _25603_/Q vssd1 vssd1 vccd1 vccd1 _12857_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18364_ _18446_/A _25744_/Q _21716_/A vssd1 vssd1 vccd1 vccd1 _18365_/C sky130_fd_sc_hd__nand3_1
X_15576_ _15574_/X hold2473/X _15464_/X vssd1 vssd1 vccd1 vccd1 _15576_/Y sky130_fd_sc_hd__a21oi_1
X_12788_ _26221_/Q _25590_/Q vssd1 vssd1 vccd1 vccd1 _14313_/A sky130_fd_sc_hd__xor2_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17315_ _21048_/B _25867_/Q _21072_/B vssd1 vssd1 vccd1 vccd1 _17316_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14527_ _14524_/Y hold132/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold133/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18295_ _18295_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18295_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17246_ _17272_/A _17246_/B vssd1 vssd1 vccd1 vccd1 _17246_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_189_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14458_ _14458_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14458_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_52_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13409_ _13220_/A _14660_/A _13242_/X _19802_/A vssd1 vssd1 vccd1 vccd1 _13409_/X
+ sky130_fd_sc_hd__a22o_1
X_17177_ _17272_/A _17177_/B vssd1 vssd1 vccd1 vccd1 _17177_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14389_ _14404_/A hold251/X vssd1 vssd1 vccd1 vccd1 hold252/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16128_ _16126_/X _16127_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _16128_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16059_ _16273_/C _15945_/X _16056_/X _16058_/X vssd1 vssd1 vccd1 vccd1 _16059_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_110_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2406 _25446_/Q vssd1 vssd1 vccd1 vccd1 _15296_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2417 _25676_/Q vssd1 vssd1 vccd1 vccd1 _13259_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2428 _12574_/Y vssd1 vssd1 vccd1 vccd1 _12576_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2439 _25646_/Q vssd1 vssd1 vccd1 vccd1 _13082_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1705 _25650_/Q vssd1 vssd1 vccd1 vccd1 _18011_/B sky130_fd_sc_hd__dlygate4sd3_1
X_19818_ _20634_/A _19816_/Y _20639_/C vssd1 vssd1 vccd1 vccd1 _19901_/B sky130_fd_sc_hd__o21a_2
Xhold1716 _20854_/Y vssd1 vssd1 vccd1 vccd1 _25795_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1727 hold2756/X vssd1 vssd1 vccd1 vccd1 _18232_/B sky130_fd_sc_hd__buf_2
Xhold1738 _25593_/Q vssd1 vssd1 vccd1 vccd1 _17177_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1749 hold2757/X vssd1 vssd1 vccd1 vccd1 _17064_/B sky130_fd_sc_hd__clkbuf_2
X_19749_ _19749_/A _19749_/B vssd1 vssd1 vccd1 vccd1 _19749_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_155_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22760_ _22760_/A _22760_/B vssd1 vssd1 vccd1 vccd1 _22761_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_67_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21711_ _21711_/A _21711_/B vssd1 vssd1 vccd1 vccd1 _21712_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_149_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22691_ _22691_/A _25900_/Q vssd1 vssd1 vccd1 vccd1 _22691_/Y sky130_fd_sc_hd__nand2_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24430_ hold2089/X hold1988/X _24433_/S vssd1 vssd1 vccd1 vccd1 _24431_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_177_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21642_ _21644_/B _21693_/B vssd1 vssd1 vccd1 vccd1 _21643_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24361_ _24361_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24362_/A sky130_fd_sc_hd__and2_1
X_21573_ _21573_/A _21573_/B vssd1 vssd1 vccd1 vccd1 _21573_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_20 _17308_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_31 _19038_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26100_ _26103_/CLK _26100_/D vssd1 vssd1 vccd1 vccd1 _26100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23312_ _23312_/A vssd1 vssd1 vccd1 vccd1 _25924_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_42 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20524_ _20526_/B vssd1 vssd1 vccd1 vccd1 _20525_/B sky130_fd_sc_hd__inv_2
XFILLER_0_90_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24292_ _24292_/A vssd1 vssd1 vccd1 vccd1 _26162_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_64 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_75 _25837_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26031_ _26032_/CLK _26031_/D vssd1 vssd1 vccd1 vccd1 _26031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23243_ _23243_/A vssd1 vssd1 vccd1 vccd1 _23244_/B sky130_fd_sc_hd__inv_2
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20455_ _20455_/A _21172_/B _20455_/C vssd1 vssd1 vccd1 vccd1 _20456_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_15_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23174_ _26083_/Q vssd1 vssd1 vccd1 vccd1 _23175_/A sky130_fd_sc_hd__inv_2
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20386_ _20386_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _20386_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_179_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22125_ _22125_/A _22821_/B vssd1 vssd1 vccd1 vccd1 _22126_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22056_ _22054_/X _22055_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _22056_/Y sky130_fd_sc_hd__a21oi_2
X_21007_ _21007_/A _21007_/B _21007_/C vssd1 vssd1 vccd1 vccd1 _21011_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_103_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25815_ _25822_/CLK _25815_/D vssd1 vssd1 vccd1 vccd1 _25815_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13760_ _13760_/A hold671/X vssd1 vssd1 vccd1 vccd1 hold672/A sky130_fd_sc_hd__nand2_1
XFILLER_0_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22958_ _23106_/A _22958_/B vssd1 vssd1 vccd1 vccd1 _22959_/B sky130_fd_sc_hd__nand2_1
X_25746_ _25748_/CLK _25746_/D vssd1 vssd1 vccd1 vccd1 _25746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12711_ _12711_/A _24983_/Q _24982_/Q _12711_/D vssd1 vssd1 vccd1 vccd1 _12712_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_35_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21909_ _21909_/A _21909_/B vssd1 vssd1 vccd1 vccd1 _21910_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_179_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13691_ _13703_/A _13691_/B vssd1 vssd1 vccd1 vccd1 _13691_/Y sky130_fd_sc_hd__nand2_1
X_22889_ _22887_/X _22888_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _22889_/Y sky130_fd_sc_hd__a21oi_1
X_25677_ _26306_/CLK _25677_/D vssd1 vssd1 vccd1 vccd1 _25677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15430_ _15430_/A _15443_/B vssd1 vssd1 vccd1 vccd1 _15430_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_168_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12642_ _24976_/Q _24977_/Q vssd1 vssd1 vccd1 vccd1 _12645_/C sky130_fd_sc_hd__nand2_1
X_24628_ _24628_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24629_/A sky130_fd_sc_hd__and2_1
XFILLER_0_66_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15361_ _15361_/A _15361_/B vssd1 vssd1 vccd1 vccd1 _15361_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_26_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12573_ _12575_/B vssd1 vssd1 vccd1 vccd1 _23596_/B sky130_fd_sc_hd__inv_2
XFILLER_0_136_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24559_ hold2567/X _26250_/Q _24587_/S vssd1 vssd1 vccd1 vccd1 _24559_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17100_ _25652_/Q _17100_/B vssd1 vssd1 vccd1 vccd1 _17652_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_108_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14312_ _14310_/Y hold141/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold142/A sky130_fd_sc_hd__a21oi_1
X_15292_ _15827_/A _15265_/A _15264_/B vssd1 vssd1 vccd1 vccd1 _15294_/A sky130_fd_sc_hd__a21o_1
X_18080_ _18080_/A _18080_/B vssd1 vssd1 vccd1 vccd1 _22247_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_136_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14243_ _25834_/Q vssd1 vssd1 vccd1 vccd1 _18895_/B sky130_fd_sc_hd__inv_2
X_17031_ _17031_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17031_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_184_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26229_ _26232_/CLK _26229_/D vssd1 vssd1 vccd1 vccd1 _26229_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_80_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14174_ _14180_/A _14174_/B vssd1 vssd1 vccd1 vccd1 _14174_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_180_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13125_ _26285_/Q _25654_/Q vssd1 vssd1 vccd1 vccd1 _14515_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18982_ _19032_/A _18982_/B vssd1 vssd1 vccd1 vccd1 _18982_/X sky130_fd_sc_hd__xor2_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ _17933_/A _19137_/A vssd1 vssd1 vccd1 vccd1 _17934_/A sky130_fd_sc_hd__xor2_2
X_13056_ _13049_/X _14476_/A _12909_/X _25641_/Q vssd1 vssd1 vccd1 vccd1 _13056_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17864_ _18535_/A _17864_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _17864_/X sky130_fd_sc_hd__and3_1
XFILLER_0_79_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19603_ _20054_/A _22120_/B _25622_/Q vssd1 vssd1 vccd1 vccd1 _20058_/C sky130_fd_sc_hd__nand3_1
X_16815_ _16935_/A _16820_/B vssd1 vssd1 vccd1 vccd1 _16817_/B sky130_fd_sc_hd__nand2_1
X_17795_ _18612_/A _25720_/Q _18083_/C vssd1 vssd1 vccd1 vccd1 _17796_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_88_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19534_ _21210_/A _19532_/Y _21214_/C vssd1 vssd1 vccd1 vccd1 _19621_/B sky130_fd_sc_hd__o21a_2
X_16746_ _16747_/B _16747_/A vssd1 vssd1 vccd1 vccd1 _16746_/X sky130_fd_sc_hd__or2_1
X_13958_ _17990_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13958_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_152_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19465_ _19457_/X _19464_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19465_/Y sky130_fd_sc_hd__o21ai_1
X_12909_ _13242_/A vssd1 vssd1 vccd1 vccd1 _12909_/X sky130_fd_sc_hd__buf_12
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16677_ _16678_/B _16678_/A vssd1 vssd1 vccd1 vccd1 _16695_/B sky130_fd_sc_hd__or2_1
XFILLER_0_5_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13889_ _25777_/Q vssd1 vssd1 vccd1 vccd1 _17931_/B sky130_fd_sc_hd__inv_2
XFILLER_0_69_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18416_ _18413_/X _18269_/X _18415_/X vssd1 vssd1 vccd1 vccd1 _18417_/A sky130_fd_sc_hd__a21o_1
X_15628_ _15615_/X _15693_/B _15627_/Y vssd1 vssd1 vccd1 vccd1 _15628_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19396_ _19452_/A _19396_/B vssd1 vssd1 vccd1 vccd1 _19396_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_5_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18347_ _18952_/A _18347_/B _18952_/C vssd1 vssd1 vccd1 vccd1 _18348_/C sky130_fd_sc_hd__nand3_1
X_15559_ _15577_/B _15560_/A vssd1 vssd1 vccd1 vccd1 _15559_/X sky130_fd_sc_hd__or2_1
XFILLER_0_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18278_ _21075_/B _19458_/A vssd1 vssd1 vccd1 vccd1 _18279_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_142_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17229_ _17229_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17229_/Y sky130_fd_sc_hd__nand2_1
Xhold802 hold802/A vssd1 vssd1 vccd1 vccd1 hold802/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold813 hold813/A vssd1 vssd1 vccd1 vccd1 hold813/X sky130_fd_sc_hd__dlygate4sd3_1
X_20240_ _20240_/A _22272_/B _20240_/C vssd1 vssd1 vccd1 vccd1 _20244_/C sky130_fd_sc_hd__nand3_1
Xhold824 hold824/A vssd1 vssd1 vccd1 vccd1 hold824/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold835 hold835/A vssd1 vssd1 vccd1 vccd1 hold835/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 hold846/A vssd1 vssd1 vccd1 vccd1 hold846/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold857 hold857/A vssd1 vssd1 vccd1 vccd1 hold857/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold868 hold868/A vssd1 vssd1 vccd1 vccd1 hold868/X sky130_fd_sc_hd__dlygate4sd3_1
X_20171_ _20171_/A _20171_/B _20171_/C vssd1 vssd1 vccd1 vccd1 _20172_/B sky130_fd_sc_hd__nand3_1
Xhold879 hold879/A vssd1 vssd1 vccd1 vccd1 hold879/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2203 _25417_/Q vssd1 vssd1 vccd1 vccd1 _14938_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2214 _26205_/Q vssd1 vssd1 vccd1 vccd1 hold2214/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2225 _23668_/X vssd1 vssd1 vccd1 vccd1 _23669_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2236 _24261_/X vssd1 vssd1 vccd1 vccd1 _24262_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2247 _14993_/Y vssd1 vssd1 vccd1 vccd1 hold2247/X sky130_fd_sc_hd__dlygate4sd3_1
X_23930_ _23930_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23931_/A sky130_fd_sc_hd__and2_1
Xhold1502 _23038_/Y vssd1 vssd1 vccd1 vccd1 _25891_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2258 _25942_/Q vssd1 vssd1 vccd1 vccd1 hold2258/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1513 _25559_/Q vssd1 vssd1 vccd1 vccd1 _16837_/B sky130_fd_sc_hd__buf_1
Xhold1524 _23182_/Y vssd1 vssd1 vccd1 vccd1 _25900_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2269 _26192_/Q vssd1 vssd1 vccd1 vccd1 hold2269/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1535 _25808_/Q vssd1 vssd1 vccd1 vccd1 _21208_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23861_ _23861_/A vssd1 vssd1 vccd1 vccd1 _26024_/D sky130_fd_sc_hd__clkbuf_1
Xhold1546 _13382_/X vssd1 vssd1 vccd1 vccd1 _25115_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1557 _25758_/Q vssd1 vssd1 vccd1 vccd1 _19810_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1568 _25780_/Q vssd1 vssd1 vccd1 vccd1 _20270_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1579 _22989_/Y vssd1 vssd1 vccd1 vccd1 _25888_/D sky130_fd_sc_hd__dlygate4sd3_1
X_22812_ _23188_/A _22812_/B vssd1 vssd1 vccd1 vccd1 _22812_/X sky130_fd_sc_hd__or2_1
X_25600_ _26109_/CLK _25600_/D vssd1 vssd1 vccd1 vccd1 _25600_/Q sky130_fd_sc_hd__dfxtp_4
X_23792_ _23792_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23793_/A sky130_fd_sc_hd__and2_1
XFILLER_0_149_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25531_ _25534_/CLK hold963/X vssd1 vssd1 vccd1 vccd1 hold962/A sky130_fd_sc_hd__dfxtp_1
X_22743_ _22743_/A _23056_/B vssd1 vssd1 vccd1 vccd1 _22744_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25462_ _26012_/CLK hold909/X vssd1 vssd1 vccd1 vccd1 hold908/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22674_ _23007_/A _23152_/B vssd1 vssd1 vccd1 vccd1 _22675_/B sky130_fd_sc_hd__nand2_1
Xascon_wrapper_15 vssd1 vssd1 vccd1 vccd1 io_oeb[1] ascon_wrapper_15/LO sky130_fd_sc_hd__conb_1
XFILLER_0_165_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24413_ _24413_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24414_/A sky130_fd_sc_hd__and2_1
XFILLER_0_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21625_ _21676_/B _21629_/B vssd1 vssd1 vccd1 vccd1 _21627_/A sky130_fd_sc_hd__nand2_1
X_25393_ _25999_/CLK _25393_/D vssd1 vssd1 vccd1 vccd1 _25393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24344_ hold2332/X hold2334/X _24356_/S vssd1 vssd1 vccd1 vccd1 _24345_/A sky130_fd_sc_hd__mux2_1
X_21556_ _21556_/A _22902_/B vssd1 vssd1 vccd1 vccd1 _21556_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20507_ _20507_/A _20507_/B vssd1 vssd1 vccd1 vccd1 _20511_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24275_ _24275_/A vssd1 vssd1 vccd1 vccd1 _26157_/D sky130_fd_sc_hd__clkbuf_1
X_21487_ _26326_/Q hold698/X vssd1 vssd1 vccd1 vccd1 _21487_/Y sky130_fd_sc_hd__nand2_1
X_26014_ _26014_/CLK _26014_/D vssd1 vssd1 vccd1 vccd1 _26014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23226_ _24858_/S vssd1 vssd1 vccd1 vccd1 _24946_/A sky130_fd_sc_hd__inv_16
X_20438_ _20438_/A _22391_/B vssd1 vssd1 vccd1 vccd1 _20439_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23157_ _15775_/B _22893_/A _22829_/A vssd1 vssd1 vccd1 vccd1 _23157_/Y sky130_fd_sc_hd__a21oi_1
X_20369_ _20369_/A _20369_/B vssd1 vssd1 vccd1 vccd1 _20371_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_105_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22108_ _22108_/A _22108_/B vssd1 vssd1 vccd1 vccd1 _23074_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_100_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23088_ _23088_/A _23088_/B vssd1 vssd1 vccd1 vccd1 _23089_/B sky130_fd_sc_hd__nand2_1
X_14930_ _25416_/Q _14931_/A vssd1 vssd1 vccd1 vccd1 _14932_/A sky130_fd_sc_hd__or2_1
X_22039_ _22039_/A _25875_/Q vssd1 vssd1 vccd1 vccd1 _22039_/Y sky130_fd_sc_hd__nand2_1
X_14861_ _22292_/B _15543_/B vssd1 vssd1 vccd1 vccd1 _14862_/A sky130_fd_sc_hd__nand2_1
X_16600_ _16574_/A _16596_/B _16577_/Y _16597_/B _16588_/A vssd1 vssd1 vccd1 vccd1
+ _16600_/X sky130_fd_sc_hd__a221o_1
X_13812_ _13807_/Y _13811_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold945/A sky130_fd_sc_hd__a21oi_1
X_17580_ _17624_/A _17580_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _17580_/X sky130_fd_sc_hd__and3_1
XFILLER_0_187_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14792_ _25848_/Q _12527_/A _14980_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14792_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16531_ _16529_/Y _16530_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 hold865/A sky130_fd_sc_hd__a21oi_1
X_25729_ _25729_/CLK _25729_/D vssd1 vssd1 vccd1 vccd1 _25729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13743_ _25754_/Q vssd1 vssd1 vccd1 vccd1 _18571_/B sky130_fd_sc_hd__inv_2
XFILLER_0_168_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19250_ _19249_/Y _21228_/A _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _19252_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16462_ _16462_/A _16487_/A vssd1 vssd1 vccd1 vccd1 _16468_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13674_ _13760_/A hold545/X vssd1 vssd1 vccd1 vccd1 hold546/A sky130_fd_sc_hd__nand2_1
XFILLER_0_168_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18201_ _18611_/A _25736_/Q vssd1 vssd1 vccd1 vccd1 _18203_/A sky130_fd_sc_hd__nand2_1
X_15413_ _15443_/A _15414_/A vssd1 vssd1 vccd1 vccd1 _15413_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12625_ _12628_/A _24836_/B _12625_/C vssd1 vssd1 vccd1 vccd1 _12626_/A sky130_fd_sc_hd__and3_1
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19181_ _19989_/A _19261_/A vssd1 vssd1 vccd1 vccd1 _19183_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_66_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16393_ _16393_/A _16393_/B vssd1 vssd1 vccd1 vccd1 _16394_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18132_ _18132_/A _18132_/B vssd1 vssd1 vccd1 vccd1 _21903_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_183_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15344_ _15331_/X _15406_/B _15343_/Y vssd1 vssd1 vccd1 vccd1 _15344_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12556_ _14267_/A _17688_/B _16996_/C _23201_/B vssd1 vssd1 vccd1 vccd1 _12556_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18063_ _20248_/B _25652_/Q vssd1 vssd1 vccd1 vccd1 _18067_/A sky130_fd_sc_hd__nand2_1
X_15275_ _15275_/A _15275_/B vssd1 vssd1 vccd1 vccd1 _15275_/Y sky130_fd_sc_hd__nand2_1
X_12487_ _14893_/A vssd1 vssd1 vccd1 vccd1 _15839_/A sky130_fd_sc_hd__buf_8
XFILLER_0_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17014_ _22586_/A vssd1 vssd1 vccd1 vccd1 _19199_/A sky130_fd_sc_hd__buf_12
Xhold109 hold109/A vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
X_14226_ _18834_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14226_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_111_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14157_ _14236_/A hold647/X vssd1 vssd1 vccd1 vccd1 hold648/A sky130_fd_sc_hd__nand2_1
XFILLER_0_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13108_ _13018_/X _13106_/X _13096_/X _13107_/X vssd1 vssd1 vccd1 vccd1 _13108_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14088_ _14118_/A hold569/X vssd1 vssd1 vccd1 vccd1 hold570/A sky130_fd_sc_hd__nand2_1
X_18965_ _18963_/Y _18964_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25692_/D sky130_fd_sc_hd__a21oi_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17916_ _17916_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _17916_/Y sky130_fd_sc_hd__nand2_1
X_13039_ _26269_/Q _25638_/Q vssd1 vssd1 vccd1 vccd1 _14464_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18896_ _20835_/B _22642_/A vssd1 vssd1 vccd1 vccd1 _20828_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17847_ _17847_/A _17847_/B _17847_/C vssd1 vssd1 vccd1 vccd1 _22310_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_179_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17778_ _17779_/B _17779_/A vssd1 vssd1 vccd1 vccd1 _17780_/A sky130_fd_sc_hd__or2_1
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19517_ _19514_/Y _19517_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19517_/X sky130_fd_sc_hd__and3b_1
X_16729_ _16858_/A _16729_/B vssd1 vssd1 vccd1 vccd1 _16729_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_159_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19448_ _19449_/B _19449_/A vssd1 vssd1 vccd1 vccd1 _19448_/X sky130_fd_sc_hd__or2_1
XFILLER_0_159_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19379_ _19377_/X _19378_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19379_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21410_ _21410_/A _21410_/B vssd1 vssd1 vccd1 vccd1 _21411_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_174_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22390_ _22390_/A _25888_/Q vssd1 vssd1 vccd1 vccd1 _22390_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21341_ _26317_/Q _21228_/X hold821/X vssd1 vssd1 vccd1 vccd1 _21344_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24060_ _24060_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24061_/A sky130_fd_sc_hd__and2_1
Xhold610 hold610/A vssd1 vssd1 vccd1 vccd1 hold610/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21272_ _21272_/A _21272_/B vssd1 vssd1 vccd1 vccd1 _21691_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_64_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold621 hold621/A vssd1 vssd1 vccd1 vccd1 hold621/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23011_ _23011_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _23011_/Y sky130_fd_sc_hd__nand2_1
Xhold632 hold632/A vssd1 vssd1 vccd1 vccd1 hold632/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_25_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold643 hold643/A vssd1 vssd1 vccd1 vccd1 hold643/X sky130_fd_sc_hd__dlygate4sd3_1
X_20223_ _20223_/A _21007_/C vssd1 vssd1 vccd1 vccd1 _20225_/A sky130_fd_sc_hd__nand2_1
Xhold654 hold654/A vssd1 vssd1 vccd1 vccd1 hold654/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold665 hold665/A vssd1 vssd1 vccd1 vccd1 hold665/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold676 hold676/A vssd1 vssd1 vccd1 vccd1 hold676/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 hold687/A vssd1 vssd1 vccd1 vccd1 hold687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 hold698/A vssd1 vssd1 vccd1 vccd1 hold698/X sky130_fd_sc_hd__dlygate4sd3_1
X_20154_ _26280_/Q _20078_/X hold851/X vssd1 vssd1 vccd1 vccd1 _20157_/B sky130_fd_sc_hd__a21oi_1
Xhold2000 _24520_/X vssd1 vssd1 vccd1 vccd1 _24521_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2011 _12707_/Y vssd1 vssd1 vccd1 vccd1 _12715_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2022 _23339_/X vssd1 vssd1 vccd1 vccd1 _23340_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2033 _23822_/X vssd1 vssd1 vccd1 vccd1 _23823_/A sky130_fd_sc_hd__dlygate4sd3_1
X_24962_ _23593_/X _24910_/X hold1981/X vssd1 vssd1 vccd1 vccd1 _24962_/Y sky130_fd_sc_hd__a21boi_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2044 _23868_/X vssd1 vssd1 vccd1 vccd1 _23869_/A sky130_fd_sc_hd__dlygate4sd3_1
X_20085_ _20660_/A _20085_/B vssd1 vssd1 vccd1 vccd1 _20085_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2055 _25933_/Q vssd1 vssd1 vccd1 vccd1 _23351_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1310 _25392_/Q vssd1 vssd1 vccd1 vccd1 _14731_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1321 _16905_/X vssd1 vssd1 vccd1 vccd1 _16906_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2066 _14936_/Y vssd1 vssd1 vccd1 vccd1 _25416_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1332 _16971_/Y vssd1 vssd1 vccd1 vccd1 _25578_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23913_ _23913_/A vssd1 vssd1 vccd1 vccd1 _26041_/D sky130_fd_sc_hd__clkbuf_1
Xhold2077 _26164_/Q vssd1 vssd1 vccd1 vccd1 hold2077/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2088 _23767_/X vssd1 vssd1 vccd1 vccd1 _23768_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1343 _25393_/Q vssd1 vssd1 vccd1 vccd1 _14740_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24893_ _15690_/B _15712_/B _24945_/S vssd1 vssd1 vccd1 vccd1 _24893_/X sky130_fd_sc_hd__mux2_1
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1354 _19753_/Y vssd1 vssd1 vccd1 vccd1 _25754_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2099 _23366_/Y vssd1 vssd1 vccd1 vccd1 _23367_/C sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1365 _25409_/Q vssd1 vssd1 vccd1 vccd1 _14882_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_174_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1376 _20234_/Y vssd1 vssd1 vccd1 vccd1 _25779_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23844_ hold2051/X _26019_/Q _23907_/S vssd1 vssd1 vccd1 vccd1 _23844_/X sky130_fd_sc_hd__mux2_1
Xhold1387 _25566_/Q vssd1 vssd1 vccd1 vccd1 _16886_/B sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1398 _20042_/Y vssd1 vssd1 vccd1 vccd1 _25774_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23775_ _23775_/A vssd1 vssd1 vccd1 vccd1 _25996_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20987_ _20985_/Y _20192_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _20987_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_68_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25514_ _25515_/CLK hold951/X vssd1 vssd1 vccd1 vccd1 hold950/A sky130_fd_sc_hd__dfxtp_1
X_22726_ _23183_/B _23040_/B vssd1 vssd1 vccd1 vccd1 _22728_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25445_ _26052_/CLK _25445_/D vssd1 vssd1 vccd1 vccd1 _25445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22657_ _22656_/A _22454_/X _22656_/B vssd1 vssd1 vccd1 vccd1 _22658_/C sky130_fd_sc_hd__o21ai_1
X_21608_ _21660_/B _21612_/A vssd1 vssd1 vccd1 vccd1 _21610_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_168_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13390_ _26328_/Q _19758_/A vssd1 vssd1 vccd1 vccd1 _14651_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_106_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22588_ _22585_/X _22587_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22588_/Y sky130_fd_sc_hd__a21oi_1
X_25376_ _26202_/CLK hold175/X vssd1 vssd1 vccd1 vccd1 hold173/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21539_ _21539_/A _21539_/B vssd1 vssd1 vccd1 vccd1 _21540_/A sky130_fd_sc_hd__nand2_1
X_24327_ _24327_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24328_/A sky130_fd_sc_hd__and2_1
XFILLER_0_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15060_ _15055_/A _15050_/A _15050_/B vssd1 vssd1 vccd1 vccd1 _15062_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_133_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24258_ hold1995/X _26152_/Q _24279_/S vssd1 vssd1 vccd1 vccd1 _24258_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14011_ _26299_/Q _13988_/X _13981_/X _14010_/Y vssd1 vssd1 vccd1 vccd1 _14012_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23209_ _23211_/B _23212_/A _23209_/C vssd1 vssd1 vccd1 vccd1 _23210_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_120_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24189_ _24189_/A vssd1 vssd1 vccd1 vccd1 _26129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18750_ _18793_/A _25763_/Q _18891_/C vssd1 vssd1 vccd1 vccd1 _18751_/C sky130_fd_sc_hd__nand3_1
X_15962_ _16000_/A _15963_/A vssd1 vssd1 vccd1 vccd1 _15962_/X sky130_fd_sc_hd__or2_1
X_17701_ _25904_/Q _25903_/Q vssd1 vssd1 vccd1 vccd1 _17752_/B sky130_fd_sc_hd__xnor2_2
X_14913_ _14913_/A _14913_/B vssd1 vssd1 vccd1 vccd1 _14925_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_175_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18681_ _18681_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18681_/Y sky130_fd_sc_hd__nand2_1
X_15893_ _15921_/B vssd1 vssd1 vccd1 vccd1 _15900_/B sky130_fd_sc_hd__inv_2
XFILLER_0_37_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17632_ _18535_/A _17632_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _17632_/X sky130_fd_sc_hd__and3_1
X_14844_ _14844_/A _22233_/A vssd1 vssd1 vccd1 vccd1 _22232_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17563_ _17563_/A _17563_/B vssd1 vssd1 vccd1 vccd1 _17563_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_81_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14775_ _25846_/Q _13466_/A _14774_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14776_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19302_ _19299_/Y _19302_/B _19980_/B vssd1 vssd1 vccd1 vccd1 _19302_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_58_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16514_ _16524_/B _16515_/A vssd1 vssd1 vccd1 vccd1 _16514_/X sky130_fd_sc_hd__or2_1
X_13726_ _18509_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13726_/Y sky130_fd_sc_hd__nor2_1
X_17494_ _17492_/X _17241_/X _17493_/X vssd1 vssd1 vccd1 vccd1 _17495_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_39_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19233_ _19248_/A _19322_/B vssd1 vssd1 vccd1 vccd1 _19234_/B sky130_fd_sc_hd__xor2_1
X_16445_ _16461_/A _16462_/A vssd1 vssd1 vccd1 vccd1 _16447_/A sky130_fd_sc_hd__or2_1
XFILLER_0_184_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13657_ _25740_/Q vssd1 vssd1 vccd1 vccd1 _18287_/B sky130_fd_sc_hd__inv_2
XFILLER_0_128_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12608_ _23245_/A vssd1 vssd1 vccd1 vccd1 _12702_/A sky130_fd_sc_hd__buf_12
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19164_ _20349_/A _18185_/B _20354_/C vssd1 vssd1 vccd1 vccd1 _19248_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_54_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _16473_/A hold914/X vssd1 vssd1 vccd1 vccd1 _16376_/Y sky130_fd_sc_hd__nand2_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13588_ _17908_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13588_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_53_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18115_ _25589_/Q _21992_/A vssd1 vssd1 vccd1 vccd1 _18117_/B sky130_fd_sc_hd__nor2_1
X_15327_ _15327_/A _15327_/B vssd1 vssd1 vccd1 vccd1 _15328_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12539_ hold6/X vssd1 vssd1 vccd1 vccd1 _12548_/C sky130_fd_sc_hd__inv_2
X_19095_ _20068_/A vssd1 vssd1 vccd1 vccd1 _19095_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_30_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18046_ _18446_/A _25732_/Q _21716_/A vssd1 vssd1 vccd1 vccd1 _18047_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_83_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15258_ _22653_/B _15812_/B vssd1 vssd1 vccd1 vccd1 _16282_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_112_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14209_ _26331_/Q _13518_/B _14170_/X _14208_/Y vssd1 vssd1 vccd1 vccd1 _14210_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15189_ _16743_/B vssd1 vssd1 vccd1 vccd1 _22555_/B sky130_fd_sc_hd__inv_2
X_19997_ _20660_/A _19997_/B vssd1 vssd1 vccd1 vccd1 _19997_/Y sky130_fd_sc_hd__nand2_1
X_18948_ _25645_/Q _22718_/B vssd1 vssd1 vccd1 vccd1 _18949_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_94_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18879_ _22704_/A vssd1 vssd1 vccd1 vccd1 _18879_/X sky130_fd_sc_hd__buf_12
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20910_ _20913_/A _20913_/C vssd1 vssd1 vccd1 vccd1 _20911_/A sky130_fd_sc_hd__nand2_1
X_21890_ _17976_/B _17080_/B _17977_/B vssd1 vssd1 vccd1 vccd1 _21891_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_96_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20841_ _20841_/A _20841_/B _21384_/C vssd1 vssd1 vccd1 vccd1 _20845_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_162_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23560_ _23557_/Y _23559_/Y _24957_/S vssd1 vssd1 vccd1 vccd1 _23560_/X sky130_fd_sc_hd__mux2_1
X_20772_ _26296_/Q hold656/X vssd1 vssd1 vccd1 vccd1 _20772_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_175_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22511_ _22509_/X _22510_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22511_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23491_ _24940_/S hold65/A _23490_/X vssd1 vssd1 vccd1 vccd1 _23491_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22442_ _22442_/A _22442_/B vssd1 vssd1 vccd1 vccd1 _23008_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_29_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25230_ _25687_/CLK hold541/X vssd1 vssd1 vccd1 vccd1 hold539/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25161_ _25743_/CLK hold676/X vssd1 vssd1 vccd1 vccd1 hold674/A sky130_fd_sc_hd__dfxtp_1
X_22373_ _19729_/A _22372_/A _22372_/Y vssd1 vssd1 vccd1 vccd1 _22375_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_115_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24112_ _24112_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24113_/A sky130_fd_sc_hd__and2_1
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21324_ _21324_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21329_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_128_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25092_ _26175_/CLK _25092_/D vssd1 vssd1 vccd1 vccd1 _25092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24043_ _24043_/A vssd1 vssd1 vccd1 vccd1 _26082_/D sky130_fd_sc_hd__clkbuf_1
X_21255_ _26313_/Q _21228_/X hold539/X vssd1 vssd1 vccd1 vccd1 _21258_/B sky130_fd_sc_hd__a21oi_1
Xhold440 hold440/A vssd1 vssd1 vccd1 vccd1 hold440/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 hold451/A vssd1 vssd1 vccd1 vccd1 hold451/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 hold462/A vssd1 vssd1 vccd1 vccd1 hold462/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 hold473/A vssd1 vssd1 vccd1 vccd1 hold473/X sky130_fd_sc_hd__dlygate4sd3_1
X_20206_ _20208_/B vssd1 vssd1 vccd1 vccd1 _20207_/B sky130_fd_sc_hd__inv_2
XFILLER_0_99_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold484 hold484/A vssd1 vssd1 vccd1 vccd1 hold484/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 hold495/A vssd1 vssd1 vccd1 vccd1 hold495/X sky130_fd_sc_hd__dlygate4sd3_1
X_21186_ _21186_/A _25872_/Q vssd1 vssd1 vccd1 vccd1 _21190_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_187_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20137_ _20139_/C vssd1 vssd1 vccd1 vccd1 _20138_/B sky130_fd_sc_hd__inv_2
XFILLER_0_110_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25994_ _25998_/CLK _25994_/D vssd1 vssd1 vccd1 vccd1 _25994_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24945_ hold958/A hold873/A _24945_/S vssd1 vssd1 vccd1 vccd1 _24946_/B sky130_fd_sc_hd__mux2_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20068_ _20068_/A _20068_/B vssd1 vssd1 vccd1 vccd1 _20069_/B sky130_fd_sc_hd__nand2_1
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 _12890_/X vssd1 vssd1 vccd1 vccd1 _25029_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1151 _25067_/Q vssd1 vssd1 vccd1 vccd1 _17864_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1162 _16772_/Y vssd1 vssd1 vccd1 vccd1 _25549_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1173 _25784_/Q vssd1 vssd1 vccd1 vccd1 _20426_/B sky130_fd_sc_hd__buf_1
X_24876_ hold880/A hold929/A _24944_/S vssd1 vssd1 vccd1 vccd1 _24877_/B sky130_fd_sc_hd__mux2_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _12840_/X _12888_/X _12827_/X _12889_/X vssd1 vssd1 vccd1 vccd1 _12890_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 _13119_/X vssd1 vssd1 vccd1 vccd1 _25072_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1195 _25095_/Q vssd1 vssd1 vccd1 vccd1 _18618_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23827_ _23827_/A vssd1 vssd1 vccd1 vccd1 _26013_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ _14560_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14560_/Y sky130_fd_sc_hd__nand2_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23758_ hold2156/X _14788_/B _23831_/S vssd1 vssd1 vccd1 vccd1 _23759_/A sky130_fd_sc_hd__mux2_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ hold937/A vssd1 vssd1 vccd1 vccd1 _18122_/B sky130_fd_sc_hd__inv_2
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22709_ _22709_/A _22709_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22711_/A sky130_fd_sc_hd__or3_1
XFILLER_0_32_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ _14491_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14491_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_165_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23689_ _23689_/A vssd1 vssd1 vccd1 vccd1 _25968_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _16227_/A _16227_/B _16245_/B _16229_/Y vssd1 vssd1 vccd1 vccd1 _16230_/X
+ sky130_fd_sc_hd__a31o_1
X_25428_ _25483_/CLK _25428_/D vssd1 vssd1 vccd1 vccd1 _25428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13442_ _13522_/A _13440_/X _23629_/B _13441_/X vssd1 vssd1 vccd1 vccd1 _13442_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16161_ _16161_/A _16161_/B vssd1 vssd1 vccd1 vccd1 _16161_/Y sky130_fd_sc_hd__nand2_1
X_13373_ _13220_/X _14641_/A _13242_/X _19715_/A vssd1 vssd1 vccd1 vccd1 _13373_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25359_ _26184_/CLK hold370/X vssd1 vssd1 vccd1 vccd1 hold368/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15112_ _15270_/A _15269_/B _15111_/Y vssd1 vssd1 vccd1 vccd1 _15112_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_90_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16092_ hold593/X vssd1 vssd1 vccd1 vccd1 _16095_/B sky130_fd_sc_hd__inv_2
XFILLER_0_50_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15043_ _15043_/A _15043_/B vssd1 vssd1 vccd1 vccd1 _15051_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_146_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19920_ _26270_/Q hold659/X vssd1 vssd1 vccd1 vccd1 _19920_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19851_ _19843_/X _19850_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19851_/Y sky130_fd_sc_hd__o21ai_1
X_18802_ _18986_/A _19574_/A vssd1 vssd1 vccd1 vccd1 _18802_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_101_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19782_ _19975_/A _19782_/B vssd1 vssd1 vccd1 vccd1 _19782_/Y sky130_fd_sc_hd__nand2_1
X_16994_ _25903_/Q _25902_/Q vssd1 vssd1 vccd1 vccd1 _17688_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_78_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18733_ _18793_/A _18733_/B _18894_/C vssd1 vssd1 vccd1 vccd1 _18734_/C sky130_fd_sc_hd__nand3_1
X_15945_ _15897_/X _15942_/A _15944_/X vssd1 vssd1 vccd1 vccd1 _15945_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18664_ _19729_/A vssd1 vssd1 vccd1 vccd1 _22370_/B sky130_fd_sc_hd__inv_2
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15876_ _15956_/A hold774/X vssd1 vssd1 vccd1 vccd1 hold775/A sky130_fd_sc_hd__nand2_1
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17615_ _17615_/A _17615_/B vssd1 vssd1 vccd1 vccd1 _17616_/B sky130_fd_sc_hd__xnor2_1
X_14827_ _14827_/A vssd1 vssd1 vccd1 vccd1 _15013_/A sky130_fd_sc_hd__inv_2
X_18595_ _18798_/A _18940_/A vssd1 vssd1 vccd1 vccd1 _18596_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_176_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17546_ _17605_/A _17546_/B vssd1 vssd1 vccd1 vccd1 _17546_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_54_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14758_ _14758_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14758_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13709_ _26251_/Q _13612_/X _13605_/X _13708_/Y vssd1 vssd1 vccd1 vccd1 _13710_/B
+ sky130_fd_sc_hd__a22o_1
X_17477_ _17526_/A _17644_/B vssd1 vssd1 vccd1 vccd1 _17478_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14689_ _14687_/Y hold276/X _14646_/X vssd1 vssd1 vccd1 vccd1 hold277/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19216_ _19216_/A _20507_/B vssd1 vssd1 vccd1 vccd1 _19216_/Y sky130_fd_sc_hd__nor2_1
X_16428_ _16428_/A _16441_/A vssd1 vssd1 vccd1 vccd1 _16430_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19147_ _19144_/X _19145_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19147_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16359_ _16374_/B _16359_/B vssd1 vssd1 vccd1 vccd1 _16360_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19078_ _19186_/A _19078_/B vssd1 vssd1 vccd1 vccd1 _19078_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_124_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18029_ _25853_/Q _22218_/A vssd1 vssd1 vccd1 vccd1 _18037_/A sky130_fd_sc_hd__or2_2
XFILLER_0_160_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21040_ _26305_/Q hold482/X vssd1 vssd1 vccd1 vccd1 _21040_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22991_ _22991_/A _22991_/B vssd1 vssd1 vccd1 vccd1 _22993_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_119_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24730_ _24730_/A vssd1 vssd1 vccd1 vccd1 _26305_/D sky130_fd_sc_hd__clkbuf_1
X_21942_ _21943_/B _21943_/A vssd1 vssd1 vccd1 vccd1 _21944_/A sky130_fd_sc_hd__or2_1
XFILLER_0_179_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21873_ _21874_/B _21874_/A vssd1 vssd1 vccd1 vccd1 _21875_/A sky130_fd_sc_hd__or2_1
X_24661_ hold2734/X hold2718/X _24664_/S vssd1 vssd1 vccd1 vccd1 _24662_/A sky130_fd_sc_hd__mux2_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23612_ _23612_/A vssd1 vssd1 vccd1 vccd1 _25943_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20824_ _20824_/A _20824_/B vssd1 vssd1 vccd1 vccd1 _20826_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24592_ _24592_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24593_/A sky130_fd_sc_hd__and2_1
XFILLER_0_148_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26331_ _26334_/CLK _26331_/D vssd1 vssd1 vccd1 vccd1 _26331_/Q sky130_fd_sc_hd__dfxtp_2
X_23543_ _23537_/X _23542_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _23543_/X sky130_fd_sc_hd__mux2_1
X_20755_ _23117_/B vssd1 vssd1 vccd1 vccd1 _22595_/B sky130_fd_sc_hd__inv_2
XFILLER_0_175_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23474_ _23471_/Y _23473_/Y _24957_/S vssd1 vssd1 vccd1 vccd1 _23474_/X sky130_fd_sc_hd__mux2_1
X_26262_ _26267_/CLK _26262_/D vssd1 vssd1 vccd1 vccd1 _26262_/Q sky130_fd_sc_hd__dfxtp_2
X_20686_ _20686_/A _20686_/B _21319_/C vssd1 vssd1 vccd1 vccd1 _20690_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_135_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22425_ _22680_/A _22425_/B vssd1 vssd1 vccd1 vccd1 _22425_/X sky130_fd_sc_hd__or2_1
X_25213_ _26292_/CLK hold658/X vssd1 vssd1 vccd1 vccd1 hold656/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26193_ _26193_/CLK _26193_/D vssd1 vssd1 vccd1 vccd1 _26193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22356_ _22792_/A _22940_/B vssd1 vssd1 vccd1 vccd1 _22359_/A sky130_fd_sc_hd__nand2_1
X_25144_ _26226_/CLK hold448/X vssd1 vssd1 vccd1 vccd1 hold446/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21307_ _22704_/A vssd1 vssd1 vccd1 vccd1 _21599_/B sky130_fd_sc_hd__buf_6
XFILLER_0_27_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25075_ _25783_/CLK _25075_/D vssd1 vssd1 vccd1 vccd1 _25075_/Q sky130_fd_sc_hd__dfxtp_1
X_22287_ _22287_/A _22287_/B _23170_/A vssd1 vssd1 vccd1 vccd1 _22287_/Y sky130_fd_sc_hd__nand3_1
X_24026_ hold2458/X hold2402/X _24047_/S vssd1 vssd1 vccd1 vccd1 _24027_/A sky130_fd_sc_hd__mux2_1
Xhold270 hold270/A vssd1 vssd1 vccd1 vccd1 hold270/X sky130_fd_sc_hd__dlygate4sd3_1
X_21238_ _21238_/A _21238_/B vssd1 vssd1 vccd1 vccd1 _21241_/B sky130_fd_sc_hd__nand2_1
Xhold281 hold281/A vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 hold292/A vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
X_21169_ _21169_/A _21169_/B _21169_/C vssd1 vssd1 vccd1 vccd1 _21173_/A sky130_fd_sc_hd__nand3_1
X_25977_ _26041_/CLK _25977_/D vssd1 vssd1 vccd1 vccd1 _25977_/Q sky130_fd_sc_hd__dfxtp_1
X_13991_ _26296_/Q _13988_/X _13981_/X _13990_/Y vssd1 vssd1 vccd1 vccd1 _13992_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15730_ _15730_/A _16946_/A vssd1 vssd1 vccd1 vccd1 _15731_/B sky130_fd_sc_hd__nor2_1
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24928_ _24867_/S _24921_/Y _24923_/Y _24927_/X vssd1 vssd1 vccd1 vccd1 _24928_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _12891_/X _14403_/A _12909_/X _25619_/Q vssd1 vssd1 vccd1 vccd1 _12942_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15661_ _15692_/A _15662_/A vssd1 vssd1 vccd1 vccd1 _15661_/X sky130_fd_sc_hd__or2_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24859_ _24855_/X _24858_/X _25910_/Q vssd1 vssd1 vccd1 vccd1 _24859_/X sky130_fd_sc_hd__mux2_1
X_12873_ _26109_/Q _12748_/X _12872_/X vssd1 vssd1 vccd1 vccd1 _12873_/X sky130_fd_sc_hd__a21o_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _19560_/A _17400_/B vssd1 vssd1 vccd1 vccd1 _17629_/B sky130_fd_sc_hd__xor2_4
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _14645_/A hold356/X vssd1 vssd1 vccd1 vccd1 hold357/A sky130_fd_sc_hd__nand2_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18380_ _21211_/B _19532_/A vssd1 vssd1 vccd1 vccd1 _18381_/B sky130_fd_sc_hd__nand2_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _15579_/X _15612_/A _15591_/Y vssd1 vssd1 vccd1 vccd1 _15592_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17331_ _17608_/A _17331_/B vssd1 vssd1 vccd1 vccd1 _17331_/X sky130_fd_sc_hd__xor2_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _14585_/A hold266/X vssd1 vssd1 vccd1 vccd1 hold267/A sky130_fd_sc_hd__nand2_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17262_ _20936_/B _25863_/Q _20962_/B vssd1 vssd1 vccd1 vccd1 _17263_/B sky130_fd_sc_hd__mux2_2
X_14474_ _14525_/A hold194/X vssd1 vssd1 vccd1 vccd1 hold195/A sky130_fd_sc_hd__nand2_1
XFILLER_0_148_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19001_ _19186_/A _19758_/A vssd1 vssd1 vccd1 vccd1 _19001_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16213_ _16211_/X _16212_/Y _16076_/X vssd1 vssd1 vccd1 vccd1 hold913/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13425_ _13522_/A _13423_/X _23629_/B _13424_/X vssd1 vssd1 vccd1 vccd1 _13425_/X
+ sky130_fd_sc_hd__o211a_1
X_17193_ _20780_/B _25858_/Q _25794_/Q vssd1 vssd1 vccd1 vccd1 _17194_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_148_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16144_ _16212_/A hold964/X vssd1 vssd1 vccd1 vccd1 _16144_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_122_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13356_ _26194_/Q _13239_/X _13355_/X vssd1 vssd1 vccd1 vccd1 _13356_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_178_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16075_ _16212_/A hold548/X vssd1 vssd1 vccd1 vccd1 hold549/A sky130_fd_sc_hd__nand2_1
X_13287_ _18719_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13287_/X sky130_fd_sc_hd__or2_1
X_15026_ _15027_/B _15027_/A vssd1 vssd1 vccd1 vccd1 _15028_/A sky130_fd_sc_hd__or2_1
X_19903_ _19896_/X _19902_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19903_/Y sky130_fd_sc_hd__o21ai_1
X_19834_ _19835_/B _19835_/A vssd1 vssd1 vccd1 vccd1 _19834_/X sky130_fd_sc_hd__or2_1
Xhold1909 _26160_/Q vssd1 vssd1 vccd1 vccd1 hold1909/X sky130_fd_sc_hd__dlygate4sd3_1
X_16977_ _16977_/A _16977_/B vssd1 vssd1 vccd1 vccd1 _16977_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19765_ _19762_/X _19763_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19765_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 io_in[4] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_2
X_15928_ _15926_/Y hold552/X _15805_/X vssd1 vssd1 vccd1 vccd1 hold553/A sky130_fd_sc_hd__a21oi_1
X_18716_ _18716_/A _20478_/A vssd1 vssd1 vccd1 vccd1 _18996_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19696_ _19694_/Y _19695_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19696_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_189_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18647_ _25886_/Q _22347_/A vssd1 vssd1 vccd1 vccd1 _18655_/A sky130_fd_sc_hd__or2_2
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15859_ _15859_/A _15869_/A vssd1 vssd1 vccd1 vccd1 _15859_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_189_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18578_ _18576_/X _18269_/X _18577_/X vssd1 vssd1 vccd1 vccd1 _18579_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17529_ _17624_/A _17529_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17529_/X sky130_fd_sc_hd__and3_1
XFILLER_0_46_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20540_ _21042_/A _20540_/B _20539_/X vssd1 vssd1 vccd1 vccd1 _20541_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_129_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20471_ _25850_/Q vssd1 vssd1 vccd1 vccd1 _22136_/B sky130_fd_sc_hd__inv_2
XFILLER_0_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22210_ _22210_/A _22210_/B vssd1 vssd1 vccd1 vccd1 _22210_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_162_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23190_ _26084_/Q vssd1 vssd1 vccd1 vccd1 _23191_/A sky130_fd_sc_hd__inv_2
XFILLER_0_15_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22141_ _22118_/X _22140_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _22141_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22072_ _22774_/B vssd1 vssd1 vccd1 vccd1 _22775_/A sky130_fd_sc_hd__inv_2
XFILLER_0_11_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25900_ _26084_/CLK _25900_/D vssd1 vssd1 vccd1 vccd1 _25900_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21023_ _21025_/B _21025_/C vssd1 vssd1 vccd1 vccd1 _21024_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25831_ _25865_/CLK _25831_/D vssd1 vssd1 vccd1 vccd1 _25831_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_57_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25762_ _25765_/CLK _25762_/D vssd1 vssd1 vccd1 vccd1 _25762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22974_ _22974_/A _22974_/B vssd1 vssd1 vccd1 vccd1 _22976_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24713_ hold2578/X _26300_/Q _24740_/S vssd1 vssd1 vccd1 vccd1 _24713_/X sky130_fd_sc_hd__mux2_1
X_21925_ _18022_/B _17096_/B _18023_/B vssd1 vssd1 vccd1 vccd1 _21926_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_96_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25693_ _26325_/CLK _25693_/D vssd1 vssd1 vccd1 vccd1 _25693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24644_ _24644_/A vssd1 vssd1 vccd1 vccd1 _26277_/D sky130_fd_sc_hd__clkbuf_1
X_21856_ _17931_/B _17064_/B _17932_/B vssd1 vssd1 vccd1 vccd1 _21857_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_78_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20807_ _20807_/A _20807_/B vssd1 vssd1 vccd1 vccd1 _20808_/A sky130_fd_sc_hd__nand2_1
X_21787_ _21788_/A _21788_/B _22909_/A vssd1 vssd1 vccd1 vccd1 _21787_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24575_ _26254_/Q hold2708/X _24587_/S vssd1 vssd1 vccd1 vccd1 _24575_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26314_ _26317_/CLK _26314_/D vssd1 vssd1 vccd1 vccd1 _26314_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_167_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23526_ _24944_/S hold305/A _23525_/X vssd1 vssd1 vccd1 vccd1 _23526_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20738_ _21235_/A _20738_/B vssd1 vssd1 vccd1 vccd1 _20738_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_92_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26245_ _26248_/CLK _26245_/D vssd1 vssd1 vccd1 vccd1 _26245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20669_ _20668_/B _20669_/B _20669_/C vssd1 vssd1 vccd1 vccd1 _20670_/B sky130_fd_sc_hd__nand3b_1
X_23457_ _23445_/X _23456_/X _24949_/S vssd1 vssd1 vccd1 vccd1 _23457_/X sky130_fd_sc_hd__mux2_4
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13210_ _13049_/X _14560_/A _13067_/X _19345_/A vssd1 vssd1 vccd1 vccd1 _13210_/X
+ sky130_fd_sc_hd__a22o_1
X_22408_ _25825_/Q _22408_/B vssd1 vssd1 vccd1 vccd1 _22408_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_34_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26176_ _26181_/CLK _26176_/D vssd1 vssd1 vccd1 vccd1 _26176_/Q sky130_fd_sc_hd__dfxtp_1
X_14190_ _18714_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14190_/Y sky130_fd_sc_hd__nor2_1
X_23388_ _23385_/Y _23387_/Y _24858_/S vssd1 vssd1 vccd1 vccd1 _23388_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25127_ _25708_/CLK _25127_/D vssd1 vssd1 vccd1 vccd1 _25127_/Q sky130_fd_sc_hd__dfxtp_1
X_13141_ _26288_/Q _25657_/Q vssd1 vssd1 vccd1 vccd1 _14524_/A sky130_fd_sc_hd__xor2_1
X_22339_ _22337_/X _22338_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _22339_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_131_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13072_ _26275_/Q _25644_/Q vssd1 vssd1 vccd1 vccd1 _14485_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_103_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25058_ _26142_/CLK _25058_/D vssd1 vssd1 vccd1 vccd1 _25058_/Q sky130_fd_sc_hd__dfxtp_1
X_16900_ _16977_/A _16900_/B vssd1 vssd1 vccd1 vccd1 _16900_/Y sky130_fd_sc_hd__nand2_1
X_24009_ _24009_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24010_/A sky130_fd_sc_hd__and2_1
XFILLER_0_40_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17880_ _17880_/A _25776_/Q vssd1 vssd1 vccd1 vccd1 _20111_/A sky130_fd_sc_hd__nand2_1
X_16831_ _16831_/A _16831_/B vssd1 vssd1 vccd1 vccd1 _16831_/Y sky130_fd_sc_hd__nand2_1
X_19550_ _19551_/B _19551_/A vssd1 vssd1 vccd1 vccd1 _19550_/X sky130_fd_sc_hd__or2_1
X_16762_ _16760_/X _16711_/X _16761_/Y _25869_/Q _14170_/X vssd1 vssd1 vccd1 vccd1
+ _16763_/A sky130_fd_sc_hd__a32o_1
X_13974_ _14000_/A hold760/X vssd1 vssd1 vccd1 vccd1 hold761/A sky130_fd_sc_hd__nand2_1
X_18501_ _22149_/B _25623_/Q vssd1 vssd1 vccd1 vccd1 _18503_/A sky130_fd_sc_hd__nand2_1
X_15713_ _15713_/A _15713_/B vssd1 vssd1 vccd1 vccd1 _15718_/B sky130_fd_sc_hd__nand2_1
X_12925_ _26247_/Q _25616_/Q vssd1 vssd1 vccd1 vccd1 _14394_/A sky130_fd_sc_hd__xor2_1
X_19481_ _19723_/A _19481_/B vssd1 vssd1 vccd1 vccd1 _19481_/Y sky130_fd_sc_hd__nand2_1
X_16693_ _16695_/C vssd1 vssd1 vccd1 vccd1 _16694_/B sky130_fd_sc_hd__inv_2
XFILLER_0_38_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18432_ _18432_/A _21264_/A vssd1 vssd1 vccd1 vccd1 _18778_/A sky130_fd_sc_hd__xor2_4
X_15644_ _15645_/B _15645_/A vssd1 vssd1 vccd1 vccd1 _15644_/X sky130_fd_sc_hd__or2_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _26234_/Q _25603_/Q vssd1 vssd1 vccd1 vccd1 _14355_/A sky130_fd_sc_hd__xor2_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _18445_/A _18367_/B vssd1 vssd1 vccd1 vccd1 _18365_/A sky130_fd_sc_hd__nand2_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _15575_/A _15577_/A vssd1 vssd1 vccd1 vccd1 _15575_/Y sky130_fd_sc_hd__nand2_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12787_ _12746_/X _12785_/X _14910_/B _12786_/X vssd1 vssd1 vccd1 vccd1 _12787_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _25611_/Q vssd1 vssd1 vccd1 vccd1 _21048_/B sky130_fd_sc_hd__inv_2
XFILLER_0_173_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _15464_/A vssd1 vssd1 vccd1 vccd1 _14526_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18294_ _18292_/X _18269_/X _18293_/X vssd1 vssd1 vccd1 vccd1 _18295_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_138_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17245_ _17245_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17245_/Y sky130_fd_sc_hd__nand2_1
X_14457_ _14455_/Y hold54/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13408_ _26331_/Q _19802_/A vssd1 vssd1 vccd1 vccd1 _14660_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_113_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17176_ _17176_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17176_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_98_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14388_ _14388_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14388_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16127_ _16127_/A _16134_/B vssd1 vssd1 vccd1 vccd1 _16127_/Y sky130_fd_sc_hd__nand2_1
X_13339_ _18880_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13339_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16058_ _16028_/Y _16053_/B _16057_/Y vssd1 vssd1 vccd1 vccd1 _16058_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15009_ _15015_/A _15010_/A vssd1 vssd1 vccd1 vccd1 _15009_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2407 _15311_/Y vssd1 vssd1 vccd1 vccd1 hold2407/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2418 _26064_/Q vssd1 vssd1 vccd1 vccd1 hold2418/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2429 _12576_/X vssd1 vssd1 vccd1 vccd1 _12577_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1706 _25880_/Q vssd1 vssd1 vccd1 vccd1 _22855_/B sky130_fd_sc_hd__dlygate4sd3_1
X_19817_ _20634_/A _22513_/B _25637_/Q vssd1 vssd1 vccd1 vccd1 _20639_/C sky130_fd_sc_hd__nand3_1
Xhold1717 _25817_/Q vssd1 vssd1 vccd1 vccd1 _21396_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1728 _25595_/Q vssd1 vssd1 vccd1 vccd1 _17203_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1739 _17178_/Y vssd1 vssd1 vccd1 vccd1 _25593_/D sky130_fd_sc_hd__dlygate4sd3_1
X_19748_ _19749_/B _19749_/A vssd1 vssd1 vccd1 vccd1 _19748_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19679_ _19677_/X _19678_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19679_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21710_ _21710_/A _21710_/B _21710_/C vssd1 vssd1 vccd1 vccd1 _21711_/B sky130_fd_sc_hd__nand3_1
X_22690_ _22688_/X _22689_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22690_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21641_ _21692_/B _21645_/B vssd1 vssd1 vccd1 vccd1 _21643_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21572_ _21572_/A _22902_/B vssd1 vssd1 vccd1 vccd1 _21572_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24360_ hold2265/X _26185_/Q _24433_/S vssd1 vssd1 vccd1 vccd1 _24360_/X sky130_fd_sc_hd__mux2_1
XANTENNA_10 _24867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_21 _17594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_32 _19038_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23311_ _23314_/A _23377_/B _23311_/C vssd1 vssd1 vccd1 vccd1 _23311_/X sky130_fd_sc_hd__and3_1
XANTENNA_43 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20523_ _20526_/A _20526_/C vssd1 vssd1 vccd1 vccd1 _20525_/A sky130_fd_sc_hd__nand2_1
XANTENNA_54 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_24291_ _24291_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24292_/A sky130_fd_sc_hd__and2_1
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_65 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_76 _25849_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26030_ _26032_/CLK _26030_/D vssd1 vssd1 vccd1 vccd1 _26030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23242_ _23242_/A vssd1 vssd1 vccd1 vccd1 _24950_/B sky130_fd_sc_hd__inv_2
XFILLER_0_127_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20454_ _21249_/C _21547_/A vssd1 vssd1 vccd1 vccd1 _20455_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_16_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23173_ _15793_/B _22893_/A _22829_/A vssd1 vssd1 vccd1 vccd1 _23173_/Y sky130_fd_sc_hd__a21oi_1
X_20385_ _20385_/A _20385_/B vssd1 vssd1 vccd1 vccd1 _20386_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22124_ _25878_/Q _22125_/A vssd1 vssd1 vccd1 vccd1 _22126_/A sky130_fd_sc_hd__or2_1
XFILLER_0_101_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22055_ _22055_/A _23042_/A _22055_/C vssd1 vssd1 vccd1 vccd1 _22055_/Y sky130_fd_sc_hd__nand3_1
X_21006_ _21532_/B _21483_/B vssd1 vssd1 vccd1 vccd1 _21007_/B sky130_fd_sc_hd__nand2_1
X_25814_ _25817_/CLK _25814_/D vssd1 vssd1 vccd1 vccd1 _25814_/Q sky130_fd_sc_hd__dfxtp_2
X_25745_ _25745_/CLK _25745_/D vssd1 vssd1 vccd1 vccd1 _25745_/Q sky130_fd_sc_hd__dfxtp_1
X_22957_ _22957_/A _22957_/B vssd1 vssd1 vccd1 vccd1 _22959_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_173_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12710_ _24987_/Q _24986_/Q _24985_/Q _24984_/Q vssd1 vssd1 vccd1 vccd1 _12711_/A
+ sky130_fd_sc_hd__and4_1
X_21908_ _21909_/B _21909_/A vssd1 vssd1 vccd1 vccd1 _21910_/A sky130_fd_sc_hd__or2_1
X_25676_ _26305_/CLK _25676_/D vssd1 vssd1 vccd1 vccd1 _25676_/Q sky130_fd_sc_hd__dfxtp_1
X_13690_ _26248_/Q _13612_/X _13605_/X _13689_/Y vssd1 vssd1 vccd1 vccd1 _13691_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_179_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22888_ _22937_/A _22888_/B vssd1 vssd1 vccd1 vccd1 _22888_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_35_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12641_ _12641_/A vssd1 vssd1 vccd1 vccd1 _24981_/D sky130_fd_sc_hd__clkbuf_1
X_24627_ hold2634/X _26272_/Q _24664_/S vssd1 vssd1 vccd1 vccd1 _24627_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_167_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21839_ _21840_/B _21840_/A vssd1 vssd1 vccd1 vccd1 _21841_/A sky130_fd_sc_hd__or2_1
XFILLER_0_155_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15360_ _15361_/B _15361_/A vssd1 vssd1 vccd1 vccd1 _15360_/X sky130_fd_sc_hd__or2_1
X_12572_ _12572_/A vssd1 vssd1 vccd1 vccd1 _24967_/D sky130_fd_sc_hd__clkbuf_1
X_24558_ _24558_/A vssd1 vssd1 vccd1 vccd1 _26249_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14311_ _14344_/A hold140/X vssd1 vssd1 vccd1 vccd1 hold141/A sky130_fd_sc_hd__nand2_1
XFILLER_0_163_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23509_ hold128/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23509_/X sky130_fd_sc_hd__or2b_1
X_15291_ _15291_/A _15290_/Y vssd1 vssd1 vccd1 vccd1 _15307_/A sky130_fd_sc_hd__or2b_1
XFILLER_0_108_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24489_ hold2555/X _26227_/Q _24510_/S vssd1 vssd1 vccd1 vccd1 _24489_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17030_ _17028_/X _23187_/B _17029_/X vssd1 vssd1 vccd1 vccd1 _17031_/A sky130_fd_sc_hd__a21o_1
X_14242_ _14260_/A hold845/X vssd1 vssd1 vccd1 vccd1 _14242_/Y sky130_fd_sc_hd__nand2_1
X_26228_ _26232_/CLK _26228_/D vssd1 vssd1 vccd1 vccd1 _26228_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_180_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26159_ _26244_/CLK _26159_/D vssd1 vssd1 vccd1 vccd1 _26159_/Q sky130_fd_sc_hd__dfxtp_1
X_14173_ _26325_/Q _13988_/X _14170_/X _14172_/Y vssd1 vssd1 vccd1 vccd1 _14174_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13124_ _13109_/X _13122_/X _13096_/X _13123_/X vssd1 vssd1 vccd1 vccd1 _13124_/X
+ sky130_fd_sc_hd__o211a_1
X_18981_ _18981_/A _19052_/B vssd1 vssd1 vccd1 vccd1 _18982_/B sky130_fd_sc_hd__xnor2_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17932_ _20141_/A _17932_/B vssd1 vssd1 vccd1 vccd1 _19137_/A sky130_fd_sc_hd__nand2_2
X_13055_ _26272_/Q _25641_/Q vssd1 vssd1 vccd1 vccd1 _14476_/A sky130_fd_sc_hd__xor2_1
X_17863_ _19025_/A _17863_/B vssd1 vssd1 vccd1 vccd1 _17863_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19602_ _19602_/A _20055_/B vssd1 vssd1 vccd1 vccd1 _19602_/Y sky130_fd_sc_hd__nor2_1
X_16814_ _16812_/Y _16813_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16814_/Y sky130_fd_sc_hd__a21oi_1
X_17794_ _17794_/A vssd1 vssd1 vccd1 vccd1 _18083_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16745_ _16980_/A _16750_/B vssd1 vssd1 vccd1 vccd1 _16747_/B sky130_fd_sc_hd__nand2_1
X_19533_ _21210_/A _21981_/B _25617_/Q vssd1 vssd1 vccd1 vccd1 _21214_/C sky130_fd_sc_hd__nand3_1
X_13957_ _25788_/Q vssd1 vssd1 vccd1 vccd1 _17990_/B sky130_fd_sc_hd__inv_2
X_19464_ _19462_/X _19463_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19464_/Y sky130_fd_sc_hd__a21oi_1
X_12908_ _26244_/Q _25613_/Q vssd1 vssd1 vccd1 vccd1 _14385_/A sky130_fd_sc_hd__xor2_1
X_16676_ _16676_/A _16676_/B vssd1 vssd1 vccd1 vccd1 _16678_/A sky130_fd_sc_hd__or2_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13888_ _14000_/A hold851/X vssd1 vssd1 vccd1 vccd1 _13888_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15627_ _15615_/X _15693_/B _15233_/X vssd1 vssd1 vccd1 vccd1 _15627_/Y sky130_fd_sc_hd__a21oi_1
X_18415_ _18535_/A _18415_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18415_/X sky130_fd_sc_hd__and3_1
X_12839_ _12746_/X _12837_/X _12827_/X _12838_/X vssd1 vssd1 vccd1 vccd1 _12839_/X
+ sky130_fd_sc_hd__o211a_1
X_19395_ _19387_/X _19394_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19395_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18346_ _18951_/A _25743_/Q vssd1 vssd1 vccd1 vccd1 _18348_/A sky130_fd_sc_hd__nand2_1
X_15558_ _15827_/A _15822_/B _15822_/A _15557_/Y vssd1 vssd1 vccd1 vccd1 _15560_/A
+ sky130_fd_sc_hd__a31o_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14509_ _14509_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14509_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18277_ _21810_/B _25612_/Q vssd1 vssd1 vccd1 vccd1 _18279_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_83_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15489_ _15489_/A _15776_/B vssd1 vssd1 vccd1 vccd1 _15490_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_182_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17228_ _17226_/X _23187_/B _17227_/X vssd1 vssd1 vccd1 vccd1 _17229_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold803 hold803/A vssd1 vssd1 vccd1 vccd1 hold803/X sky130_fd_sc_hd__buf_1
X_17159_ _17485_/A _17562_/A vssd1 vssd1 vccd1 vccd1 _17160_/B sky130_fd_sc_hd__xnor2_1
Xhold814 hold814/A vssd1 vssd1 vccd1 vccd1 hold814/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 hold825/A vssd1 vssd1 vccd1 vccd1 hold825/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold836 hold836/A vssd1 vssd1 vccd1 vccd1 hold836/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 hold847/A vssd1 vssd1 vccd1 vccd1 hold847/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 hold858/A vssd1 vssd1 vccd1 vccd1 hold858/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20170_ _20170_/A _20170_/B vssd1 vssd1 vccd1 vccd1 _20172_/A sky130_fd_sc_hd__nand2_1
Xhold869 hold869/A vssd1 vssd1 vccd1 vccd1 hold869/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2204 _14942_/Y vssd1 vssd1 vccd1 vccd1 hold2204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2215 _24424_/X vssd1 vssd1 vccd1 vccd1 _24425_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2226 _26100_/Q vssd1 vssd1 vccd1 vccd1 hold2226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2237 _26150_/Q vssd1 vssd1 vccd1 vccd1 hold2237/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1503 _25105_/Q vssd1 vssd1 vccd1 vccd1 _18819_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2248 _14994_/Y vssd1 vssd1 vccd1 vccd1 _25423_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1514 _16840_/Y vssd1 vssd1 vccd1 vccd1 _25559_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2259 _25977_/Q vssd1 vssd1 vccd1 vccd1 hold2259/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1525 _25796_/Q vssd1 vssd1 vccd1 vccd1 _20880_/B sky130_fd_sc_hd__clkbuf_2
Xhold1536 _21209_/Y vssd1 vssd1 vccd1 vccd1 _25808_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23860_ _23860_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23861_/A sky130_fd_sc_hd__and2_1
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1547 _25602_/Q vssd1 vssd1 vccd1 vccd1 _17299_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1558 _19811_/Y vssd1 vssd1 vccd1 vccd1 _25758_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1569 _20271_/Y vssd1 vssd1 vccd1 vccd1 _25780_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22811_ _22811_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22811_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23791_ _14875_/B _14884_/B _23831_/S vssd1 vssd1 vccd1 vccd1 _23792_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_95_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25530_ _25534_/CLK hold919/X vssd1 vssd1 vccd1 vccd1 hold918/A sky130_fd_sc_hd__dfxtp_1
X_22742_ _23055_/B _22742_/B vssd1 vssd1 vccd1 vccd1 _22744_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_149_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25461_ _26012_/CLK _25461_/D vssd1 vssd1 vccd1 vccd1 _25461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22673_ _23151_/B _23008_/B vssd1 vssd1 vccd1 vccd1 _22675_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_109_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xascon_wrapper_16 vssd1 vssd1 vccd1 vccd1 io_oeb[2] ascon_wrapper_16/LO sky130_fd_sc_hd__conb_1
XFILLER_0_165_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24412_ hold2276/X hold1989/X _24433_/S vssd1 vssd1 vccd1 vccd1 _24413_/A sky130_fd_sc_hd__mux2_1
X_21624_ _21622_/Y _21623_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21624_/Y sky130_fd_sc_hd__a21oi_1
X_25392_ _26001_/CLK _25392_/D vssd1 vssd1 vccd1 vccd1 _25392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24343_ _24343_/A vssd1 vssd1 vccd1 vccd1 _26179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21555_ _21555_/A _21555_/B vssd1 vssd1 vccd1 vccd1 _21556_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_173_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20506_ _20506_/A _22160_/B vssd1 vssd1 vccd1 vccd1 _20507_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_106_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21486_ _26326_/Q _21228_/X hold698/X vssd1 vssd1 vccd1 vccd1 _21489_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24274_ _24274_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24275_/A sky130_fd_sc_hd__and2_1
XFILLER_0_133_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26013_ _26014_/CLK _26013_/D vssd1 vssd1 vccd1 vccd1 _26013_/Q sky130_fd_sc_hd__dfxtp_1
X_23225_ _25909_/Q vssd1 vssd1 vccd1 vccd1 _24858_/S sky130_fd_sc_hd__buf_12
XFILLER_0_121_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20437_ _21249_/C vssd1 vssd1 vccd1 vccd1 _21252_/B sky130_fd_sc_hd__inv_2
XFILLER_0_31_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23156_ _23188_/A _23156_/B vssd1 vssd1 vccd1 vccd1 _23156_/X sky130_fd_sc_hd__or2_1
X_20368_ _20370_/B vssd1 vssd1 vccd1 vccd1 _20369_/B sky130_fd_sc_hd__inv_2
XFILLER_0_105_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22107_ _17859_/B _25593_/Q _17860_/B vssd1 vssd1 vccd1 vccd1 _22108_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23087_ _23087_/A _23087_/B vssd1 vssd1 vccd1 vccd1 _23089_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_140_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20299_ _20299_/A _20299_/B vssd1 vssd1 vccd1 vccd1 _20300_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22038_ _22038_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _22038_/X sky130_fd_sc_hd__and2_1
X_14860_ _14860_/A _22293_/A vssd1 vssd1 vccd1 vccd1 _22292_/B sky130_fd_sc_hd__xnor2_2
X_13811_ _13823_/A _13811_/B vssd1 vssd1 vccd1 vccd1 _13811_/Y sky130_fd_sc_hd__nand2_1
X_14791_ _14791_/A vssd1 vssd1 vccd1 vccd1 _14980_/A sky130_fd_sc_hd__inv_2
X_23989_ hold2418/X hold2053/X _24001_/S vssd1 vssd1 vccd1 vccd1 _23990_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16530_ _16698_/A hold864/X vssd1 vssd1 vccd1 vccd1 _16530_/Y sky130_fd_sc_hd__nand2_1
X_25728_ _25729_/CLK _25728_/D vssd1 vssd1 vccd1 vccd1 _25728_/Q sky130_fd_sc_hd__dfxtp_1
X_13742_ _13760_/A hold584/X vssd1 vssd1 vccd1 vccd1 hold585/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16461_ _16461_/A _16461_/B vssd1 vssd1 vccd1 vccd1 _16487_/A sky130_fd_sc_hd__and2_1
XFILLER_0_112_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25659_ _26292_/CLK _25659_/D vssd1 vssd1 vccd1 vccd1 _25659_/Q sky130_fd_sc_hd__dfxtp_1
X_13673_ hold792/X _13672_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold793/A sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_191_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _26283_/CLK sky130_fd_sc_hd__clkbuf_16
X_18200_ _18200_/A _20991_/B _18200_/C vssd1 vssd1 vccd1 vccd1 _20973_/B sky130_fd_sc_hd__nand3_2
X_15412_ _15827_/A _15822_/B _15553_/A vssd1 vssd1 vccd1 vccd1 _15414_/A sky130_fd_sc_hd__a21o_1
X_12624_ _12624_/A _12645_/B vssd1 vssd1 vccd1 vccd1 _12625_/C sky130_fd_sc_hd__nand2_1
X_19180_ _20389_/A _17671_/A _20394_/C vssd1 vssd1 vccd1 vccd1 _19261_/A sky130_fd_sc_hd__o21ai_4
X_16392_ _16394_/B vssd1 vssd1 vccd1 vccd1 _16416_/B sky130_fd_sc_hd__inv_2
XFILLER_0_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18131_ _20909_/B _19373_/A vssd1 vssd1 vccd1 vccd1 _18132_/B sky130_fd_sc_hd__nand2_1
X_15343_ _15331_/X _15406_/B _15233_/X vssd1 vssd1 vccd1 vccd1 _15343_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12555_ _17685_/C vssd1 vssd1 vccd1 vccd1 _23201_/B sky130_fd_sc_hd__inv_2
XFILLER_0_0_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18062_ _18060_/Y _18061_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _25651_/D sky130_fd_sc_hd__a21oi_1
X_15274_ _15220_/X _15268_/A _15273_/X vssd1 vssd1 vccd1 vccd1 _15275_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12486_ _12733_/A _23191_/C vssd1 vssd1 vccd1 vccd1 _14893_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17013_ _23199_/A vssd1 vssd1 vccd1 vccd1 _22586_/A sky130_fd_sc_hd__clkinv_8
X_14225_ _25831_/Q vssd1 vssd1 vccd1 vccd1 _18834_/B sky130_fd_sc_hd__inv_2
XFILLER_0_184_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14156_ _14150_/Y _14154_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold826/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ _18008_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13107_/X sky130_fd_sc_hd__or2_1
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _14082_/Y _14086_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold790/A sky130_fd_sc_hd__a21oi_1
X_18964_ _18986_/A _19687_/A vssd1 vssd1 vccd1 vccd1 _18964_/Y sky130_fd_sc_hd__nand2_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17915_ _17913_/X _17528_/X _17914_/X vssd1 vssd1 vccd1 vccd1 _17916_/A sky130_fd_sc_hd__a21o_1
X_13038_ _13018_/X _13036_/X _13005_/X _13037_/X vssd1 vssd1 vccd1 vccd1 _13038_/X
+ sky130_fd_sc_hd__o211a_1
X_18895_ _18895_/A _18895_/B _18895_/C vssd1 vssd1 vccd1 vccd1 _22642_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17846_ _18529_/A _17846_/B _18529_/C vssd1 vssd1 vccd1 vccd1 _17847_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_179_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14989_ _14989_/A _14989_/B vssd1 vssd1 vccd1 vccd1 _14990_/B sky130_fd_sc_hd__nand2_1
X_17777_ _17764_/X _17722_/A _17763_/Y _22786_/A vssd1 vssd1 vccd1 vccd1 _17779_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19516_ _19515_/Y _19272_/X _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19517_/B
+ sky130_fd_sc_hd__a211o_1
X_16728_ _16728_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16728_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16659_ _16681_/A _16659_/B vssd1 vssd1 vccd1 vccd1 _16670_/A sky130_fd_sc_hd__nand2_1
X_19447_ _19463_/B _19537_/B vssd1 vssd1 vccd1 vccd1 _19449_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_182_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _25802_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19378_ _19378_/A _19378_/B vssd1 vssd1 vccd1 vccd1 _19378_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18329_ _21136_/C _21880_/A vssd1 vssd1 vccd1 vccd1 _21128_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21340_ _21340_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21345_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21271_ _21270_/B _21271_/B _21271_/C vssd1 vssd1 vccd1 vccd1 _21272_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_13_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold600 hold600/A vssd1 vssd1 vccd1 vccd1 hold600/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 hold611/A vssd1 vssd1 vccd1 vccd1 hold611/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_130_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold622 hold622/A vssd1 vssd1 vccd1 vccd1 hold622/X sky130_fd_sc_hd__dlygate4sd3_1
X_23010_ _23010_/A _23010_/B vssd1 vssd1 vccd1 vccd1 _23011_/A sky130_fd_sc_hd__xor2_1
Xhold633 hold633/A vssd1 vssd1 vccd1 vccd1 hold633/X sky130_fd_sc_hd__dlygate4sd3_1
X_20222_ _20224_/A _20224_/B vssd1 vssd1 vccd1 vccd1 _20223_/A sky130_fd_sc_hd__nand2_1
Xhold644 hold644/A vssd1 vssd1 vccd1 vccd1 hold644/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold655 hold655/A vssd1 vssd1 vccd1 vccd1 hold655/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold666 hold666/A vssd1 vssd1 vccd1 vccd1 hold666/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 hold677/A vssd1 vssd1 vccd1 vccd1 hold677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 hold688/A vssd1 vssd1 vccd1 vccd1 hold688/X sky130_fd_sc_hd__dlygate4sd3_1
X_20153_ _20153_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20158_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_110_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold699 hold699/A vssd1 vssd1 vccd1 vccd1 hold699/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2001 _26136_/Q vssd1 vssd1 vccd1 vccd1 hold2001/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2012 _12715_/X vssd1 vssd1 vccd1 vccd1 _12716_/A sky130_fd_sc_hd__dlygate4sd3_1
X_24961_ _24930_/Y _24950_/Y _24870_/B _24959_/B _24960_/X vssd1 vssd1 vccd1 vccd1
+ _24961_/X sky130_fd_sc_hd__a41o_1
Xhold2023 _25943_/Q vssd1 vssd1 vccd1 vccd1 hold2023/X sky130_fd_sc_hd__dlygate4sd3_1
X_20084_ _20084_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _20084_/Y sky130_fd_sc_hd__nand2_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2034 _26103_/Q vssd1 vssd1 vccd1 vccd1 hold2034/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2045 _25975_/Q vssd1 vssd1 vccd1 vccd1 hold2045/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1300 _25056_/Q vssd1 vssd1 vccd1 vccd1 _17587_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2056 _23350_/X vssd1 vssd1 vccd1 vccd1 _23352_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1311 _14732_/Y vssd1 vssd1 vccd1 vccd1 _25392_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1322 _16908_/Y vssd1 vssd1 vccd1 vccd1 _25569_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23912_ _23912_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23913_/A sky130_fd_sc_hd__and2_1
Xhold2067 _26005_/Q vssd1 vssd1 vccd1 vccd1 hold2067/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24892_ _24881_/X _24891_/X _23255_/A vssd1 vssd1 vccd1 vccd1 _24892_/X sky130_fd_sc_hd__a21o_1
Xhold1333 _25391_/Q vssd1 vssd1 vccd1 vccd1 _14721_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2078 _24299_/X vssd1 vssd1 vccd1 vccd1 _24300_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1344 _14742_/Y vssd1 vssd1 vccd1 vccd1 _25393_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2089 _26207_/Q vssd1 vssd1 vccd1 vccd1 hold2089/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1355 _25760_/Q vssd1 vssd1 vccd1 vccd1 _19838_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1366 _14883_/Y vssd1 vssd1 vccd1 vccd1 _25409_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23843_ _23843_/A vssd1 vssd1 vccd1 vccd1 _26018_/D sky130_fd_sc_hd__clkbuf_1
Xhold1377 _25390_/Q vssd1 vssd1 vccd1 vccd1 _14712_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1388 _16887_/Y vssd1 vssd1 vccd1 vccd1 _25566_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1399 _25726_/Q vssd1 vssd1 vccd1 vccd1 _19353_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23774_ _23774_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23775_/A sky130_fd_sc_hd__and2_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20986_ _20986_/A vssd1 vssd1 vccd1 vccd1 _20986_/X sky130_fd_sc_hd__buf_8
XFILLER_0_71_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25513_ _25515_/CLK hold969/X vssd1 vssd1 vccd1 vccd1 hold968/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22725_ _23184_/B vssd1 vssd1 vccd1 vccd1 _23183_/B sky130_fd_sc_hd__inv_2
XFILLER_0_165_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_173_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _26226_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25444_ _26051_/CLK _25444_/D vssd1 vssd1 vccd1 vccd1 _25444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22656_ _22656_/A _22656_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22658_/A sky130_fd_sc_hd__or3_1
XFILLER_0_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21607_ _21605_/Y _21606_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21607_/Y sky130_fd_sc_hd__a21oi_1
X_25375_ _26200_/CLK hold289/X vssd1 vssd1 vccd1 vccd1 hold287/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22587_ _22937_/A _22587_/B vssd1 vssd1 vccd1 vccd1 _22587_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_168_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24326_ hold2436/X hold2400/X _24356_/S vssd1 vssd1 vccd1 vccd1 _24327_/A sky130_fd_sc_hd__mux2_1
X_21538_ _21636_/A _21538_/B _21537_/X vssd1 vssd1 vccd1 vccd1 _21539_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_44_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24257_ _24257_/A vssd1 vssd1 vccd1 vccd1 _26151_/D sky130_fd_sc_hd__clkbuf_1
X_21469_ _21469_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21474_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_105_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14010_ _18053_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14010_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_142_1228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23208_ _23208_/A _23208_/B vssd1 vssd1 vccd1 vccd1 _23209_/C sky130_fd_sc_hd__nand2_1
X_24188_ _24188_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24189_/A sky130_fd_sc_hd__and2_1
X_23139_ _23139_/A _23187_/B vssd1 vssd1 vccd1 vccd1 _23139_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_101_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15961_ _15961_/A _15961_/B vssd1 vssd1 vccd1 vccd1 _15963_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14912_ _14913_/B _14913_/A vssd1 vssd1 vccd1 vccd1 _14914_/A sky130_fd_sc_hd__or2_1
X_17700_ _17705_/A _17705_/B vssd1 vssd1 vccd1 vccd1 _17703_/A sky130_fd_sc_hd__nand2_1
X_15892_ _15909_/B _15892_/B vssd1 vssd1 vccd1 vccd1 _15921_/B sky130_fd_sc_hd__nand2_1
X_18680_ _18678_/X _18269_/X _18679_/X vssd1 vssd1 vccd1 vccd1 _18681_/A sky130_fd_sc_hd__a21o_1
Xhold2590 _24763_/X vssd1 vssd1 vccd1 vccd1 _24764_/A sky130_fd_sc_hd__dlygate4sd3_1
X_14843_ _14893_/A _14843_/B vssd1 vssd1 vccd1 vccd1 _22233_/A sky130_fd_sc_hd__nand2_1
X_17631_ _19082_/A vssd1 vssd1 vccd1 vccd1 _18535_/A sky130_fd_sc_hd__buf_8
XFILLER_0_37_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17562_ _17562_/A _17615_/A vssd1 vssd1 vccd1 vccd1 _17563_/B sky130_fd_sc_hd__xnor2_1
X_14774_ _25846_/Q _12527_/A _14962_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14774_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16513_ _16513_/A _16513_/B vssd1 vssd1 vccd1 vccd1 _16515_/A sky130_fd_sc_hd__nand2_1
X_19301_ _19300_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19302_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13725_ _25751_/Q vssd1 vssd1 vccd1 vccd1 _18509_/B sky130_fd_sc_hd__inv_2
X_17493_ _17624_/A _17493_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17493_/X sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_164_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _26296_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16444_ _16394_/A _16440_/X _16491_/B vssd1 vssd1 vccd1 vccd1 _16462_/A sky130_fd_sc_hd__a21bo_1
X_19232_ _20546_/A _19230_/Y _20551_/C vssd1 vssd1 vccd1 vccd1 _19322_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_2_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13656_ _13760_/A hold629/X vssd1 vssd1 vccd1 vccd1 hold630/A sky130_fd_sc_hd__nand2_1
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12607_ _12607_/A vssd1 vssd1 vccd1 vccd1 _24974_/D sky130_fd_sc_hd__clkbuf_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19163_ _20349_/A _22051_/A _25591_/Q vssd1 vssd1 vccd1 vccd1 _20354_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_186_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16375_ _16373_/X _16374_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _16375_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_171_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13587_ _25729_/Q vssd1 vssd1 vccd1 vccd1 _17908_/B sky130_fd_sc_hd__inv_2
XFILLER_0_171_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18114_ _25653_/Q vssd1 vssd1 vccd1 vccd1 _21992_/A sky130_fd_sc_hd__inv_2
XFILLER_0_109_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15326_ _15326_/A _15326_/B vssd1 vssd1 vccd1 vccd1 _15327_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_155_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12538_ _15621_/A _12537_/Y _12558_/B vssd1 vssd1 vccd1 vccd1 _24997_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19094_ _20067_/B _20067_/A vssd1 vssd1 vccd1 vccd1 _20068_/A sky130_fd_sc_hd__or2_1
XFILLER_0_42_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18045_ _18529_/A vssd1 vssd1 vccd1 vccd1 _18446_/A sky130_fd_sc_hd__buf_6
X_15257_ _22656_/B _15257_/B vssd1 vssd1 vccd1 vccd1 _22653_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_124_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14208_ _18774_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14208_/Y sky130_fd_sc_hd__nor2_1
X_15188_ _15112_/X _15271_/B _15272_/A vssd1 vssd1 vccd1 vccd1 _15188_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14139_ _25817_/Q vssd1 vssd1 vccd1 vccd1 _18551_/B sky130_fd_sc_hd__inv_2
XFILLER_0_120_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19996_ _19996_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _19996_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18947_ _25709_/Q vssd1 vssd1 vccd1 vccd1 _22718_/B sky130_fd_sc_hd__inv_2
XFILLER_0_158_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18878_ _18878_/A _18878_/B vssd1 vssd1 vccd1 vccd1 _18878_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_146_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17829_ _17829_/A vssd1 vssd1 vccd1 vccd1 _23203_/B sky130_fd_sc_hd__inv_2
X_20840_ _21708_/B _21435_/B vssd1 vssd1 vccd1 vccd1 _20841_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20771_ _26296_/Q _20731_/X hold656/X vssd1 vssd1 vccd1 vccd1 _20774_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_155_clk clkbuf_4_11__f_clk/X vssd1 vssd1 vccd1 vccd1 _26306_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_187_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22510_ _22561_/A _22510_/B vssd1 vssd1 vccd1 vccd1 _22510_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_18_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23490_ hold20/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23490_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22441_ _22441_/A _22441_/B vssd1 vssd1 vccd1 vccd1 _22442_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_134_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25160_ _25743_/CLK hold631/X vssd1 vssd1 vccd1 vccd1 hold629/A sky130_fd_sc_hd__dfxtp_1
X_22372_ _22372_/A _22372_/B vssd1 vssd1 vccd1 vccd1 _22372_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24111_ hold2034/X _26104_/Q _24126_/S vssd1 vssd1 vccd1 vccd1 _24111_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21323_ _21323_/A _21323_/B vssd1 vssd1 vccd1 vccd1 _21324_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_130_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25091_ _26301_/CLK _25091_/D vssd1 vssd1 vccd1 vccd1 _25091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24042_ _24042_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24043_/A sky130_fd_sc_hd__and2_1
X_21254_ _21254_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _21259_/A sky130_fd_sc_hd__nand2_1
Xhold430 hold430/A vssd1 vssd1 vccd1 vccd1 hold430/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold441 hold441/A vssd1 vssd1 vccd1 vccd1 hold441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 hold452/A vssd1 vssd1 vccd1 vccd1 hold452/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 hold463/A vssd1 vssd1 vccd1 vccd1 hold463/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20205_ _20208_/A _20208_/C vssd1 vssd1 vccd1 vccd1 _20207_/A sky130_fd_sc_hd__nand2_1
Xhold474 hold474/A vssd1 vssd1 vccd1 vccd1 hold474/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21185_ _21187_/B _21187_/C vssd1 vssd1 vccd1 vccd1 _21186_/A sky130_fd_sc_hd__nand2_1
Xhold485 hold485/A vssd1 vssd1 vccd1 vccd1 hold485/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 hold496/A vssd1 vssd1 vccd1 vccd1 hold496/X sky130_fd_sc_hd__dlygate4sd3_1
X_20136_ _20139_/A _20139_/B vssd1 vssd1 vccd1 vccd1 _20138_/A sky130_fd_sc_hd__nand2_1
X_25993_ _25998_/CLK _25993_/D vssd1 vssd1 vccd1 vccd1 _25993_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24944_ _16285_/B _16292_/Y _24944_/S vssd1 vssd1 vccd1 vccd1 _24944_/X sky130_fd_sc_hd__mux2_1
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20067_ _20067_/A _20067_/B vssd1 vssd1 vccd1 vccd1 _20068_/B sky130_fd_sc_hd__nand2_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 _13340_/X vssd1 vssd1 vccd1 vccd1 _25108_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 _25021_/Q vssd1 vssd1 vccd1 vccd1 _17282_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1152 _13092_/X vssd1 vssd1 vccd1 vccd1 _25067_/D sky130_fd_sc_hd__dlygate4sd3_1
X_24875_ _24875_/A _24957_/S vssd1 vssd1 vccd1 vccd1 _24875_/Y sky130_fd_sc_hd__nand2_1
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1163 _25030_/Q vssd1 vssd1 vccd1 vccd1 _17383_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1174 _20427_/Y vssd1 vssd1 vccd1 vccd1 _25784_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1185 _25089_/Q vssd1 vssd1 vccd1 vccd1 _18495_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1196 _13258_/X vssd1 vssd1 vccd1 vccd1 _25095_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23826_ _23826_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23827_/A sky130_fd_sc_hd__and2_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23757_ _23920_/S vssd1 vssd1 vccd1 vccd1 _23831_/S sky130_fd_sc_hd__buf_12
XFILLER_0_138_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_146_clk clkbuf_4_11__f_clk/X vssd1 vssd1 vccd1 vccd1 _26317_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20969_ _20969_/A _21977_/B _20969_/C vssd1 vssd1 vccd1 vccd1 _20973_/C sky130_fd_sc_hd__nand3_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13510_ _13522_/A hold768/X vssd1 vssd1 vccd1 vccd1 hold769/A sky130_fd_sc_hd__nand2_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22708_ _26055_/Q vssd1 vssd1 vccd1 vccd1 _22709_/A sky130_fd_sc_hd__inv_2
XFILLER_0_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14490_ _14488_/Y hold81/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__a21oi_1
X_23688_ _23688_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23689_/A sky130_fd_sc_hd__and2_1
XFILLER_0_138_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25427_ _25491_/CLK _25427_/D vssd1 vssd1 vccd1 vccd1 _25427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13441_ _19054_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13441_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22639_ _22639_/A _25898_/Q vssd1 vssd1 vccd1 vccd1 _22639_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_64_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16160_ _16160_/A _16160_/B vssd1 vssd1 vccd1 vccd1 _16171_/A sky130_fd_sc_hd__nand2_1
X_13372_ _26325_/Q _19715_/A vssd1 vssd1 vccd1 vccd1 _14641_/A sky130_fd_sc_hd__xor2_1
X_25358_ _26184_/CLK hold160/X vssd1 vssd1 vccd1 vccd1 hold158/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15111_ _15111_/A _15111_/B vssd1 vssd1 vccd1 vccd1 _15111_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24309_ _24309_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24310_/A sky130_fd_sc_hd__and2_1
X_16091_ _16089_/Y hold764/X _16076_/X vssd1 vssd1 vccd1 vccd1 hold765/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25289_ _26240_/CLK hold244/X vssd1 vssd1 vccd1 vccd1 hold242/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15042_ _15042_/A _15042_/B vssd1 vssd1 vccd1 vccd1 _15043_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_121_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19850_ _19848_/X _19849_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19850_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18801_ _18801_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18801_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19781_ _19773_/X _19780_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19781_/Y sky130_fd_sc_hd__o21ai_1
X_16993_ _17608_/A _16993_/B vssd1 vssd1 vccd1 vccd1 _16993_/X sky130_fd_sc_hd__xor2_1
X_18732_ _18792_/A _25762_/Q vssd1 vssd1 vccd1 vccd1 _18734_/A sky130_fd_sc_hd__nand2_1
X_15944_ _15922_/Y _15941_/A _15943_/Y vssd1 vssd1 vccd1 vccd1 _15944_/X sky130_fd_sc_hd__a21o_1
X_15875_ _15875_/A _16697_/B _15884_/B vssd1 vssd1 vccd1 vccd1 _15875_/Y sky130_fd_sc_hd__nand3_1
X_18663_ _18660_/Y _18662_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25677_/D sky130_fd_sc_hd__a21oi_1
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14826_ _22173_/B _15778_/B vssd1 vssd1 vccd1 vccd1 _14827_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17614_ _17611_/Y _17613_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _25639_/D sky130_fd_sc_hd__a21oi_1
X_18594_ _18594_/A _20235_/A vssd1 vssd1 vccd1 vccd1 _18940_/A sky130_fd_sc_hd__xor2_4
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14757_ _25844_/Q _13466_/A _14756_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14758_/A
+ sky130_fd_sc_hd__a22o_1
X_17545_ _17545_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17545_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_175_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_137_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _25835_/CLK sky130_fd_sc_hd__clkbuf_16
X_13708_ _18449_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13708_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17476_ _17473_/Y _17475_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _25620_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14688_ _14688_/A hold275/X vssd1 vssd1 vccd1 vccd1 hold276/A sky130_fd_sc_hd__nand2_1
XFILLER_0_129_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19215_ _19213_/Y _19214_/Y _19086_/X vssd1 vssd1 vccd1 vccd1 _19215_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_183_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16427_ _16427_/A _16442_/A vssd1 vssd1 vccd1 vccd1 _16441_/B sky130_fd_sc_hd__or2_1
X_13639_ _26240_/Q _13612_/X _13605_/X _13638_/Y vssd1 vssd1 vccd1 vccd1 _13640_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16358_ _16358_/A _16358_/B vssd1 vssd1 vccd1 vccd1 _16359_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_26_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19146_ _21789_/A vssd1 vssd1 vccd1 vccd1 _19146_/X sky130_fd_sc_hd__buf_8
XFILLER_0_143_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15309_ _15827_/A _15327_/A _15308_/X vssd1 vssd1 vccd1 vccd1 _15311_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16289_ _16287_/B _16309_/A _16288_/Y vssd1 vssd1 vccd1 vccd1 _16289_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19077_ _19077_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _19077_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18028_ _18028_/A _18028_/B vssd1 vssd1 vccd1 vccd1 _22218_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_112_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19979_ _26275_/Q _19134_/X hold806/X vssd1 vssd1 vccd1 vccd1 _19980_/C sky130_fd_sc_hd__a21o_1
X_22990_ _23138_/A vssd1 vssd1 vccd1 vccd1 _22991_/A sky130_fd_sc_hd__inv_2
X_21941_ _19388_/A _21940_/A _21940_/Y vssd1 vssd1 vccd1 vccd1 _21943_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24660_ _24660_/A vssd1 vssd1 vccd1 vccd1 _26282_/D sky130_fd_sc_hd__clkbuf_1
X_21872_ _19359_/A _21871_/A _21871_/Y vssd1 vssd1 vccd1 vccd1 _21874_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23611_ _23611_/A _23629_/B vssd1 vssd1 vccd1 vccd1 _23612_/A sky130_fd_sc_hd__and2_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20823_ _20825_/B _20825_/C vssd1 vssd1 vccd1 vccd1 _20824_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_128_clk clkbuf_4_14__f_clk/X vssd1 vssd1 vccd1 vccd1 _26335_/CLK sky130_fd_sc_hd__clkbuf_16
X_24591_ _26259_/Q hold2739/X _24664_/S vssd1 vssd1 vccd1 vccd1 _24591_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26330_ _26330_/CLK _26330_/D vssd1 vssd1 vccd1 vccd1 _26330_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23542_ _23539_/Y _23541_/Y _24858_/S vssd1 vssd1 vccd1 vccd1 _23542_/X sky130_fd_sc_hd__mux2_1
X_20754_ _20754_/A _25896_/Q vssd1 vssd1 vccd1 vccd1 _20759_/B sky130_fd_sc_hd__nand2_1
X_26261_ _26273_/CLK _26261_/D vssd1 vssd1 vccd1 vccd1 _26261_/Q sky130_fd_sc_hd__dfxtp_2
X_23473_ _24956_/S hold194/A _23472_/X vssd1 vssd1 vccd1 vccd1 _23473_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20685_ _21644_/B _21371_/B vssd1 vssd1 vccd1 vccd1 _20686_/B sky130_fd_sc_hd__nand2_1
X_25212_ _26292_/CLK hold720/X vssd1 vssd1 vccd1 vccd1 hold718/A sky130_fd_sc_hd__dfxtp_1
X_22424_ _25540_/Q _22424_/B vssd1 vssd1 vccd1 vccd1 _22424_/X sky130_fd_sc_hd__or2_1
XFILLER_0_45_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26192_ _26193_/CLK _26192_/D vssd1 vssd1 vccd1 vccd1 _26192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25143_ _26234_/CLK hold583/X vssd1 vssd1 vccd1 vccd1 hold581/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22355_ _22941_/B vssd1 vssd1 vccd1 vccd1 _22940_/B sky130_fd_sc_hd__inv_2
XFILLER_0_115_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21306_ _21306_/A _21306_/B vssd1 vssd1 vccd1 vccd1 _21308_/A sky130_fd_sc_hd__nand2_1
X_25074_ _26248_/CLK _25074_/D vssd1 vssd1 vccd1 vccd1 _25074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22286_ _22287_/A _22287_/B _23170_/A vssd1 vssd1 vccd1 vccd1 _22286_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24025_ _24025_/A vssd1 vssd1 vccd1 vccd1 _26076_/D sky130_fd_sc_hd__clkbuf_1
X_21237_ _21237_/A _22015_/B vssd1 vssd1 vccd1 vccd1 _21238_/A sky130_fd_sc_hd__nand2_1
Xhold260 hold260/A vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 hold271/A vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 hold282/A vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 hold293/A vssd1 vssd1 vccd1 vccd1 hold293/X sky130_fd_sc_hd__dlygate4sd3_1
X_21168_ _21627_/C _21580_/B vssd1 vssd1 vccd1 vccd1 _21169_/B sky130_fd_sc_hd__nand2_1
X_20119_ _21709_/A _21402_/A vssd1 vssd1 vccd1 vccd1 _20120_/C sky130_fd_sc_hd__nand2_1
X_25976_ _26040_/CLK _25976_/D vssd1 vssd1 vccd1 vccd1 _25976_/Q sky130_fd_sc_hd__dfxtp_1
X_13990_ _17909_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13990_/Y sky130_fd_sc_hd__nor2_1
X_21099_ _21099_/A vssd1 vssd1 vccd1 vccd1 _21099_/X sky130_fd_sc_hd__buf_6
XFILLER_0_102_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24927_ _24946_/A _24924_/X _24958_/B _24926_/Y vssd1 vssd1 vccd1 vccd1 _24927_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12941_ _26250_/Q _25619_/Q vssd1 vssd1 vccd1 vccd1 _14403_/A sky130_fd_sc_hd__xor2_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15660_ _15615_/X _15693_/B _15693_/C _15659_/X vssd1 vssd1 vccd1 vccd1 _15662_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24858_ _24856_/X _24857_/X _24858_/S vssd1 vssd1 vccd1 vccd1 _24858_/X sky130_fd_sc_hd__mux2_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _12726_/B _14364_/A _12752_/X _25606_/Q vssd1 vssd1 vccd1 vccd1 _12872_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14611_ _14611_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14611_/Y sky130_fd_sc_hd__nand2_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23809_ hold2123/X hold2036/X _23831_/S vssd1 vssd1 vccd1 vccd1 _23810_/A sky130_fd_sc_hd__mux2_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15591_ _15579_/X _15612_/A _15233_/X vssd1 vssd1 vccd1 vccd1 _15591_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_clk clkbuf_4_14__f_clk/X vssd1 vssd1 vccd1 vccd1 _26200_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24789_ _24789_/A vssd1 vssd1 vccd1 vccd1 _26324_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17330_ _17527_/A _17578_/A vssd1 vssd1 vccd1 vccd1 _17331_/B sky130_fd_sc_hd__xnor2_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _14542_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14542_/Y sky130_fd_sc_hd__nand2_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _25607_/Q vssd1 vssd1 vccd1 vccd1 _20936_/B sky130_fd_sc_hd__inv_2
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14473_ _14473_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14473_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16212_ _16212_/A hold912/X vssd1 vssd1 vccd1 vccd1 _16212_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19000_ _19000_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _19000_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_102_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13424_ _19033_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13424_/X sky130_fd_sc_hd__or2_1
X_17192_ _25602_/Q vssd1 vssd1 vccd1 vccd1 _20780_/B sky130_fd_sc_hd__inv_2
XFILLER_0_102_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16143_ _16132_/Y _16135_/Y _16156_/A _16142_/Y vssd1 vssd1 vccd1 vccd1 _16143_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13355_ _13220_/X _14632_/A _13242_/X _19673_/A vssd1 vssd1 vccd1 vccd1 _13355_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16074_ _16072_/X _16073_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _16074_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_122_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13286_ _26183_/Q _13239_/X _13285_/X vssd1 vssd1 vccd1 vccd1 _13286_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_87_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15025_ _15023_/X hold1953/X _14928_/X vssd1 vssd1 vccd1 vccd1 _15025_/Y sky130_fd_sc_hd__a21oi_1
X_19902_ _19900_/X _19901_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19902_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19833_ _19849_/B _19914_/B vssd1 vssd1 vccd1 vccd1 _19835_/A sky130_fd_sc_hd__xnor2_1
X_19764_ _21789_/A vssd1 vssd1 vccd1 vccd1 _19764_/X sky130_fd_sc_hd__buf_8
X_16976_ _16976_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16976_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_78_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18715_ _20487_/B _22410_/A vssd1 vssd1 vccd1 vccd1 _20478_/A sky130_fd_sc_hd__nand2_2
X_15927_ _15956_/A hold551/X vssd1 vssd1 vccd1 vccd1 hold552/A sky130_fd_sc_hd__nand2_1
Xinput6 io_in[5] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
X_19695_ _19723_/A _19695_/B vssd1 vssd1 vccd1 vccd1 _19695_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18646_ _18646_/A _18646_/B vssd1 vssd1 vccd1 vccd1 _22347_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_189_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ _15869_/A _15859_/A vssd1 vssd1 vccd1 vccd1 _15858_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14809_ _14809_/A vssd1 vssd1 vccd1 vccd1 _14996_/A sky130_fd_sc_hd__inv_2
XFILLER_0_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18577_ _19026_/A _18577_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18577_/X sky130_fd_sc_hd__and3_1
X_15789_ _15789_/A _15789_/B vssd1 vssd1 vccd1 vccd1 _15789_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_148_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17528_ _22704_/A vssd1 vssd1 vccd1 vccd1 _17528_/X sky130_fd_sc_hd__buf_12
XFILLER_0_15_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17459_ _17459_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17459_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_89_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20470_ _20470_/A _25850_/Q vssd1 vssd1 vccd1 vccd1 _20475_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19129_ _26215_/Q hold715/A vssd1 vssd1 vccd1 vccd1 _19129_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22140_ _22138_/X _22139_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _22140_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22071_ _22071_/A _22071_/B vssd1 vssd1 vccd1 vccd1 _22774_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_125_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21022_ _21022_/A _21022_/B vssd1 vssd1 vccd1 vccd1 _21025_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_10_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25830_ _25838_/CLK _25830_/D vssd1 vssd1 vccd1 vccd1 _25830_/Q sky130_fd_sc_hd__dfxtp_4
X_25761_ _25761_/CLK _25761_/D vssd1 vssd1 vccd1 vccd1 _25761_/Q sky130_fd_sc_hd__dfxtp_1
X_22973_ _23122_/A vssd1 vssd1 vccd1 vccd1 _22974_/A sky130_fd_sc_hd__inv_2
X_24712_ _24712_/A vssd1 vssd1 vccd1 vccd1 _26299_/D sky130_fd_sc_hd__clkbuf_1
X_21924_ _21924_/A _21924_/B vssd1 vssd1 vccd1 vccd1 _21926_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_97_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25692_ _26325_/CLK _25692_/D vssd1 vssd1 vccd1 vccd1 _25692_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24643_ _24643_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24644_/A sky130_fd_sc_hd__and2_1
XFILLER_0_167_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21855_ _21855_/A _21855_/B vssd1 vssd1 vccd1 vccd1 _21857_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_132_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20806_ _20806_/A _21371_/B _20806_/C vssd1 vssd1 vccd1 vccd1 _20807_/B sky130_fd_sc_hd__nand3_1
X_24574_ _24574_/A vssd1 vssd1 vccd1 vccd1 _26254_/D sky130_fd_sc_hd__clkbuf_1
X_21786_ _21786_/A _21786_/B vssd1 vssd1 vccd1 vccd1 _22909_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_148_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26313_ _26313_/CLK _26313_/D vssd1 vssd1 vccd1 vccd1 _26313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23525_ hold119/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23525_/X sky130_fd_sc_hd__or2b_1
X_20737_ _20737_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _20737_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26244_ _26244_/CLK _26244_/D vssd1 vssd1 vccd1 vccd1 _26244_/Q sky130_fd_sc_hd__dfxtp_2
X_23456_ _23450_/X _23455_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _23456_/X sky130_fd_sc_hd__mux2_1
X_20668_ _20668_/A _20668_/B vssd1 vssd1 vccd1 vccd1 _20670_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22407_ _22407_/A _25889_/Q vssd1 vssd1 vccd1 vccd1 _22407_/Y sky130_fd_sc_hd__nand2_1
X_26175_ _26175_/CLK _26175_/D vssd1 vssd1 vccd1 vccd1 _26175_/Q sky130_fd_sc_hd__dfxtp_1
X_23387_ _24942_/S hold101/A _23386_/X vssd1 vssd1 vccd1 vccd1 _23387_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20599_ _20599_/A _25892_/Q vssd1 vssd1 vccd1 vccd1 _20605_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25126_ _26335_/CLK _25126_/D vssd1 vssd1 vccd1 vccd1 _25126_/Q sky130_fd_sc_hd__dfxtp_1
X_13140_ _13109_/X _13137_/X _13096_/X _13139_/X vssd1 vssd1 vccd1 vccd1 _13140_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22338_ _22338_/A _23055_/A _22338_/C vssd1 vssd1 vccd1 vccd1 _22338_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_115_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25057_ _26142_/CLK _25057_/D vssd1 vssd1 vccd1 vccd1 _25057_/Q sky130_fd_sc_hd__dfxtp_1
X_13071_ _13018_/X _13069_/X _13005_/X _13070_/X vssd1 vssd1 vccd1 vccd1 _13071_/X
+ sky130_fd_sc_hd__o211a_1
X_22269_ _22269_/A _22269_/B vssd1 vssd1 vccd1 vccd1 _22269_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24008_ hold2430/X hold2425/X _24047_/S vssd1 vssd1 vccd1 vccd1 _24009_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16830_ _16831_/B _16831_/A vssd1 vssd1 vccd1 vccd1 _16830_/X sky130_fd_sc_hd__or2_1
X_16761_ _16761_/A _16761_/B vssd1 vssd1 vccd1 vccd1 _16761_/Y sky130_fd_sc_hd__nand2_1
X_13973_ hold639/X _13972_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold640/A sky130_fd_sc_hd__a21oi_1
X_25959_ _26023_/CLK _25959_/D vssd1 vssd1 vccd1 vccd1 _25959_/Q sky130_fd_sc_hd__dfxtp_1
X_18500_ _19616_/A vssd1 vssd1 vccd1 vccd1 _22149_/B sky130_fd_sc_hd__inv_2
X_15712_ _16937_/A _15712_/B vssd1 vssd1 vccd1 vccd1 _15713_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_38_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12924_ _12840_/X _12922_/X _12917_/X _12923_/X vssd1 vssd1 vccd1 vccd1 _12924_/X
+ sky130_fd_sc_hd__o211a_1
X_16692_ _16692_/A _16692_/B vssd1 vssd1 vccd1 vccd1 _16695_/C sky130_fd_sc_hd__xor2_1
X_19480_ _19472_/X _19479_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19480_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18431_ _21270_/B _22042_/A vssd1 vssd1 vccd1 vccd1 _21264_/A sky130_fd_sc_hd__nand2_2
X_15643_ _15615_/X _15693_/B _15626_/B vssd1 vssd1 vccd1 vccd1 _15645_/A sky130_fd_sc_hd__a21o_1
X_12855_ _12840_/X _12853_/X _12827_/X _12854_/X vssd1 vssd1 vccd1 vccd1 _12855_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15574_ _15577_/A _15575_/A vssd1 vssd1 vccd1 vccd1 _15574_/X sky130_fd_sc_hd__or2_1
XFILLER_0_111_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18362_ _25872_/Q _21946_/A vssd1 vssd1 vccd1 vccd1 _18370_/A sky130_fd_sc_hd__or2_2
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _17122_/B _14264_/A vssd1 vssd1 vccd1 vccd1 _12786_/X sky130_fd_sc_hd__or2_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17313_ _17311_/Y _17312_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _25603_/D sky130_fd_sc_hd__a21oi_1
X_14525_ _14525_/A hold131/X vssd1 vssd1 vccd1 vccd1 hold132/A sky130_fd_sc_hd__nand2_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18293_ _18535_/A _18293_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _18293_/X sky130_fd_sc_hd__and3_1
XFILLER_0_56_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17244_ _21791_/A vssd1 vssd1 vccd1 vccd1 _17444_/B sky130_fd_sc_hd__clkbuf_8
X_14456_ _14465_/A hold53/X vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__nand2_1
XFILLER_0_114_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13407_ _13407_/A vssd1 vssd1 vccd1 vccd1 _19802_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17175_ _17173_/X _23187_/B _17174_/X vssd1 vssd1 vccd1 vccd1 _17176_/A sky130_fd_sc_hd__a21o_1
X_14387_ _14385_/Y hold327/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold328/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16126_ _16134_/B _16127_/A vssd1 vssd1 vccd1 vccd1 _16126_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13338_ _26191_/Q _13239_/X _13337_/X vssd1 vssd1 vccd1 vccd1 _13338_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_84_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16057_ _16040_/B _16052_/B _16039_/A vssd1 vssd1 vccd1 vccd1 _16057_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13269_ _18658_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13269_/X sky130_fd_sc_hd__or2_1
X_15008_ _15003_/A _14997_/A _14997_/B vssd1 vssd1 vccd1 vccd1 _15010_/A sky130_fd_sc_hd__a21bo_1
Xhold2408 _15312_/Y vssd1 vssd1 vccd1 vccd1 _25446_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2419 _24977_/Q vssd1 vssd1 vccd1 vccd1 _12616_/A sky130_fd_sc_hd__dlygate4sd3_1
X_19816_ _19816_/A _20635_/B vssd1 vssd1 vccd1 vccd1 _19816_/Y sky130_fd_sc_hd__nor2_1
Xhold1707 _22857_/Y vssd1 vssd1 vccd1 vccd1 _25880_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1718 _21397_/Y vssd1 vssd1 vccd1 vccd1 _25817_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1729 _17205_/Y vssd1 vssd1 vccd1 vccd1 _25595_/D sky130_fd_sc_hd__dlygate4sd3_1
X_19747_ _19763_/B _19835_/B vssd1 vssd1 vccd1 vccd1 _19749_/A sky130_fd_sc_hd__xnor2_1
X_16959_ _16960_/B _16960_/A vssd1 vssd1 vccd1 vccd1 _16959_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19678_ _19678_/A _19678_/B vssd1 vssd1 vccd1 vccd1 _19678_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_154_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18629_ _18952_/A _25757_/Q _18891_/C vssd1 vssd1 vccd1 vccd1 _18630_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_176_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21640_ _21638_/Y _21639_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21640_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_164_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21571_ _21571_/A _21571_/B vssd1 vssd1 vccd1 vccd1 _21572_/A sky130_fd_sc_hd__nand2_1
XANTENNA_11 _23457_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _17863_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23310_ _23310_/A _23310_/B vssd1 vssd1 vccd1 vccd1 _23310_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20522_ _20522_/A _22441_/B _20522_/C vssd1 vssd1 vccd1 vccd1 _20526_/C sky130_fd_sc_hd__nand3_1
XANTENNA_33 _25837_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_44 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_24290_ hold2166/X hold1949/X _24356_/S vssd1 vssd1 vccd1 vccd1 _24291_/A sky130_fd_sc_hd__mux2_1
XANTENNA_55 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_66 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23241_ _23242_/A _23243_/A vssd1 vssd1 vccd1 vccd1 _23241_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_77 _25581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20453_ _21252_/B _21546_/A vssd1 vssd1 vccd1 vccd1 _20455_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_104_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23172_ _23188_/A _23172_/B vssd1 vssd1 vccd1 vccd1 _23172_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20384_ _21042_/A _20384_/B _20383_/X vssd1 vssd1 vccd1 vccd1 _20385_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22123_ _19602_/A _22122_/A _22122_/Y vssd1 vssd1 vccd1 vccd1 _22125_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22054_ _22055_/A _22055_/C _23042_/A vssd1 vssd1 vccd1 vccd1 _22054_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_11_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21005_ _21529_/C vssd1 vssd1 vccd1 vccd1 _21532_/B sky130_fd_sc_hd__inv_2
X_25813_ _25835_/CLK _25813_/D vssd1 vssd1 vccd1 vccd1 _25813_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_98_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25744_ _25781_/CLK _25744_/D vssd1 vssd1 vccd1 vccd1 _25744_/Q sky130_fd_sc_hd__dfxtp_1
X_22956_ _23106_/A vssd1 vssd1 vccd1 vccd1 _22957_/A sky130_fd_sc_hd__inv_2
XFILLER_0_186_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21907_ _19373_/A _21906_/A _21906_/Y vssd1 vssd1 vccd1 vccd1 _21909_/A sky130_fd_sc_hd__o21ai_1
X_25675_ _26306_/CLK _25675_/D vssd1 vssd1 vccd1 vccd1 _25675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22887_ _22878_/Y _22886_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22887_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_70_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12640_ _12640_/A _24836_/B _12640_/C vssd1 vssd1 vccd1 vccd1 _12640_/X sky130_fd_sc_hd__and3_1
X_24626_ _24626_/A vssd1 vssd1 vccd1 vccd1 _26271_/D sky130_fd_sc_hd__clkbuf_1
X_21838_ _19345_/A _21837_/A _21837_/Y vssd1 vssd1 vccd1 vccd1 _21840_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_183_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12571_ _12574_/A _24836_/B _12571_/C vssd1 vssd1 vccd1 vccd1 _12572_/A sky130_fd_sc_hd__and3_1
X_24557_ _24557_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24558_/A sky130_fd_sc_hd__and2_1
X_21769_ _21769_/A _21769_/B vssd1 vssd1 vccd1 vccd1 _21770_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_109_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_50_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _26014_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_148_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14310_ _14310_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14310_/Y sky130_fd_sc_hd__nand2_1
X_23508_ _23496_/X _23507_/X _24949_/S vssd1 vssd1 vccd1 vccd1 _23508_/X sky130_fd_sc_hd__mux2_1
X_15290_ _15290_/A _15290_/B vssd1 vssd1 vccd1 vccd1 _15290_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_124_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24488_ _24488_/A vssd1 vssd1 vccd1 vccd1 _26226_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_1231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14241_ hold633/X _14240_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold634/A sky130_fd_sc_hd__a21oi_1
X_26227_ _26232_/CLK _26227_/D vssd1 vssd1 vccd1 vccd1 _26227_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_124_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23439_ _23434_/Y _23437_/Y _24957_/S vssd1 vssd1 vccd1 vccd1 _23439_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26158_ _26244_/CLK _26158_/D vssd1 vssd1 vccd1 vccd1 _26158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14172_ _18653_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14172_/Y sky130_fd_sc_hd__nor2_1
X_13123_ _18144_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13123_/X sky130_fd_sc_hd__or2_1
X_25109_ _26193_/CLK _25109_/D vssd1 vssd1 vccd1 vccd1 _25109_/Q sky130_fd_sc_hd__dfxtp_1
X_18980_ _18978_/Y _18979_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25694_/D sky130_fd_sc_hd__a21oi_1
X_26089_ _26089_/CLK _26089_/D vssd1 vssd1 vccd1 vccd1 _26089_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17931_ _17931_/A _17931_/B vssd1 vssd1 vccd1 vccd1 _17932_/B sky130_fd_sc_hd__nand2_1
X_13054_ _13018_/X _13052_/X _13005_/X _13053_/X vssd1 vssd1 vccd1 vccd1 _13054_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17862_ _18392_/A _19045_/B vssd1 vssd1 vccd1 vccd1 _17863_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19601_ _19598_/Y _19601_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19601_/X sky130_fd_sc_hd__and3b_1
X_16813_ _16858_/A _16813_/B vssd1 vssd1 vccd1 vccd1 _16813_/Y sky130_fd_sc_hd__nand2_1
X_17793_ _18100_/A vssd1 vssd1 vccd1 vccd1 _18612_/A sky130_fd_sc_hd__buf_8
X_19532_ _19532_/A _21211_/B vssd1 vssd1 vccd1 vccd1 _19532_/Y sky130_fd_sc_hd__nor2_1
X_16744_ _16742_/Y _16743_/Y _16594_/X vssd1 vssd1 vccd1 vccd1 _16744_/Y sky130_fd_sc_hd__a21oi_1
X_13956_ _14000_/A hold777/X vssd1 vssd1 vccd1 vccd1 hold778/A sky130_fd_sc_hd__nand2_1
XFILLER_0_159_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12907_ _14262_/B vssd1 vssd1 vccd1 vccd1 _12907_/X sky130_fd_sc_hd__buf_12
X_19463_ _19463_/A _19463_/B vssd1 vssd1 vccd1 vccd1 _19463_/Y sky130_fd_sc_hd__nand2_1
X_16675_ hold608/X vssd1 vssd1 vccd1 vccd1 _16678_/B sky130_fd_sc_hd__inv_2
XFILLER_0_158_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13887_ _14125_/A vssd1 vssd1 vccd1 vccd1 _14000_/A sky130_fd_sc_hd__buf_8
XFILLER_0_158_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18414_ _22786_/A vssd1 vssd1 vccd1 vccd1 _18976_/C sky130_fd_sc_hd__clkbuf_8
X_15626_ _15626_/A _15626_/B vssd1 vssd1 vccd1 vccd1 _15693_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12838_ _17256_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12838_/X sky130_fd_sc_hd__or2_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19394_ _19392_/X _19393_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19394_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18345_ _18345_/A _25807_/Q _18345_/C vssd1 vssd1 vccd1 vccd1 _21164_/C sky130_fd_sc_hd__nand3_2
X_15557_ _15557_/A _15557_/B vssd1 vssd1 vccd1 vccd1 _15557_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_139_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12769_ _12726_/B _14301_/A _12752_/X _25586_/Q vssd1 vssd1 vccd1 vccd1 _12769_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_41_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _26041_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14508_ _14506_/Y hold21/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__a21oi_1
X_15488_ _26026_/Q _25962_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15489_/A sky130_fd_sc_hd__mux2_1
X_18276_ _19458_/A vssd1 vssd1 vccd1 vccd1 _21810_/B sky130_fd_sc_hd__inv_2
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17227_ _17393_/A _17227_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17227_/X sky130_fd_sc_hd__and3_1
X_14439_ _14437_/Y hold123/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold124/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17158_ _19758_/A _17158_/B vssd1 vssd1 vccd1 vccd1 _17562_/A sky130_fd_sc_hd__xor2_4
Xhold804 hold804/A vssd1 vssd1 vccd1 vccd1 hold804/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold815 hold815/A vssd1 vssd1 vccd1 vccd1 hold815/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold826 hold826/A vssd1 vssd1 vccd1 vccd1 hold826/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 hold837/A vssd1 vssd1 vccd1 vccd1 hold837/X sky130_fd_sc_hd__dlygate4sd3_1
X_16109_ _16109_/A vssd1 vssd1 vccd1 vccd1 _16133_/B sky130_fd_sc_hd__inv_2
Xhold848 hold848/A vssd1 vssd1 vccd1 vccd1 hold848/X sky130_fd_sc_hd__dlygate4sd3_1
X_17089_ _20273_/B _25884_/Q _25820_/Q vssd1 vssd1 vccd1 vccd1 _17090_/B sky130_fd_sc_hd__mux2_2
Xhold859 hold859/A vssd1 vssd1 vccd1 vccd1 hold859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2205 _14943_/Y vssd1 vssd1 vccd1 vccd1 _25417_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2216 _25996_/Q vssd1 vssd1 vccd1 vccd1 hold2216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2227 _24982_/Q vssd1 vssd1 vccd1 vccd1 _12654_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2238 _26016_/Q vssd1 vssd1 vccd1 vccd1 hold2238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2249 _26144_/Q vssd1 vssd1 vccd1 vccd1 hold2249/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1504 _13321_/X vssd1 vssd1 vccd1 vccd1 _25105_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1515 _25114_/Q vssd1 vssd1 vccd1 vccd1 _18976_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1526 _20881_/Y vssd1 vssd1 vccd1 vccd1 _25796_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1537 _25777_/Q vssd1 vssd1 vccd1 vccd1 _20160_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1548 _17300_/Y vssd1 vssd1 vccd1 vccd1 _25602_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1559 _25117_/Q vssd1 vssd1 vccd1 vccd1 _18998_/B sky130_fd_sc_hd__dlygate4sd3_1
X_22810_ _22960_/A _22810_/B vssd1 vssd1 vccd1 vccd1 _22811_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23790_ _23790_/A vssd1 vssd1 vccd1 vccd1 _26001_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22741_ _22739_/X _22740_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22741_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_177_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25460_ _26009_/CLK _25460_/D vssd1 vssd1 vccd1 vccd1 _25460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22672_ _23152_/B vssd1 vssd1 vccd1 vccd1 _23151_/B sky130_fd_sc_hd__inv_2
XFILLER_0_176_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xascon_wrapper_17 vssd1 vssd1 vccd1 vccd1 io_oeb[3] ascon_wrapper_17/LO sky130_fd_sc_hd__conb_1
X_24411_ _24411_/A vssd1 vssd1 vccd1 vccd1 _26201_/D sky130_fd_sc_hd__clkbuf_1
X_21623_ _22058_/A _21623_/B vssd1 vssd1 vccd1 vccd1 _21623_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25391_ _26004_/CLK _25391_/D vssd1 vssd1 vccd1 vccd1 _25391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _25893_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24342_ _24342_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24343_/A sky130_fd_sc_hd__and2_1
X_21554_ _21636_/A _21554_/B _21553_/X vssd1 vssd1 vccd1 vccd1 _21555_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_7_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20505_ _20503_/Y _20504_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _20505_/Y sky130_fd_sc_hd__a21oi_1
X_24273_ hold2182/X hold1985/X _24279_/S vssd1 vssd1 vccd1 vccd1 _24274_/A sky130_fd_sc_hd__mux2_1
X_21485_ _21485_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21490_/A sky130_fd_sc_hd__nand2_1
X_26012_ _26012_/CLK _26012_/D vssd1 vssd1 vccd1 vccd1 _26012_/Q sky130_fd_sc_hd__dfxtp_1
X_23224_ _23240_/A vssd1 vssd1 vccd1 vccd1 _23231_/A sky130_fd_sc_hd__inv_2
XFILLER_0_133_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20436_ _20436_/A _20436_/B vssd1 vssd1 vccd1 vccd1 _21249_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23155_ _23155_/A _23187_/B vssd1 vssd1 vccd1 vccd1 _23155_/Y sky130_fd_sc_hd__nand2_1
X_20367_ _20370_/A _20370_/C vssd1 vssd1 vccd1 vccd1 _20369_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22106_ _22106_/A _22106_/B vssd1 vssd1 vccd1 vccd1 _22108_/A sky130_fd_sc_hd__xor2_4
X_23086_ _23084_/X _23085_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _23086_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20298_ _20298_/A _20298_/B _21059_/C vssd1 vssd1 vccd1 vccd1 _20299_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_101_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_99_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _25495_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22037_ _22035_/X _15839_/B _22036_/Y _14786_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _22038_/A sky130_fd_sc_hd__a32o_1
Xhold2750 _25907_/Q vssd1 vssd1 vccd1 vccd1 _14694_/A sky130_fd_sc_hd__dlygate4sd3_1
X_13810_ _26267_/Q _13801_/X _13793_/X _13809_/Y vssd1 vssd1 vccd1 vccd1 _13811_/B
+ sky130_fd_sc_hd__a22o_1
X_14790_ _22060_/B _15778_/B vssd1 vssd1 vccd1 vccd1 _14791_/A sky130_fd_sc_hd__nand2_1
X_23988_ _23988_/A vssd1 vssd1 vccd1 vccd1 _26064_/D sky130_fd_sc_hd__clkbuf_1
X_13741_ hold366/X _13740_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold367/A sky130_fd_sc_hd__a21oi_1
X_22939_ _23090_/A vssd1 vssd1 vccd1 vccd1 _22940_/A sky130_fd_sc_hd__inv_2
X_25727_ _25727_/CLK _25727_/D vssd1 vssd1 vccd1 vccd1 _25727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16460_ _16461_/B _16438_/A _16452_/B vssd1 vssd1 vccd1 vccd1 _16468_/B sky130_fd_sc_hd__a21oi_1
X_13672_ _13703_/A _13672_/B vssd1 vssd1 vccd1 vccd1 _13672_/Y sky130_fd_sc_hd__nand2_1
X_25658_ _26289_/CLK _25658_/D vssd1 vssd1 vccd1 vccd1 _25658_/Q sky130_fd_sc_hd__dfxtp_1
X_15411_ _15411_/A _15411_/B vssd1 vssd1 vccd1 vccd1 _15553_/A sky130_fd_sc_hd__nand2_1
X_12623_ _12629_/A vssd1 vssd1 vccd1 vccd1 _12628_/A sky130_fd_sc_hd__inv_2
X_16391_ _16404_/B _16391_/B vssd1 vssd1 vccd1 vccd1 _16394_/B sky130_fd_sc_hd__and2_1
XFILLER_0_66_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24609_ hold2719/X hold2700/X _24664_/S vssd1 vssd1 vccd1 vccd1 _24610_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_109_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25589_ _26221_/CLK _25589_/D vssd1 vssd1 vccd1 vccd1 _25589_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_94_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_clk _25759_/CLK vssd1 vssd1 vccd1 vccd1 _26251_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_171_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15342_ _15342_/A _15342_/B vssd1 vssd1 vccd1 vccd1 _15406_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_136_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18130_ _21904_/B _25606_/Q vssd1 vssd1 vccd1 vccd1 _18132_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12554_ _23211_/A vssd1 vssd1 vccd1 vccd1 _16996_/C sky130_fd_sc_hd__inv_1
XFILLER_0_53_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15273_ _15266_/A _15232_/B _15248_/A vssd1 vssd1 vccd1 vccd1 _15273_/X sky130_fd_sc_hd__a21o_1
X_18061_ _18252_/A _19176_/A vssd1 vssd1 vccd1 vccd1 _18061_/Y sky130_fd_sc_hd__nand2_1
X_12485_ _14277_/A _14277_/B vssd1 vssd1 vccd1 vccd1 _23191_/C sky130_fd_sc_hd__nand2_8
XFILLER_0_81_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14224_ _14236_/A hold566/X vssd1 vssd1 vccd1 vccd1 hold567/A sky130_fd_sc_hd__nand2_1
X_17012_ _17012_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17012_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_184_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14155_ _14345_/A vssd1 vssd1 vccd1 vccd1 _14155_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ _26153_/Q _13065_/X _13105_/X vssd1 vssd1 vccd1 vccd1 _13106_/X sky130_fd_sc_hd__a21o_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14086_ _14180_/A _14086_/B vssd1 vssd1 vccd1 vccd1 _14086_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_95_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18963_ _18963_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18963_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_120_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17914_ _18535_/A _17914_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _17914_/X sky130_fd_sc_hd__and3_1
X_13037_ _17595_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13037_/X sky130_fd_sc_hd__or2_1
X_18894_ _18955_/A _18894_/B _18894_/C vssd1 vssd1 vccd1 vccd1 _18895_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17845_ _18528_/A _25728_/Q vssd1 vssd1 vccd1 vccd1 _17847_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_89_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17776_ _16996_/C _17764_/A _17794_/A vssd1 vssd1 vccd1 vccd1 _17779_/B sky130_fd_sc_hd__o21ai_1
X_14988_ _14989_/B _14989_/A vssd1 vssd1 vccd1 vccd1 _14990_/A sky130_fd_sc_hd__or2_1
X_19515_ _26241_/Q hold596/X vssd1 vssd1 vccd1 vccd1 _19515_/Y sky130_fd_sc_hd__nand2_1
X_16727_ _16725_/X _16711_/X _16726_/Y _25864_/Q _14170_/X vssd1 vssd1 vccd1 vccd1
+ _16728_/A sky130_fd_sc_hd__a32o_1
X_13939_ _17859_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13939_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_44_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19446_ _21047_/A _19444_/Y _21051_/C vssd1 vssd1 vccd1 vccd1 _19537_/B sky130_fd_sc_hd__o21a_2
X_16658_ _16658_/A _16658_/B vssd1 vssd1 vccd1 vccd1 _16681_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_159_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15609_ _15609_/A _15609_/B vssd1 vssd1 vccd1 vccd1 _15609_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_174_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19377_ _19378_/B _19378_/A vssd1 vssd1 vccd1 vccd1 _19377_/X sky130_fd_sc_hd__or2_1
X_16589_ _16555_/A _16597_/A _16577_/Y vssd1 vssd1 vccd1 vccd1 _16589_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _26148_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18328_ _18328_/A _18328_/B _18328_/C vssd1 vssd1 vccd1 vccd1 _21880_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18259_ _18445_/A _18263_/B vssd1 vssd1 vccd1 vccd1 _18261_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21270_ _21270_/A _21270_/B vssd1 vssd1 vccd1 vccd1 _21272_/A sky130_fd_sc_hd__nand2_1
Xhold601 hold601/A vssd1 vssd1 vccd1 vccd1 hold601/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold612 hold612/A vssd1 vssd1 vccd1 vccd1 hold612/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold623 hold623/A vssd1 vssd1 vccd1 vccd1 hold623/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20221_ _21450_/A _21086_/C vssd1 vssd1 vccd1 vccd1 _20224_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_130_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold634 hold634/A vssd1 vssd1 vccd1 vccd1 hold634/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold645 hold645/A vssd1 vssd1 vccd1 vccd1 hold645/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold656 hold656/A vssd1 vssd1 vccd1 vccd1 hold656/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_12_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold667 hold667/A vssd1 vssd1 vccd1 vccd1 hold667/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold678 hold678/A vssd1 vssd1 vccd1 vccd1 hold678/X sky130_fd_sc_hd__dlygate4sd3_1
X_20152_ _20152_/A _20152_/B vssd1 vssd1 vccd1 vccd1 _20153_/A sky130_fd_sc_hd__nand2_1
Xhold689 hold689/A vssd1 vssd1 vccd1 vccd1 hold689/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2002 _24213_/X vssd1 vssd1 vccd1 vccd1 _24214_/A sky130_fd_sc_hd__dlygate4sd3_1
X_24960_ _24954_/X _24958_/Y _24959_/X _23484_/B vssd1 vssd1 vccd1 vccd1 _24960_/X
+ sky130_fd_sc_hd__a31o_1
Xhold2013 _24981_/Q vssd1 vssd1 vccd1 vccd1 _12654_/C sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold2024 _23613_/X vssd1 vssd1 vccd1 vccd1 _23614_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20083_ _20083_/A _20083_/B vssd1 vssd1 vccd1 vccd1 _20084_/A sky130_fd_sc_hd__nand2_1
Xhold2035 _24111_/X vssd1 vssd1 vccd1 vccd1 _24112_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2046 _26121_/Q vssd1 vssd1 vccd1 vccd1 hold2046/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1301 _13033_/X vssd1 vssd1 vccd1 vccd1 _25056_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2057 _23352_/X vssd1 vssd1 vccd1 vccd1 _23353_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23911_ hold1912/X _26041_/Q _23920_/S vssd1 vssd1 vccd1 vccd1 _23911_/X sky130_fd_sc_hd__mux2_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1312 _25075_/Q vssd1 vssd1 vccd1 vccd1 _18208_/B sky130_fd_sc_hd__dlygate4sd3_1
X_24891_ _24958_/B _24883_/X _24885_/Y _24890_/X vssd1 vssd1 vccd1 vccd1 _24891_/X
+ sky130_fd_sc_hd__a31o_1
Xhold2068 _25955_/Q vssd1 vssd1 vccd1 vccd1 hold2068/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1323 _25015_/Q vssd1 vssd1 vccd1 vccd1 _17200_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1334 _14722_/Y vssd1 vssd1 vccd1 vccd1 _25391_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2079 _25978_/Q vssd1 vssd1 vccd1 vccd1 hold2079/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1345 _25800_/Q vssd1 vssd1 vccd1 vccd1 _20991_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23842_ _23842_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23843_/A sky130_fd_sc_hd__and2_1
Xhold1356 _19839_/Y vssd1 vssd1 vccd1 vccd1 _25760_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1367 _25050_/Q vssd1 vssd1 vccd1 vccd1 _17543_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1378 _14713_/Y vssd1 vssd1 vccd1 vccd1 _25390_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1389 _25017_/Q vssd1 vssd1 vccd1 vccd1 _17227_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23773_ _14824_/B _25996_/Q _23831_/S vssd1 vssd1 vccd1 vccd1 _23773_/X sky130_fd_sc_hd__mux2_1
X_20985_ _26303_/Q hold710/X vssd1 vssd1 vccd1 vccd1 _20985_/Y sky130_fd_sc_hd__nand2_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25512_ _25515_/CLK hold907/X vssd1 vssd1 vccd1 vccd1 hold906/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22724_ _22724_/A _22724_/B vssd1 vssd1 vccd1 vccd1 _23184_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_178_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25443_ _25501_/CLK _25443_/D vssd1 vssd1 vccd1 vccd1 _25443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22655_ _26053_/Q vssd1 vssd1 vccd1 vccd1 _22656_/A sky130_fd_sc_hd__inv_2
XFILLER_0_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21606_ _22058_/A _21606_/B vssd1 vssd1 vccd1 vccd1 _21606_/Y sky130_fd_sc_hd__nand2_1
X_25374_ _26200_/CLK hold154/X vssd1 vssd1 vccd1 vccd1 hold152/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22586_ _22586_/A vssd1 vssd1 vccd1 vccd1 _22937_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24325_ _24325_/A vssd1 vssd1 vccd1 vccd1 _26173_/D sky130_fd_sc_hd__clkbuf_1
X_21537_ _21536_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21537_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_168_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24256_ _24256_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24257_/A sky130_fd_sc_hd__and2_1
XFILLER_0_161_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21468_ _21468_/A _21468_/B vssd1 vssd1 vccd1 vccd1 _21469_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_160_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23207_ _23208_/B _23208_/A vssd1 vssd1 vccd1 vccd1 _23211_/B sky130_fd_sc_hd__nor2_1
X_20419_ _20419_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20424_/A sky130_fd_sc_hd__nand2_1
X_24187_ hold2159/X hold2189/X _24203_/S vssd1 vssd1 vccd1 vccd1 _24188_/A sky130_fd_sc_hd__mux2_1
X_21399_ _21449_/A _21402_/A vssd1 vssd1 vccd1 vccd1 _21400_/B sky130_fd_sc_hd__nand2_1
X_23138_ _23138_/A _23138_/B vssd1 vssd1 vccd1 vccd1 _23139_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_105_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15960_ _15960_/A _15960_/B vssd1 vssd1 vccd1 vccd1 _16000_/A sky130_fd_sc_hd__nand2_1
X_23069_ _23197_/A _23069_/B vssd1 vssd1 vccd1 vccd1 _23069_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_179_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14911_ _14911_/A vssd1 vssd1 vccd1 vccd1 _25413_/D sky130_fd_sc_hd__inv_2
XFILLER_0_41_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15891_ _15891_/A _15891_/B vssd1 vssd1 vccd1 vccd1 _15892_/B sky130_fd_sc_hd__nand2_1
Xhold2580 _26297_/Q vssd1 vssd1 vccd1 vccd1 hold2580/X sky130_fd_sc_hd__dlygate4sd3_1
X_17630_ _17630_/A _17630_/B vssd1 vssd1 vccd1 vccd1 _17630_/X sky130_fd_sc_hd__xor2_1
X_14842_ _14900_/A _14844_/A vssd1 vssd1 vccd1 vccd1 _14842_/Y sky130_fd_sc_hd__nand2_1
Xhold2591 _26286_/Q vssd1 vssd1 vccd1 vccd1 hold2591/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1890 _25704_/Q vssd1 vssd1 vccd1 vccd1 _19050_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17561_ _17559_/Y _17560_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _17561_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14773_ _14773_/A vssd1 vssd1 vccd1 vccd1 _14962_/A sky130_fd_sc_hd__inv_2
XFILLER_0_98_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19300_ _26226_/Q hold581/X vssd1 vssd1 vccd1 vccd1 _19300_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_105_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16512_ _16512_/A vssd1 vssd1 vccd1 vccd1 _16524_/B sky130_fd_sc_hd__inv_2
X_13724_ _13760_/A hold515/X vssd1 vssd1 vccd1 vccd1 hold516/A sky130_fd_sc_hd__nand2_1
X_17492_ _17492_/A _17492_/B vssd1 vssd1 vccd1 vccd1 _17492_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_39_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19231_ _20546_/A _22190_/B _25596_/Q vssd1 vssd1 vccd1 vccd1 _20551_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16443_ _16417_/Y _16439_/X _16442_/Y vssd1 vssd1 vccd1 vccd1 _16491_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_168_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13655_ hold417/X _13654_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold418/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12606_ _12606_/A _24836_/B _12606_/C vssd1 vssd1 vccd1 vccd1 _12606_/X sky130_fd_sc_hd__and3_1
X_19162_ _25655_/Q vssd1 vssd1 vccd1 vccd1 _22051_/A sky130_fd_sc_hd__inv_2
XFILLER_0_39_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16374_ _16374_/A _16374_/B _16378_/B vssd1 vssd1 vccd1 vccd1 _16374_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_184_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13586_ _13944_/A vssd1 vssd1 vccd1 vccd1 _13703_/A sky130_fd_sc_hd__buf_6
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18113_ _18109_/Y _18110_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25652_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15325_ _15323_/X hold2669/X _15090_/X vssd1 vssd1 vccd1 vccd1 _15325_/Y sky130_fd_sc_hd__a21oi_1
X_12537_ _23199_/C _12537_/B vssd1 vssd1 vccd1 vccd1 _12537_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_48_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19093_ _19093_/A _21784_/A vssd1 vssd1 vccd1 vccd1 _20067_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18044_ _18445_/A _18052_/B vssd1 vssd1 vccd1 vccd1 _18047_/A sky130_fd_sc_hd__nand2_1
X_15256_ _15256_/A _15810_/B vssd1 vssd1 vccd1 vccd1 _15257_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_2_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14207_ _25828_/Q vssd1 vssd1 vccd1 vccd1 _18774_/B sky130_fd_sc_hd__inv_2
XFILLER_0_112_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15187_ _15185_/B _15165_/B _15186_/Y vssd1 vssd1 vccd1 vccd1 _15272_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14138_ _14236_/A hold748/X vssd1 vssd1 vccd1 vccd1 hold749/A sky130_fd_sc_hd__nand2_1
X_19995_ _19990_/X _18879_/X _19994_/X vssd1 vssd1 vccd1 vccd1 _19996_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_120_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14069_ hold621/X _14068_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold622/A sky130_fd_sc_hd__a21oi_1
X_18946_ _25709_/Q _20088_/B vssd1 vssd1 vccd1 vccd1 _18949_/A sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_3_clk _26093_/CLK vssd1 vssd1 vccd1 vccd1 _25135_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18877_ _19003_/A _19052_/B vssd1 vssd1 vccd1 vccd1 _18878_/B sky130_fd_sc_hd__xnor2_1
X_17828_ _17828_/A _17828_/B _20069_/A vssd1 vssd1 vccd1 vccd1 _17836_/A sky130_fd_sc_hd__and3_2
XFILLER_0_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17759_ _17759_/A _17925_/B _17759_/C vssd1 vssd1 vccd1 vccd1 _17973_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_89_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20770_ _20770_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _20775_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_119_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19429_ _19426_/Y _19429_/B _19980_/B vssd1 vssd1 vccd1 vccd1 _19429_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_174_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22440_ _22441_/B _22441_/A vssd1 vssd1 vccd1 vccd1 _22442_/A sky130_fd_sc_hd__or2_1
XFILLER_0_17_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22371_ _18676_/A _25823_/Q _22369_/Y _22370_/Y vssd1 vssd1 vccd1 vccd1 _22372_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24110_ _24110_/A vssd1 vssd1 vccd1 vccd1 _26103_/D sky130_fd_sc_hd__clkbuf_1
X_21322_ _21322_/A _21322_/B _21322_/C vssd1 vssd1 vccd1 vccd1 _21323_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_142_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25090_ _26301_/CLK _25090_/D vssd1 vssd1 vccd1 vccd1 _25090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24041_ hold2523/X _26082_/Q _24047_/S vssd1 vssd1 vccd1 vccd1 _24041_/X sky130_fd_sc_hd__mux2_1
Xhold420 hold420/A vssd1 vssd1 vccd1 vccd1 hold420/X sky130_fd_sc_hd__dlygate4sd3_1
X_21253_ _21253_/A _21253_/B vssd1 vssd1 vccd1 vccd1 _21254_/A sky130_fd_sc_hd__nand2_1
Xhold431 hold431/A vssd1 vssd1 vccd1 vccd1 hold431/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 hold442/A vssd1 vssd1 vccd1 vccd1 hold442/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold453 hold453/A vssd1 vssd1 vccd1 vccd1 hold453/X sky130_fd_sc_hd__dlygate4sd3_1
X_20204_ _20204_/A _20204_/B _20204_/C vssd1 vssd1 vccd1 vccd1 _20208_/C sky130_fd_sc_hd__nand3_1
Xhold464 hold464/A vssd1 vssd1 vccd1 vccd1 hold464/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 hold475/A vssd1 vssd1 vccd1 vccd1 hold475/X sky130_fd_sc_hd__dlygate4sd3_1
X_21184_ _21184_/A _21184_/B vssd1 vssd1 vccd1 vccd1 _21187_/B sky130_fd_sc_hd__nand2_1
Xhold486 hold486/A vssd1 vssd1 vccd1 vccd1 hold486/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold497 hold497/A vssd1 vssd1 vccd1 vccd1 hold497/X sky130_fd_sc_hd__dlygate4sd3_1
X_20135_ _25880_/Q _20135_/B _20135_/C vssd1 vssd1 vccd1 vccd1 _20139_/B sky130_fd_sc_hd__nand3b_1
X_25992_ _25992_/CLK _25992_/D vssd1 vssd1 vccd1 vccd1 _25992_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24943_ _24957_/S _24943_/B vssd1 vssd1 vccd1 vccd1 _24943_/Y sky130_fd_sc_hd__nor2_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20066_ _21385_/A _21693_/A vssd1 vssd1 vccd1 vccd1 _20072_/B sky130_fd_sc_hd__nand2_1
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1120 _19468_/Y vssd1 vssd1 vccd1 vccd1 _25734_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 _25803_/Q vssd1 vssd1 vccd1 vccd1 _21072_/B sky130_fd_sc_hd__buf_1
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 _12850_/X vssd1 vssd1 vccd1 vccd1 _25021_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1153 _25749_/Q vssd1 vssd1 vccd1 vccd1 _19681_/B sky130_fd_sc_hd__dlygate4sd3_1
X_24874_ _16023_/B _16038_/B _24956_/S vssd1 vssd1 vccd1 vccd1 _24875_/A sky130_fd_sc_hd__mux2_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 _12896_/X vssd1 vssd1 vccd1 vccd1 _25030_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1175 _25574_/Q vssd1 vssd1 vccd1 vccd1 _16940_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 _13219_/X vssd1 vssd1 vccd1 vccd1 _25089_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23825_ hold2314/X hold2165/X _23831_/S vssd1 vssd1 vccd1 vccd1 _23826_/A sky130_fd_sc_hd__mux2_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1197 _25121_/Q vssd1 vssd1 vccd1 vccd1 _19026_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23756_ _23756_/A vssd1 vssd1 vccd1 vccd1 _25990_/D sky130_fd_sc_hd__clkbuf_1
X_20968_ _25864_/Q vssd1 vssd1 vccd1 vccd1 _21977_/B sky130_fd_sc_hd__inv_2
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22707_ _15300_/B _22680_/X _14273_/X vssd1 vssd1 vccd1 vccd1 _22707_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23687_ hold1974/X _25968_/Q _23754_/S vssd1 vssd1 vccd1 vccd1 _23687_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20899_ _20899_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _20904_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_95_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13440_ _26208_/Q _13426_/X _13439_/X vssd1 vssd1 vccd1 vccd1 _13440_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_36_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25426_ _25992_/CLK _25426_/D vssd1 vssd1 vccd1 vccd1 _25426_/Q sky130_fd_sc_hd__dfxtp_1
X_22638_ _22636_/X _22637_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22638_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13371_ _13371_/A vssd1 vssd1 vccd1 vccd1 _19715_/A sky130_fd_sc_hd__clkbuf_8
X_25357_ _26184_/CLK hold388/X vssd1 vssd1 vccd1 vccd1 hold386/A sky130_fd_sc_hd__dfxtp_1
X_22569_ _22569_/A _22569_/B vssd1 vssd1 vccd1 vccd1 _22570_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15110_ _15110_/A _15110_/B vssd1 vssd1 vccd1 vccd1 _15111_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_23_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16090_ _16212_/A hold763/X vssd1 vssd1 vccd1 vccd1 hold764/A sky130_fd_sc_hd__nand2_1
X_24308_ hold1920/X _26168_/Q _24356_/S vssd1 vssd1 vccd1 vccd1 _24308_/X sky130_fd_sc_hd__mux2_1
X_25288_ _26240_/CLK hold88/X vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15041_ _15042_/B _15042_/A vssd1 vssd1 vccd1 vccd1 _15043_/A sky130_fd_sc_hd__or2_1
XFILLER_0_160_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24239_ _24239_/A vssd1 vssd1 vccd1 vccd1 _26145_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18800_ _18798_/X _18269_/X _18799_/X vssd1 vssd1 vccd1 vccd1 _18801_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19780_ _19778_/X _19779_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19780_/Y sky130_fd_sc_hd__a21oi_1
X_16992_ _17402_/A _17491_/A vssd1 vssd1 vccd1 vccd1 _16993_/B sky130_fd_sc_hd__xnor2_1
X_18731_ _18731_/A _25826_/Q _18731_/C vssd1 vssd1 vccd1 vccd1 _20526_/B sky130_fd_sc_hd__nand3_2
X_15943_ _15934_/B _15940_/B _15933_/A vssd1 vssd1 vccd1 vccd1 _15943_/Y sky130_fd_sc_hd__o21ai_1
X_18662_ _18986_/A _19473_/A vssd1 vssd1 vccd1 vccd1 _18662_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ _15874_/A _15874_/B vssd1 vssd1 vccd1 vccd1 _15884_/B sky130_fd_sc_hd__nand2_1
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17613_ _18252_/A _17613_/B vssd1 vssd1 vccd1 vccd1 _17613_/Y sky130_fd_sc_hd__nand2_1
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ _14831_/B _22175_/A vssd1 vssd1 vccd1 vccd1 _22173_/B sky130_fd_sc_hd__xnor2_2
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18593_ _20244_/B _22269_/A vssd1 vssd1 vccd1 vccd1 _20235_/A sky130_fd_sc_hd__nand2_2
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17544_ _17542_/X _17528_/X _17543_/X vssd1 vssd1 vccd1 vccd1 _17545_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_54_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756_ _25844_/Q _12527_/A _14945_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14756_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13707_ _25748_/Q vssd1 vssd1 vccd1 vccd1 _18449_/B sky130_fd_sc_hd__inv_2
X_17475_ _17605_/A _17475_/B vssd1 vssd1 vccd1 vccd1 _17475_/Y sky130_fd_sc_hd__nand2_1
X_14687_ _14687_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _14687_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19214_ _19452_/A _19214_/B vssd1 vssd1 vccd1 vccd1 _19214_/Y sky130_fd_sc_hd__nand2_1
X_16426_ _16426_/A hold933/X vssd1 vssd1 vccd1 vccd1 _16442_/A sky130_fd_sc_hd__and2_1
XFILLER_0_172_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13638_ _18223_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13638_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19145_ _19145_/A _19961_/B vssd1 vssd1 vccd1 vccd1 _19145_/Y sky130_fd_sc_hd__nand2_1
X_16357_ _16358_/B _16358_/A vssd1 vssd1 vccd1 vccd1 _16374_/B sky130_fd_sc_hd__or2_1
XFILLER_0_82_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13569_ _18086_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13569_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_171_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15308_ _15264_/B _15290_/Y _15291_/A vssd1 vssd1 vccd1 vccd1 _15308_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19076_ _19074_/X _18879_/X _19075_/X vssd1 vssd1 vccd1 vccd1 _19077_/A sky130_fd_sc_hd__a21o_1
X_16288_ _16297_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16288_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_152_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18027_ _20586_/B _19244_/A vssd1 vssd1 vccd1 vccd1 _18028_/B sky130_fd_sc_hd__nand2_1
X_15239_ _16764_/B vssd1 vssd1 vccd1 vccd1 _22631_/B sky130_fd_sc_hd__inv_2
XFILLER_0_151_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19978_ _19977_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19980_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18929_ _18929_/A _18929_/B vssd1 vssd1 vccd1 vccd1 _22691_/A sky130_fd_sc_hd__or2_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21940_ _21940_/A _21940_/B vssd1 vssd1 vccd1 vccd1 _21940_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_55_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21871_ _21871_/A _21871_/B vssd1 vssd1 vccd1 vccd1 _21871_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23610_ hold2258/X hold2023/X _23677_/S vssd1 vssd1 vccd1 vccd1 _23611_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_89_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20822_ _20822_/A _21806_/B _20822_/C vssd1 vssd1 vccd1 vccd1 _20825_/C sky130_fd_sc_hd__nand3_1
X_24590_ _24743_/A vssd1 vssd1 vccd1 vccd1 _24664_/S sky130_fd_sc_hd__clkbuf_16
X_23541_ _24942_/S hold356/A _23540_/X vssd1 vssd1 vccd1 vccd1 _23541_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_159_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20753_ _20756_/A _20756_/C vssd1 vssd1 vccd1 vccd1 _20754_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26260_ _26273_/CLK _26260_/D vssd1 vssd1 vccd1 vccd1 _26260_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23472_ hold68/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23472_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20684_ _21645_/B vssd1 vssd1 vccd1 vccd1 _21644_/B sky130_fd_sc_hd__inv_2
XFILLER_0_135_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25211_ _26292_/CLK hold762/X vssd1 vssd1 vccd1 vccd1 hold760/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22423_ _22424_/B _22423_/B vssd1 vssd1 vccd1 vccd1 _22423_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_128_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26191_ _26193_/CLK _26191_/D vssd1 vssd1 vccd1 vccd1 _26191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25142_ _26234_/CLK hold421/X vssd1 vssd1 vccd1 vccd1 hold419/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22354_ _22354_/A _22354_/B vssd1 vssd1 vccd1 vccd1 _22941_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_66_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21305_ _21305_/A _21305_/B _21305_/C vssd1 vssd1 vccd1 vccd1 _21306_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_130_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25073_ _26284_/CLK _25073_/D vssd1 vssd1 vccd1 vccd1 _25073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22285_ _23023_/B vssd1 vssd1 vccd1 vccd1 _23170_/A sky130_fd_sc_hd__inv_2
X_24024_ _24024_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24025_/A sky130_fd_sc_hd__and2_1
XFILLER_0_131_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold250 hold250/A vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
X_21236_ _21234_/Y _21235_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21236_/Y sky130_fd_sc_hd__a21oi_1
Xhold261 hold261/A vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 hold272/A vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 hold283/A vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 hold294/A vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
X_21167_ _21630_/B vssd1 vssd1 vccd1 vccd1 _21627_/C sky130_fd_sc_hd__inv_2
XFILLER_0_141_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20118_ _21708_/A _21401_/A vssd1 vssd1 vccd1 vccd1 _20120_/A sky130_fd_sc_hd__nand2_1
X_25975_ _26079_/CLK _25975_/D vssd1 vssd1 vccd1 vccd1 _25975_/Q sky130_fd_sc_hd__dfxtp_1
X_21098_ _21235_/A _21098_/B vssd1 vssd1 vccd1 vccd1 _21098_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24926_ _24946_/A _24926_/B vssd1 vssd1 vccd1 vccd1 _24926_/Y sky130_fd_sc_hd__nor2_1
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20049_ _20051_/B _20051_/C vssd1 vssd1 vccd1 vccd1 _20050_/A sky130_fd_sc_hd__nand2_1
X_12940_ _12930_/X _12938_/X _12917_/X _12939_/X vssd1 vssd1 vccd1 vccd1 _12940_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24857_ _15515_/A _15530_/A _24863_/S vssd1 vssd1 vccd1 vccd1 _24857_/X sky130_fd_sc_hd__mux2_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _26237_/Q _25606_/Q vssd1 vssd1 vccd1 vccd1 _14364_/A sky130_fd_sc_hd__xor2_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _14608_/Y hold24/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__a21oi_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23808_ _23808_/A vssd1 vssd1 vccd1 vccd1 _26007_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _15590_/A _15590_/B vssd1 vssd1 vccd1 vccd1 _15612_/A sky130_fd_sc_hd__nor2_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24788_ _24788_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24789_/A sky130_fd_sc_hd__and2_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14541_ _14539_/Y hold96/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__a21oi_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23739_ _14723_/B _25985_/Q _23754_/S vssd1 vssd1 vccd1 vccd1 _23739_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17260_ _17258_/Y _17259_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _17260_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14472_ _14469_/Y hold192/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold193/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16211_ _16209_/X _16210_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _16211_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_181_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25409_ _26001_/CLK _25409_/D vssd1 vssd1 vccd1 vccd1 _25409_/Q sky130_fd_sc_hd__dfxtp_1
X_13423_ _26205_/Q _13239_/X _13422_/X vssd1 vssd1 vccd1 vccd1 _13423_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17191_ _17189_/Y _17190_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _17191_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16142_ _16150_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16142_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_183_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13354_ _26322_/Q _19673_/A vssd1 vssd1 vccd1 vccd1 _14632_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16073_ _16073_/A _16084_/B vssd1 vssd1 vccd1 vccd1 _16073_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_45_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13285_ _13220_/X _14599_/A _13242_/X _19518_/A vssd1 vssd1 vccd1 vccd1 _13285_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15024_ _15024_/A _15024_/B vssd1 vssd1 vccd1 vccd1 _15024_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_121_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19901_ _19901_/A _19901_/B vssd1 vssd1 vccd1 vccd1 _19901_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_20_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19832_ _20672_/A _19830_/Y _20677_/C vssd1 vssd1 vccd1 vccd1 _19914_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_20_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19763_ _19763_/A _19763_/B vssd1 vssd1 vccd1 vccd1 _19763_/Y sky130_fd_sc_hd__nand2_1
X_16975_ _16973_/X _16711_/A _16974_/Y _25900_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16976_/A sky130_fd_sc_hd__a32o_1
X_18714_ _18714_/A _18714_/B _18714_/C vssd1 vssd1 vccd1 vccd1 _22410_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_21_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15926_ _15926_/A _16697_/B _15934_/A vssd1 vssd1 vccd1 vccd1 _15926_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19694_ _19686_/X _19693_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19694_/Y sky130_fd_sc_hd__o21ai_1
Xinput7 rst vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_155_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18645_ _20362_/B _19715_/A vssd1 vssd1 vccd1 vccd1 _18646_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ _15857_/A _15857_/B vssd1 vssd1 vccd1 vccd1 _15859_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_91_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14808_ _22115_/B _15543_/B vssd1 vssd1 vccd1 vccd1 _14809_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18576_ _18576_/A _18576_/B vssd1 vssd1 vccd1 vccd1 _18576_/X sky130_fd_sc_hd__xor2_1
X_15788_ _15762_/A _15786_/A _15781_/A vssd1 vssd1 vccd1 vccd1 _15789_/B sky130_fd_sc_hd__o21a_1
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17527_ _17527_/A _17527_/B vssd1 vssd1 vccd1 vccd1 _17527_/X sky130_fd_sc_hd__xor2_1
X_14739_ _14739_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14739_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17458_ _17456_/X _17241_/X _17457_/X vssd1 vssd1 vccd1 vccd1 _17459_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_27_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16409_ _16407_/X _16408_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 hold967/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17389_ _21238_/B _25874_/Q _25810_/Q vssd1 vssd1 vccd1 vccd1 _17390_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_171_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19128_ _19126_/Y hold669/X _19086_/X vssd1 vssd1 vccd1 vccd1 hold670/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19059_ _19059_/A _19059_/B vssd1 vssd1 vccd1 vccd1 _19060_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22070_ _22070_/A _22789_/B vssd1 vssd1 vccd1 vccd1 _22071_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_11_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21021_ _21021_/A _21738_/B vssd1 vssd1 vccd1 vccd1 _21022_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22972_ _22970_/X _22971_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _22972_/Y sky130_fd_sc_hd__a21oi_1
X_25760_ _25898_/CLK _25760_/D vssd1 vssd1 vccd1 vccd1 _25760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24711_ _24711_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24712_/A sky130_fd_sc_hd__and2_1
X_21923_ _25843_/Q _25779_/Q vssd1 vssd1 vccd1 vccd1 _21924_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25691_ _26324_/CLK _25691_/D vssd1 vssd1 vccd1 vccd1 _25691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21854_ _25841_/Q _25777_/Q vssd1 vssd1 vccd1 vccd1 _21855_/B sky130_fd_sc_hd__nor2_2
X_24642_ hold2632/X _26277_/Q _24664_/S vssd1 vssd1 vccd1 vccd1 _24642_/X sky130_fd_sc_hd__mux2_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20805_ _21419_/B _21693_/B vssd1 vssd1 vccd1 vccd1 _20806_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_77_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24573_ _24573_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24574_/A sky130_fd_sc_hd__and2_1
XFILLER_0_93_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21785_ _17834_/B _17032_/B _17835_/B vssd1 vssd1 vccd1 vccd1 _21786_/B sky130_fd_sc_hd__o21ai_2
X_26312_ _26313_/CLK _26312_/D vssd1 vssd1 vccd1 vccd1 _26312_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_163_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20736_ _20736_/A _20736_/B vssd1 vssd1 vccd1 vccd1 _20737_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23524_ _23521_/Y _23523_/Y _24946_/A vssd1 vssd1 vccd1 vccd1 _23524_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26243_ _26244_/CLK _26243_/D vssd1 vssd1 vccd1 vccd1 _26243_/Q sky130_fd_sc_hd__dfxtp_2
X_23455_ _23452_/Y _23454_/Y _24946_/A vssd1 vssd1 vccd1 vccd1 _23455_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20667_ _20669_/B _20669_/C vssd1 vssd1 vccd1 vccd1 _20668_/A sky130_fd_sc_hd__nand2_1
X_22406_ _22404_/Y _22405_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _22406_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23386_ hold182/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23386_/X sky130_fd_sc_hd__or2b_1
X_26174_ _26175_/CLK _26174_/D vssd1 vssd1 vccd1 vccd1 _26174_/Q sky130_fd_sc_hd__dfxtp_1
X_20598_ _20601_/A _20601_/C vssd1 vssd1 vccd1 vccd1 _20599_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_162_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22337_ _22338_/A _22338_/C _23055_/A vssd1 vssd1 vccd1 vccd1 _22337_/X sky130_fd_sc_hd__a21o_1
X_25125_ _26335_/CLK _25125_/D vssd1 vssd1 vccd1 vccd1 _25125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25056_ _26142_/CLK _25056_/D vssd1 vssd1 vccd1 vccd1 _25056_/Q sky130_fd_sc_hd__dfxtp_1
X_13070_ _17639_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13070_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22268_ _18594_/A _25819_/Q _22266_/Y _22267_/Y vssd1 vssd1 vccd1 vccd1 _22269_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24007_ _24007_/A vssd1 vssd1 vccd1 vccd1 _26070_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21219_ _21659_/C vssd1 vssd1 vccd1 vccd1 _21662_/B sky130_fd_sc_hd__inv_4
X_22199_ _22197_/X _22198_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _22199_/Y sky130_fd_sc_hd__a21oi_4
X_16760_ _16761_/B _16761_/A vssd1 vssd1 vccd1 vccd1 _16760_/X sky130_fd_sc_hd__or2_1
X_25958_ _26023_/CLK _25958_/D vssd1 vssd1 vccd1 vccd1 _25958_/Q sky130_fd_sc_hd__dfxtp_1
X_13972_ _14061_/A _13972_/B vssd1 vssd1 vccd1 vccd1 _13972_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_38_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15711_ _15712_/B _16937_/A vssd1 vssd1 vccd1 vccd1 _15713_/A sky130_fd_sc_hd__or2_1
X_24909_ _24870_/Y _24959_/B _24892_/X _24908_/Y _23581_/B vssd1 vssd1 vccd1 vccd1
+ _24909_/X sky130_fd_sc_hd__a41o_1
X_12923_ _17435_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12923_/X sky130_fd_sc_hd__or2_1
X_16691_ _16691_/A _16691_/B vssd1 vssd1 vccd1 vccd1 _16692_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25889_ _26084_/CLK _25889_/D vssd1 vssd1 vccd1 vccd1 _25889_/Q sky130_fd_sc_hd__dfxtp_2
X_18430_ _18430_/A _18430_/B _18430_/C vssd1 vssd1 vccd1 vccd1 _22042_/A sky130_fd_sc_hd__nand3_2
X_15642_ _15693_/C vssd1 vssd1 vccd1 vccd1 _15645_/B sky130_fd_sc_hd__inv_2
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12854_ _17296_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12854_/X sky130_fd_sc_hd__or2_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _18361_/A _18361_/B vssd1 vssd1 vccd1 vccd1 _21946_/A sky130_fd_sc_hd__nand2_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15573_ _15560_/A _15549_/A _15548_/B vssd1 vssd1 vccd1 vccd1 _15575_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_150_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12785_ _26092_/Q _12748_/X _12784_/X vssd1 vssd1 vccd1 vccd1 _12785_/X sky130_fd_sc_hd__a21o_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17312_ _17467_/A _17312_/B vssd1 vssd1 vccd1 vccd1 _17312_/Y sky130_fd_sc_hd__nand2_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14524_ _14524_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14524_/Y sky130_fd_sc_hd__nand2_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18292_ _19059_/A _18292_/B vssd1 vssd1 vccd1 vccd1 _18292_/X sky130_fd_sc_hd__xor2_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17243_ _17239_/X _17241_/X _17242_/X vssd1 vssd1 vccd1 vccd1 _17245_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_71_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14455_ _14455_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14455_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_142_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13406_ _13315_/X _13404_/X _23629_/B _13405_/X vssd1 vssd1 vccd1 vccd1 hold996/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17174_ _17393_/A hold977/X _19994_/B vssd1 vssd1 vccd1 vccd1 _17174_/X sky130_fd_sc_hd__and3_1
XFILLER_0_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14386_ _14404_/A hold326/X vssd1 vssd1 vccd1 vccd1 hold327/A sky130_fd_sc_hd__nand2_1
XFILLER_0_109_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16125_ _16125_/A _16125_/B vssd1 vssd1 vccd1 vccd1 _16127_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13337_ _13220_/X _14623_/A _13242_/X _19630_/A vssd1 vssd1 vccd1 vccd1 _13337_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16056_ _16056_/A _16056_/B vssd1 vssd1 vccd1 vccd1 _16056_/X sky130_fd_sc_hd__and2_1
XFILLER_0_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13268_ _26180_/Q _13239_/X _13267_/X vssd1 vssd1 vccd1 vccd1 _13268_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_161_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15007_ _15007_/A _15007_/B vssd1 vssd1 vccd1 vccd1 _15015_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13199_ _18435_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13199_/X sky130_fd_sc_hd__or2_1
Xhold2409 _26188_/Q vssd1 vssd1 vccd1 vccd1 hold2409/X sky130_fd_sc_hd__dlygate4sd3_1
X_19815_ _19812_/Y _19815_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19815_/X sky130_fd_sc_hd__and3b_1
Xhold1708 _25869_/Q vssd1 vssd1 vccd1 vccd1 _22637_/B sky130_fd_sc_hd__buf_1
Xhold1719 _25833_/Q vssd1 vssd1 vccd1 vccd1 _21655_/B sky130_fd_sc_hd__dlygate4sd3_1
X_16958_ _22145_/B _16963_/B vssd1 vssd1 vccd1 vccd1 _16960_/B sky130_fd_sc_hd__nand2_1
X_19746_ _20438_/A _19744_/Y _20443_/C vssd1 vssd1 vccd1 vccd1 _19835_/B sky130_fd_sc_hd__o21a_2
X_15909_ _15909_/A _15909_/B vssd1 vssd1 vccd1 vccd1 _15911_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19677_ _19678_/B _19678_/A vssd1 vssd1 vccd1 vccd1 _19677_/X sky130_fd_sc_hd__or2_1
X_16889_ _16890_/B _16890_/A vssd1 vssd1 vccd1 vccd1 _16889_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_200_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _26235_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_177_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18628_ _18951_/A _18632_/B vssd1 vssd1 vccd1 vccd1 _18630_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18559_ _18559_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18559_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21570_ _21636_/A _21570_/B _21569_/X vssd1 vssd1 vccd1 vccd1 _21571_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_118_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 _23481_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20521_ _23021_/B vssd1 vssd1 vccd1 vccd1 _22441_/B sky130_fd_sc_hd__inv_2
XANTENNA_23 _18007_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 _25581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_45 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_56 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23240_ _23240_/A _24949_/S _24958_/B vssd1 vssd1 vccd1 vccd1 _23243_/A sky130_fd_sc_hd__and3_1
XANTENNA_67 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_78 _25837_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20452_ _20452_/A _20452_/B _21169_/C vssd1 vssd1 vccd1 vccd1 _20456_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23171_ _23171_/A _23187_/B vssd1 vssd1 vccd1 vccd1 _23171_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20383_ _20382_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20383_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22122_ _22122_/A _22122_/B vssd1 vssd1 vccd1 vccd1 _22122_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_141_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22053_ _22053_/A _22053_/B vssd1 vssd1 vccd1 vccd1 _23042_/A sky130_fd_sc_hd__xor2_4
X_21004_ _21480_/C _21529_/C vssd1 vssd1 vccd1 vccd1 _21007_/A sky130_fd_sc_hd__nand2_1
X_25812_ _25812_/CLK _25812_/D vssd1 vssd1 vccd1 vccd1 _25812_/Q sky130_fd_sc_hd__dfxtp_2
X_25743_ _25743_/CLK _25743_/D vssd1 vssd1 vccd1 vccd1 _25743_/Q sky130_fd_sc_hd__dfxtp_1
X_22955_ _22953_/X _22954_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _22955_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21906_ _21906_/A _21906_/B vssd1 vssd1 vccd1 vccd1 _21906_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_69_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25674_ _26305_/CLK _25674_/D vssd1 vssd1 vccd1 vccd1 _25674_/Q sky130_fd_sc_hd__dfxtp_1
X_22886_ _22886_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _22886_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24625_ _24625_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24626_/A sky130_fd_sc_hd__and2_1
X_21837_ _21837_/A _21837_/B vssd1 vssd1 vccd1 vccd1 _21837_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_182_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12570_ _12570_/A _23598_/A vssd1 vssd1 vccd1 vccd1 _12571_/C sky130_fd_sc_hd__nand2_1
X_21768_ _21769_/B _21769_/A vssd1 vssd1 vccd1 vccd1 _21770_/A sky130_fd_sc_hd__or2_1
X_24556_ hold2688/X hold2567/X _24587_/S vssd1 vssd1 vccd1 vccd1 _24557_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_26_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20719_ _20719_/A _20719_/B vssd1 vssd1 vccd1 vccd1 _20721_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_19_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23507_ _23501_/X _23506_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _23507_/X sky130_fd_sc_hd__mux2_1
X_21699_ _21698_/Y _21203_/X _20986_/A _20957_/A vssd1 vssd1 vccd1 vccd1 _21699_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24487_ _24487_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24488_/A sky130_fd_sc_hd__and2_1
XFILLER_0_80_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14240_ _14264_/A _14240_/B vssd1 vssd1 vccd1 vccd1 _14240_/Y sky130_fd_sc_hd__nand2_1
X_26226_ _26226_/CLK _26226_/D vssd1 vssd1 vccd1 vccd1 _26226_/Q sky130_fd_sc_hd__dfxtp_2
X_23438_ _24858_/S vssd1 vssd1 vccd1 vccd1 _24957_/S sky130_fd_sc_hd__buf_12
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14171_ _25822_/Q vssd1 vssd1 vccd1 vccd1 _18653_/B sky130_fd_sc_hd__inv_2
X_23369_ _23369_/A vssd1 vssd1 vccd1 vccd1 _23372_/B sky130_fd_sc_hd__inv_2
XFILLER_0_1_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26157_ _26248_/CLK _26157_/D vssd1 vssd1 vccd1 vccd1 _26157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13122_ _26156_/Q _13065_/X _13121_/X vssd1 vssd1 vccd1 vccd1 _13122_/X sky130_fd_sc_hd__a21o_1
X_25108_ _26317_/CLK _25108_/D vssd1 vssd1 vccd1 vccd1 _25108_/Q sky130_fd_sc_hd__dfxtp_1
X_26088_ _26089_/CLK _26088_/D vssd1 vssd1 vccd1 vccd1 _26088_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17930_ _17930_/A _25777_/Q vssd1 vssd1 vccd1 vccd1 _20141_/A sky130_fd_sc_hd__nand2_1
X_13053_ _17617_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13053_/X sky130_fd_sc_hd__or2_1
XFILLER_0_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25039_ _26122_/CLK _25039_/D vssd1 vssd1 vccd1 vccd1 _25039_/Q sky130_fd_sc_hd__dfxtp_1
X_17861_ _17861_/A _20428_/A vssd1 vssd1 vccd1 vccd1 _19045_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16812_ _16812_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16812_/Y sky130_fd_sc_hd__nand2_1
X_19600_ _19599_/Y _19272_/X _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19601_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_108_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17792_ _18611_/A _17800_/B vssd1 vssd1 vccd1 vccd1 _17796_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19531_ _19528_/Y _19531_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19531_/X sky130_fd_sc_hd__and3b_1
X_16743_ _16858_/A _16743_/B vssd1 vssd1 vccd1 vccd1 _16743_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13955_ hold729/X _13954_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold730/A sky130_fd_sc_hd__a21oi_1
X_12906_ _12840_/X _12904_/X _12827_/X _12905_/X vssd1 vssd1 vccd1 vccd1 _12906_/X
+ sky130_fd_sc_hd__o211a_1
X_19462_ _19463_/B _19463_/A vssd1 vssd1 vccd1 vccd1 _19462_/X sky130_fd_sc_hd__or2_1
X_16674_ _16672_/Y hold690/X _16594_/X vssd1 vssd1 vccd1 vccd1 hold691/A sky130_fd_sc_hd__a21oi_1
X_13886_ hold708/X _13885_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold709/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18413_ _18413_/A _18413_/B vssd1 vssd1 vccd1 vccd1 _18413_/X sky130_fd_sc_hd__xor2_1
X_15625_ _15625_/A _16904_/A vssd1 vssd1 vccd1 vccd1 _15626_/B sky130_fd_sc_hd__nor2_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12837_ _26102_/Q _12748_/X _12836_/X vssd1 vssd1 vccd1 vccd1 _12837_/X sky130_fd_sc_hd__a21o_1
X_19393_ _19393_/A _19393_/B vssd1 vssd1 vccd1 vccd1 _19393_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_68_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18344_ _18446_/A _25743_/Q _18952_/C vssd1 vssd1 vccd1 vccd1 _18345_/C sky130_fd_sc_hd__nand3_1
X_15556_ _15469_/Y _15552_/B _15555_/Y vssd1 vssd1 vccd1 vccd1 _15557_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12768_ _26217_/Q _25586_/Q vssd1 vssd1 vccd1 vccd1 _14301_/A sky130_fd_sc_hd__xor2_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14507_ _14525_/A hold20/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__nand2_1
X_18275_ _18272_/Y _18274_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25658_/D sky130_fd_sc_hd__a21oi_1
X_15487_ _25562_/Q vssd1 vssd1 vccd1 vccd1 _22896_/B sky130_fd_sc_hd__inv_2
XFILLER_0_127_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12699_ _12699_/A vssd1 vssd1 vccd1 vccd1 _12704_/A sky130_fd_sc_hd__inv_2
XFILLER_0_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17226_ _17470_/A _17226_/B vssd1 vssd1 vccd1 vccd1 _17226_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_181_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14438_ _14465_/A hold122/X vssd1 vssd1 vccd1 vccd1 hold123/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17157_ _20479_/B _25889_/Q _25825_/Q vssd1 vssd1 vccd1 vccd1 _17158_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_123_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14369_ _14367_/Y hold84/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__a21oi_1
Xhold805 hold805/A vssd1 vssd1 vccd1 vccd1 hold805/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold816 hold816/A vssd1 vssd1 vccd1 vccd1 hold816/X sky130_fd_sc_hd__dlygate4sd3_1
X_16108_ _16097_/B _16103_/B _16106_/Y _16107_/Y _16096_/A vssd1 vssd1 vccd1 vccd1
+ _16109_/A sky130_fd_sc_hd__o221ai_4
XFILLER_0_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold827 hold827/A vssd1 vssd1 vccd1 vccd1 hold827/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 hold838/A vssd1 vssd1 vccd1 vccd1 hold838/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold849 hold849/A vssd1 vssd1 vccd1 vccd1 hold849/X sky130_fd_sc_hd__dlygate4sd3_1
X_17088_ _25628_/Q vssd1 vssd1 vccd1 vccd1 _20273_/B sky130_fd_sc_hd__inv_2
XFILLER_0_126_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16039_ _16039_/A _16039_/B vssd1 vssd1 vccd1 vccd1 _16052_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2206 _25419_/Q vssd1 vssd1 vccd1 vccd1 _14955_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2217 _23776_/X vssd1 vssd1 vccd1 vccd1 _23777_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2228 _12651_/Y vssd1 vssd1 vccd1 vccd1 _12661_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2239 _26086_/Q vssd1 vssd1 vccd1 vccd1 hold2239/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1505 _25096_/Q vssd1 vssd1 vccd1 vccd1 _18638_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1516 _13376_/X vssd1 vssd1 vccd1 vccd1 _25114_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1527 _25728_/Q vssd1 vssd1 vccd1 vccd1 _19381_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1538 _20161_/Y vssd1 vssd1 vccd1 vccd1 _25777_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1549 _25118_/Q vssd1 vssd1 vccd1 vccd1 _19005_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19729_ _19729_/A _20401_/B vssd1 vssd1 vccd1 vccd1 _19729_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22740_ _22937_/A _22740_/B vssd1 vssd1 vccd1 vccd1 _22740_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22671_ _22671_/A _22671_/B vssd1 vssd1 vccd1 vccd1 _23152_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_149_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24410_ _24410_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24411_/A sky130_fd_sc_hd__and2_1
X_21622_ _21622_/A _22902_/B vssd1 vssd1 vccd1 vccd1 _21622_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xascon_wrapper_18 vssd1 vssd1 vccd1 vccd1 io_oeb[4] ascon_wrapper_18/LO sky130_fd_sc_hd__conb_1
XFILLER_0_34_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25390_ _26004_/CLK _25390_/D vssd1 vssd1 vccd1 vccd1 _25390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21553_ _21552_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21553_/X
+ sky130_fd_sc_hd__a211o_1
X_24341_ _26178_/Q hold2332/X _24356_/S vssd1 vssd1 vccd1 vccd1 _24341_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_145_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20504_ _20660_/A _20504_/B vssd1 vssd1 vccd1 vccd1 _20504_/Y sky130_fd_sc_hd__nand2_1
X_24272_ _24272_/A vssd1 vssd1 vccd1 vccd1 _26156_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21484_ _21484_/A _21484_/B vssd1 vssd1 vccd1 vccd1 _21485_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_172_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23223_ _24871_/B _23253_/C vssd1 vssd1 vccd1 vccd1 _23240_/A sky130_fd_sc_hd__nor2_1
X_26011_ _26012_/CLK _26011_/D vssd1 vssd1 vccd1 vccd1 _26011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20435_ _20434_/B _20435_/B _20435_/C vssd1 vssd1 vccd1 vccd1 _20436_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_160_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23154_ _23154_/A _23154_/B vssd1 vssd1 vccd1 vccd1 _23155_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_30_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20366_ _20366_/A _22353_/B _20366_/C vssd1 vssd1 vccd1 vccd1 _20370_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_105_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22105_ _25849_/Q _25785_/Q vssd1 vssd1 vccd1 vccd1 _22106_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_105_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23085_ _23197_/A _23085_/B vssd1 vssd1 vccd1 vccd1 _23085_/Y sky130_fd_sc_hd__nand2_1
X_20297_ _20297_/A _21062_/B vssd1 vssd1 vccd1 vccd1 _20299_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22036_ _22036_/A _22145_/B vssd1 vssd1 vccd1 vccd1 _22036_/Y sky130_fd_sc_hd__nand2_1
Xhold2740 _24591_/X vssd1 vssd1 vccd1 vccd1 _24592_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2751 _25916_/Q vssd1 vssd1 vccd1 vccd1 _23276_/C sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23987_ _23987_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23988_/A sky130_fd_sc_hd__and2_1
X_25726_ _25729_/CLK _25726_/D vssd1 vssd1 vccd1 vccd1 _25726_/Q sky130_fd_sc_hd__dfxtp_1
X_13740_ _13823_/A _13740_/B vssd1 vssd1 vccd1 vccd1 _13740_/Y sky130_fd_sc_hd__nand2_1
X_22938_ _22936_/X _22937_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _22938_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25657_ _26289_/CLK _25657_/D vssd1 vssd1 vccd1 vccd1 _25657_/Q sky130_fd_sc_hd__dfxtp_4
X_13671_ _26245_/Q _13612_/X _13605_/X _13670_/Y vssd1 vssd1 vccd1 vccd1 _13672_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22869_ _16842_/B _22421_/X _22863_/X _22864_/Y _22868_/X vssd1 vssd1 vccd1 vccd1
+ _22870_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_35_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15410_ _15375_/X _15406_/A _15409_/X vssd1 vssd1 vccd1 vccd1 _15411_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12622_ _12645_/B _12624_/A vssd1 vssd1 vccd1 vccd1 _12629_/A sky130_fd_sc_hd__nor2_1
X_24608_ _24608_/A vssd1 vssd1 vccd1 vccd1 _26265_/D sky130_fd_sc_hd__clkbuf_1
X_16390_ _16390_/A _16390_/B vssd1 vssd1 vccd1 vccd1 _16391_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_149_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25588_ _25594_/CLK _25588_/D vssd1 vssd1 vccd1 vccd1 _25588_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_183_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15341_ _15341_/A _16796_/A vssd1 vssd1 vccd1 vccd1 _15342_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_164_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24539_ _24539_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24540_/A sky130_fd_sc_hd__and2_1
X_12553_ _17748_/B vssd1 vssd1 vccd1 vccd1 _17688_/B sky130_fd_sc_hd__inv_2
XFILLER_0_109_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18060_ _18060_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _18060_/Y sky130_fd_sc_hd__nand2_1
X_15272_ _15272_/A _15272_/B vssd1 vssd1 vccd1 vccd1 _15275_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12484_ _15773_/S vssd1 vssd1 vccd1 vccd1 _14277_/B sky130_fd_sc_hd__inv_6
XFILLER_0_108_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17011_ _21791_/A vssd1 vssd1 vccd1 vccd1 _17229_/B sky130_fd_sc_hd__buf_8
X_26209_ _26336_/CLK _26209_/D vssd1 vssd1 vccd1 vccd1 _26209_/Q sky130_fd_sc_hd__dfxtp_1
X_14223_ hold399/X _14222_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold400/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14154_ _14180_/A _14154_/B vssd1 vssd1 vccd1 vccd1 _14154_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_132_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13105_ _13049_/X _14503_/A _13067_/X _25650_/Q vssd1 vssd1 vccd1 vccd1 _13105_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14085_ _26311_/Q _13988_/X _13981_/X _14084_/Y vssd1 vssd1 vccd1 vccd1 _14086_/B
+ sky130_fd_sc_hd__a22o_1
X_18962_ _18960_/X _18879_/X _18961_/X vssd1 vssd1 vccd1 vccd1 _18963_/A sky130_fd_sc_hd__a21o_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17913_ _19032_/A _17913_/B vssd1 vssd1 vccd1 vccd1 _17913_/X sky130_fd_sc_hd__xor2_1
X_13036_ _26140_/Q _12907_/X _13035_/X vssd1 vssd1 vccd1 vccd1 _13036_/X sky130_fd_sc_hd__a21o_1
X_18893_ _18954_/A _25770_/Q vssd1 vssd1 vccd1 vccd1 _18895_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17844_ _17844_/A _20738_/B _17844_/C vssd1 vssd1 vccd1 vccd1 _20707_/B sky130_fd_sc_hd__nand3_2
X_17775_ _17775_/A _18118_/B _17775_/C vssd1 vssd1 vccd1 vccd1 _18118_/A sky130_fd_sc_hd__nand3_4
X_14987_ _14985_/X hold2231/X _14928_/X vssd1 vssd1 vccd1 vccd1 _14987_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16726_ _16726_/A _16726_/B vssd1 vssd1 vccd1 vccd1 _16726_/Y sky130_fd_sc_hd__nand2_1
X_19514_ _26241_/Q _19483_/X hold596/X vssd1 vssd1 vccd1 vccd1 _19514_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13938_ _25785_/Q vssd1 vssd1 vccd1 vccd1 _17859_/B sky130_fd_sc_hd__inv_2
XFILLER_0_53_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19445_ _21047_/A _21773_/B _25611_/Q vssd1 vssd1 vccd1 vccd1 _21051_/C sky130_fd_sc_hd__nand3_1
X_16657_ _16659_/B vssd1 vssd1 vccd1 vccd1 _16680_/B sky130_fd_sc_hd__inv_2
XFILLER_0_187_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13869_ _20041_/B vssd1 vssd1 vccd1 vccd1 _17665_/B sky130_fd_sc_hd__inv_2
XFILLER_0_88_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15608_ _15609_/B _15609_/A vssd1 vssd1 vccd1 vccd1 _15608_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19376_ _19393_/B _19463_/B vssd1 vssd1 vccd1 vccd1 _19378_/A sky130_fd_sc_hd__xnor2_1
X_16588_ _16588_/A _16588_/B vssd1 vssd1 vccd1 vccd1 _16596_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_173_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18327_ _18952_/A _18327_/B _18952_/C vssd1 vssd1 vccd1 vccd1 _18328_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_174_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15539_ _15539_/A _15774_/B vssd1 vssd1 vccd1 vccd1 _15540_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_127_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18258_ _25867_/Q _21772_/A vssd1 vssd1 vccd1 vccd1 _18266_/A sky130_fd_sc_hd__or2_2
XFILLER_0_72_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17209_ _25637_/Q vssd1 vssd1 vccd1 vccd1 _20635_/B sky130_fd_sc_hd__inv_2
XFILLER_0_4_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18189_ _18189_/A _18189_/B vssd1 vssd1 vccd1 vccd1 _18191_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold602 hold602/A vssd1 vssd1 vccd1 vccd1 hold602/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold613 hold613/A vssd1 vssd1 vccd1 vccd1 hold613/X sky130_fd_sc_hd__dlygate4sd3_1
X_20220_ _21449_/A _21089_/B vssd1 vssd1 vccd1 vccd1 _20224_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold624 hold624/A vssd1 vssd1 vccd1 vccd1 hold624/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold635 hold635/A vssd1 vssd1 vccd1 vccd1 hold635/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 hold646/A vssd1 vssd1 vccd1 vccd1 hold646/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold657 hold657/A vssd1 vssd1 vccd1 vccd1 hold657/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20151_ _20151_/A _20151_/B _20952_/B vssd1 vssd1 vccd1 vccd1 _20152_/B sky130_fd_sc_hd__nand3_1
Xhold668 hold668/A vssd1 vssd1 vccd1 vccd1 hold668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 hold679/A vssd1 vssd1 vccd1 vccd1 hold679/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2003 _26039_/Q vssd1 vssd1 vccd1 vccd1 hold2003/X sky130_fd_sc_hd__dlygate4sd3_1
X_20082_ _21042_/A _20082_/B _20081_/X vssd1 vssd1 vccd1 vccd1 _20083_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_110_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2014 _12639_/Y vssd1 vssd1 vccd1 vccd1 _12640_/C sky130_fd_sc_hd__dlygate4sd3_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2025 _25985_/Q vssd1 vssd1 vccd1 vccd1 _14733_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2036 _26008_/Q vssd1 vssd1 vccd1 vccd1 hold2036/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23910_ _23910_/A vssd1 vssd1 vccd1 vccd1 _26040_/D sky130_fd_sc_hd__clkbuf_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2047 _24166_/X vssd1 vssd1 vccd1 vccd1 _24167_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1302 _25058_/Q vssd1 vssd1 vccd1 vccd1 _17602_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1313 _13134_/X vssd1 vssd1 vccd1 vccd1 _25075_/D sky130_fd_sc_hd__dlygate4sd3_1
X_24890_ _24887_/Y _24889_/Y _24867_/S _24959_/C vssd1 vssd1 vccd1 vccd1 _24890_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_176_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2058 _26166_/Q vssd1 vssd1 vccd1 vccd1 hold2058/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2069 _23650_/X vssd1 vssd1 vccd1 vccd1 _23651_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1324 _12817_/X vssd1 vssd1 vccd1 vccd1 _25015_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1335 _25789_/Q vssd1 vssd1 vccd1 vccd1 _20622_/B sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1346 _20992_/Y vssd1 vssd1 vccd1 vccd1 _25800_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23841_ hold2119/X hold2051/X _23907_/S vssd1 vssd1 vccd1 vccd1 _23842_/A sky130_fd_sc_hd__mux2_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1357 _25090_/Q vssd1 vssd1 vccd1 vccd1 _18515_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1368 _13001_/X vssd1 vssd1 vccd1 vccd1 _25050_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1379 _25787_/Q vssd1 vssd1 vccd1 vccd1 _20544_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23772_ _23772_/A vssd1 vssd1 vccd1 vccd1 _25995_/D sky130_fd_sc_hd__clkbuf_1
X_20984_ _26303_/Q _20731_/X hold710/X vssd1 vssd1 vccd1 vccd1 _20988_/B sky130_fd_sc_hd__a21oi_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25511_ _25511_/CLK hold874/X vssd1 vssd1 vccd1 vccd1 hold873/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22723_ _22723_/A _22723_/B vssd1 vssd1 vccd1 vccd1 _22724_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25442_ _26052_/CLK hold886/X vssd1 vssd1 vccd1 vccd1 hold885/A sky130_fd_sc_hd__dfxtp_1
X_22654_ _15257_/B _22387_/B _14273_/X vssd1 vssd1 vccd1 vccd1 _22654_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_164_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21605_ _21605_/A _22902_/B vssd1 vssd1 vccd1 vccd1 _21605_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22585_ _22576_/Y _22584_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22585_/X sky130_fd_sc_hd__a21o_1
X_25373_ _26198_/CLK hold469/X vssd1 vssd1 vccd1 vccd1 hold467/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24324_ _24324_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24325_/A sky130_fd_sc_hd__and2_1
XFILLER_0_91_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21536_ _26329_/Q hold827/X vssd1 vssd1 vccd1 vccd1 _21536_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_118_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24255_ hold2237/X hold1995/X _24279_/S vssd1 vssd1 vccd1 vccd1 _24256_/A sky130_fd_sc_hd__mux2_1
X_21467_ _21467_/A _21467_/B _21467_/C vssd1 vssd1 vccd1 vccd1 _21468_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_105_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23206_ _23206_/A vssd1 vssd1 vccd1 vccd1 _25904_/D sky130_fd_sc_hd__inv_2
XFILLER_0_31_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20418_ _20418_/A _20418_/B vssd1 vssd1 vccd1 vccd1 _20419_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_160_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24186_ _24186_/A vssd1 vssd1 vccd1 vccd1 _26128_/D sky130_fd_sc_hd__clkbuf_1
X_21398_ _21401_/A _21450_/A vssd1 vssd1 vccd1 vccd1 _21400_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23137_ _23137_/A _23137_/B vssd1 vssd1 vccd1 vccd1 _23138_/B sky130_fd_sc_hd__nand2_1
X_20349_ _20349_/A _22051_/A vssd1 vssd1 vccd1 vccd1 _20350_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_105_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23068_ _23059_/Y _23067_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _23068_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_175_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14910_ _14910_/A _14910_/B _14910_/C vssd1 vssd1 vccd1 vccd1 _14910_/Y sky130_fd_sc_hd__nand3_1
X_22019_ _25874_/Q _22020_/A vssd1 vssd1 vccd1 vccd1 _22021_/A sky130_fd_sc_hd__or2_1
XFILLER_0_175_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15890_ _15891_/B _15891_/A vssd1 vssd1 vccd1 vccd1 _15909_/B sky130_fd_sc_hd__or2_1
XFILLER_0_179_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2570 _15610_/Y vssd1 vssd1 vccd1 vccd1 _25463_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14841_ _14839_/Y _14840_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 hold956/A sky130_fd_sc_hd__a21oi_1
Xhold2581 _24707_/X vssd1 vssd1 vccd1 vccd1 _24708_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2592 _26216_/Q vssd1 vssd1 vccd1 vccd1 hold2592/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1880 _25845_/Q vssd1 vssd1 vccd1 vccd1 _21999_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17560_ _17605_/A _17560_/B vssd1 vssd1 vccd1 vccd1 _17560_/Y sky130_fd_sc_hd__nand2_1
X_14772_ _22001_/B _15778_/B vssd1 vssd1 vccd1 vccd1 _14773_/A sky130_fd_sc_hd__nand2_1
Xhold1891 _26175_/Q vssd1 vssd1 vccd1 vccd1 hold1891/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16511_ _16511_/A _16511_/B vssd1 vssd1 vccd1 vccd1 _16512_/A sky130_fd_sc_hd__nor2_1
X_13723_ _13718_/Y _13722_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold926/A sky130_fd_sc_hd__a21oi_1
X_25709_ _25709_/CLK _25709_/D vssd1 vssd1 vccd1 vccd1 _25709_/Q sky130_fd_sc_hd__dfxtp_4
X_17491_ _17491_/A _17541_/A vssd1 vssd1 vccd1 vccd1 _17492_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19230_ _19230_/A _20547_/B vssd1 vssd1 vccd1 vccd1 _19230_/Y sky130_fd_sc_hd__nor2_1
X_16442_ _16442_/A _16442_/B vssd1 vssd1 vccd1 vccd1 _16442_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_168_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ _13703_/A _13654_/B vssd1 vssd1 vccd1 vccd1 _13654_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12605_ _12610_/A _12643_/B vssd1 vssd1 vccd1 vccd1 _12605_/Y sky130_fd_sc_hd__nand2_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19161_ _19159_/A _19158_/Y _20175_/A vssd1 vssd1 vccd1 vccd1 _19983_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_109_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16373_ _16374_/A _16374_/B _16378_/B vssd1 vssd1 vccd1 vccd1 _16373_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_155_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _13642_/A hold590/X vssd1 vssd1 vccd1 vccd1 hold591/A sky130_fd_sc_hd__nand2_1
XFILLER_0_171_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18112_ _21099_/A vssd1 vssd1 vccd1 vccd1 _18112_/X sky130_fd_sc_hd__buf_8
X_15324_ _15324_/A _15326_/A vssd1 vssd1 vccd1 vccd1 _15324_/Y sky130_fd_sc_hd__nand2_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12536_ _15795_/A vssd1 vssd1 vccd1 vccd1 _15621_/A sky130_fd_sc_hd__buf_8
XFILLER_0_147_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19092_ _19093_/A vssd1 vssd1 vccd1 vccd1 _19092_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18043_ _18528_/A vssd1 vssd1 vccd1 vccd1 _18445_/A sky130_fd_sc_hd__buf_12
XFILLER_0_83_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15255_ _26013_/Q _25949_/Q _15773_/S vssd1 vssd1 vccd1 vccd1 _15256_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_151_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14206_ _14236_/A hold473/X vssd1 vssd1 vccd1 vccd1 hold474/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15186_ _15184_/A _15161_/B _15178_/A vssd1 vssd1 vccd1 vccd1 _15186_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14137_ _14132_/Y _14136_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold732/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19994_ _19994_/A _19994_/B _19994_/C vssd1 vssd1 vccd1 vccd1 _19994_/X sky130_fd_sc_hd__and3_1
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14068_ _14180_/A _14068_/B vssd1 vssd1 vccd1 vccd1 _14068_/Y sky130_fd_sc_hd__nand2_1
X_18945_ _18943_/Y _18944_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _18945_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_183_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13019_ _26265_/Q _25634_/Q vssd1 vssd1 vccd1 vccd1 _14452_/A sky130_fd_sc_hd__xor2_2
X_18876_ _18876_/A _20790_/A vssd1 vssd1 vccd1 vccd1 _19052_/B sky130_fd_sc_hd__xor2_4
X_17827_ _25839_/Q vssd1 vssd1 vccd1 vccd1 _20069_/A sky130_fd_sc_hd__inv_2
X_17758_ _17924_/B _17924_/A vssd1 vssd1 vccd1 vccd1 _17925_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16709_ _16980_/A _16715_/B vssd1 vssd1 vccd1 vccd1 _16712_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_76_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17689_ _17693_/C vssd1 vssd1 vccd1 vccd1 _17690_/C sky130_fd_sc_hd__inv_2
XFILLER_0_147_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19428_ _19427_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19429_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19359_ _19359_/A _20883_/B vssd1 vssd1 vccd1 vccd1 _19359_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_45_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22370_ _25823_/Q _22370_/B vssd1 vssd1 vccd1 vccd1 _22370_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21321_ _21675_/C _21370_/A vssd1 vssd1 vccd1 vccd1 _21322_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold410 hold410/A vssd1 vssd1 vccd1 vccd1 hold410/X sky130_fd_sc_hd__dlygate4sd3_1
X_24040_ _24040_/A vssd1 vssd1 vccd1 vccd1 _26081_/D sky130_fd_sc_hd__clkbuf_1
X_21252_ _21252_/A _21252_/B _21252_/C vssd1 vssd1 vccd1 vccd1 _21253_/B sky130_fd_sc_hd__nand3_1
Xhold421 hold421/A vssd1 vssd1 vccd1 vccd1 hold421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 hold432/A vssd1 vssd1 vccd1 vccd1 hold432/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 hold443/A vssd1 vssd1 vccd1 vccd1 hold443/X sky130_fd_sc_hd__dlygate4sd3_1
X_20203_ _25882_/Q vssd1 vssd1 vccd1 vccd1 _20204_/B sky130_fd_sc_hd__inv_2
XFILLER_0_130_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold454 hold454/A vssd1 vssd1 vccd1 vccd1 hold454/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21183_ _21183_/A _21947_/B vssd1 vssd1 vccd1 vccd1 _21184_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_141_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold465 hold465/A vssd1 vssd1 vccd1 vccd1 hold465/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 hold476/A vssd1 vssd1 vccd1 vccd1 hold476/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold487 hold487/A vssd1 vssd1 vccd1 vccd1 hold487/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 hold498/A vssd1 vssd1 vccd1 vccd1 hold498/X sky130_fd_sc_hd__dlygate4sd3_1
X_20134_ _20134_/A _25880_/Q vssd1 vssd1 vccd1 vccd1 _20139_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25991_ _25991_/CLK _25991_/D vssd1 vssd1 vccd1 vccd1 _25991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24942_ hold906/A hold968/A _24942_/S vssd1 vssd1 vccd1 vccd1 _24943_/B sky130_fd_sc_hd__mux2_1
X_20065_ _21386_/A vssd1 vssd1 vccd1 vccd1 _21385_/A sky130_fd_sc_hd__inv_2
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 _13054_/X vssd1 vssd1 vccd1 vccd1 _25060_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 _25128_/Q vssd1 vssd1 vccd1 vccd1 _19075_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1132 _21073_/Y vssd1 vssd1 vccd1 vccd1 _25803_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24873_ _24873_/A _24946_/A vssd1 vssd1 vccd1 vccd1 _24873_/Y sky130_fd_sc_hd__nand2_1
Xhold1143 _25011_/Q vssd1 vssd1 vccd1 vccd1 _17148_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1154 _19682_/Y vssd1 vssd1 vccd1 vccd1 _25749_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1165 _25091_/Q vssd1 vssd1 vccd1 vccd1 _18535_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 _16942_/Y vssd1 vssd1 vccd1 vccd1 _25574_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23824_ _23824_/A vssd1 vssd1 vccd1 vccd1 _26012_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1187 _25032_/Q vssd1 vssd1 vccd1 vccd1 _17404_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1198 _13418_/X vssd1 vssd1 vccd1 vccd1 _25121_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23755_ _23755_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23756_/A sky130_fd_sc_hd__and2_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20967_ _20967_/A _25864_/Q vssd1 vssd1 vccd1 vccd1 _20973_/A sky130_fd_sc_hd__nand2_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22706_ _23188_/A _22706_/B vssd1 vssd1 vccd1 vccd1 _22706_/X sky130_fd_sc_hd__or2_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23686_ _23686_/A vssd1 vssd1 vccd1 vccd1 _25967_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20898_ _20898_/A _20898_/B vssd1 vssd1 vccd1 vccd1 _20899_/A sky130_fd_sc_hd__nand2_1
X_25425_ _25425_/CLK _25425_/D vssd1 vssd1 vccd1 vccd1 _25425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22637_ _22937_/A _22637_/B vssd1 vssd1 vccd1 vccd1 _22637_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_119_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25356_ _26308_/CLK hold187/X vssd1 vssd1 vccd1 vccd1 hold185/A sky130_fd_sc_hd__dfxtp_1
X_13370_ _13315_/X _13368_/X _13300_/X _13369_/X vssd1 vssd1 vccd1 vccd1 _13370_/X
+ sky130_fd_sc_hd__o211a_1
X_22568_ _22569_/B _22569_/A vssd1 vssd1 vccd1 vccd1 _22570_/A sky130_fd_sc_hd__or2_1
XFILLER_0_152_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24307_ _24307_/A vssd1 vssd1 vccd1 vccd1 _26167_/D sky130_fd_sc_hd__clkbuf_1
X_21519_ _26328_/Q _21228_/X hold422/X vssd1 vssd1 vccd1 vccd1 _21522_/B sky130_fd_sc_hd__a21oi_1
X_25287_ _26240_/CLK hold220/X vssd1 vssd1 vccd1 vccd1 hold218/A sky130_fd_sc_hd__dfxtp_1
X_22499_ _23168_/A _22499_/B vssd1 vssd1 vccd1 vccd1 _22500_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15040_ _15038_/X hold2375/X _14928_/X vssd1 vssd1 vccd1 vccd1 _15040_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24238_ _24238_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24239_/A sky130_fd_sc_hd__and2_1
XFILLER_0_43_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24169_ hold2302/X _26123_/Q _24203_/S vssd1 vssd1 vccd1 vccd1 _24169_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16991_ _19616_/A _16991_/B vssd1 vssd1 vccd1 vccd1 _17491_/A sky130_fd_sc_hd__xor2_4
X_15942_ _15942_/A _15942_/B vssd1 vssd1 vccd1 vccd1 _16273_/B sky130_fd_sc_hd__and2_1
X_18730_ _18793_/A _25762_/Q _18891_/C vssd1 vssd1 vccd1 vccd1 _18731_/C sky130_fd_sc_hd__nand3_1
X_18661_ _19199_/A vssd1 vssd1 vccd1 vccd1 _18986_/A sky130_fd_sc_hd__clkbuf_8
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ _16660_/B vssd1 vssd1 vccd1 vccd1 _16697_/B sky130_fd_sc_hd__buf_8
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14824_ _15839_/A _14824_/B vssd1 vssd1 vccd1 vccd1 _22175_/A sky130_fd_sc_hd__nand2_1
X_17612_ _19199_/A vssd1 vssd1 vccd1 vccd1 _18252_/A sky130_fd_sc_hd__buf_8
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18592_ _18592_/A _18592_/B _18592_/C vssd1 vssd1 vccd1 vccd1 _22269_/A sky130_fd_sc_hd__nand3_2
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17543_ _17624_/A _17543_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17543_/X sky130_fd_sc_hd__and3_1
XFILLER_0_59_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ _14755_/A vssd1 vssd1 vccd1 vccd1 _14945_/A sky130_fd_sc_hd__inv_2
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13706_ _13944_/A vssd1 vssd1 vccd1 vccd1 _13823_/A sky130_fd_sc_hd__buf_6
XFILLER_0_169_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17474_ _19199_/A vssd1 vssd1 vccd1 vccd1 _17605_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14686_ _14684_/Y hold318/X _14646_/X vssd1 vssd1 vccd1 vccd1 hold319/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16425_ hold933/X _16426_/A vssd1 vssd1 vccd1 vccd1 _16427_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_6_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19213_ _19205_/X _19212_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19213_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_184_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13637_ _25737_/Q vssd1 vssd1 vccd1 vccd1 _18223_/B sky130_fd_sc_hd__inv_2
XFILLER_0_172_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19144_ _19961_/B _19145_/A vssd1 vssd1 vccd1 vccd1 _19144_/X sky130_fd_sc_hd__or2_1
X_16356_ _16356_/A _16401_/C vssd1 vssd1 vccd1 vccd1 _16358_/A sky130_fd_sc_hd__nand2_1
X_13568_ _25726_/Q vssd1 vssd1 vccd1 vccd1 _18086_/B sky130_fd_sc_hd__inv_2
XFILLER_0_171_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15307_ _15307_/A _15307_/B vssd1 vssd1 vccd1 vccd1 _15327_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_136_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12519_ _12537_/B _12497_/Y _12518_/Y _23278_/B vssd1 vssd1 vccd1 vccd1 _12519_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19075_ _19082_/A _19075_/B _22786_/A vssd1 vssd1 vccd1 vccd1 _19075_/X sky130_fd_sc_hd__and3_1
XFILLER_0_70_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16287_ _16309_/A _16287_/B vssd1 vssd1 vccd1 vccd1 _16297_/A sky130_fd_sc_hd__or2_1
XFILLER_0_41_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13499_ _25715_/Q vssd1 vssd1 vccd1 vccd1 _13500_/A sky130_fd_sc_hd__inv_2
XFILLER_0_180_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18026_ _22219_/B _25597_/Q vssd1 vssd1 vccd1 vccd1 _18028_/A sky130_fd_sc_hd__nand2_1
X_15238_ _15238_/A vssd1 vssd1 vccd1 vccd1 _15247_/B sky130_fd_sc_hd__inv_2
XFILLER_0_164_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169_ _15169_/A vssd1 vssd1 vccd1 vccd1 _15177_/B sky130_fd_sc_hd__inv_2
XFILLER_0_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19977_ _26275_/Q hold806/X vssd1 vssd1 vccd1 vccd1 _19977_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18928_ _25644_/Q _22692_/B vssd1 vssd1 vccd1 vccd1 _18929_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_66_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18859_ _19026_/A _18859_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18859_/X sky130_fd_sc_hd__and3_1
XFILLER_0_98_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21870_ _18104_/A _25797_/Q _21868_/Y _21869_/Y vssd1 vssd1 vccd1 vccd1 _21871_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20821_ _25859_/Q vssd1 vssd1 vccd1 vccd1 _21806_/B sky130_fd_sc_hd__inv_2
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23540_ hold74/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23540_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_148_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20752_ _20752_/A _20752_/B vssd1 vssd1 vccd1 vccd1 _20756_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_175_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20683_ _21368_/C _21645_/B vssd1 vssd1 vccd1 vccd1 _20686_/A sky130_fd_sc_hd__nand2_1
X_23471_ _24956_/S hold479/A _23470_/X vssd1 vssd1 vccd1 vccd1 _23471_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25210_ _26292_/CLK hold640/X vssd1 vssd1 vccd1 vccd1 hold638/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22422_ _23191_/C vssd1 vssd1 vccd1 vccd1 _22424_/B sky130_fd_sc_hd__inv_2
XFILLER_0_169_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26190_ _26190_/CLK _26190_/D vssd1 vssd1 vccd1 vccd1 _26190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25141_ _26234_/CLK hold460/X vssd1 vssd1 vccd1 vccd1 hold458/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22353_ _22353_/A _22353_/B vssd1 vssd1 vccd1 vccd1 _22354_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_72_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21304_ _21659_/C _21707_/C vssd1 vssd1 vccd1 vccd1 _21305_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_131_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22284_ _22284_/A _22284_/B vssd1 vssd1 vccd1 vccd1 _23023_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_60_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25072_ _26284_/CLK _25072_/D vssd1 vssd1 vccd1 vccd1 _25072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24023_ hold2487/X hold2458/X _24047_/S vssd1 vssd1 vccd1 vccd1 _24024_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_41_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21235_ _21235_/A _21235_/B vssd1 vssd1 vccd1 vccd1 _21235_/Y sky130_fd_sc_hd__nand2_1
Xhold240 hold240/A vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 hold251/A vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 hold262/A vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold273 hold273/A vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold284 hold284/A vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
X_21166_ _21577_/C _21630_/B vssd1 vssd1 vccd1 vccd1 _21169_/A sky130_fd_sc_hd__nand2_1
Xhold295 hold295/A vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20117_ _20117_/A _20117_/B _21010_/B vssd1 vssd1 vccd1 vccd1 _20121_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_102_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25974_ _26040_/CLK _25974_/D vssd1 vssd1 vccd1 vccd1 _25974_/Q sky130_fd_sc_hd__dfxtp_1
X_21097_ _21097_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _21097_/Y sky130_fd_sc_hd__nand2_1
X_24925_ hold864/A _25527_/Q _24944_/S vssd1 vssd1 vccd1 vccd1 _24926_/B sky130_fd_sc_hd__mux2_1
X_20048_ _20048_/A _25900_/Q _20048_/C vssd1 vssd1 vccd1 vccd1 _20051_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_77_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24856_ _15480_/A _15495_/B _24860_/S vssd1 vssd1 vccd1 vccd1 _24856_/X sky130_fd_sc_hd__mux2_1
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _12840_/X _12868_/X _12827_/X _12869_/X vssd1 vssd1 vccd1 vccd1 hold984/A
+ sky130_fd_sc_hd__o211a_1
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23807_ _23807_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23808_/A sky130_fd_sc_hd__and2_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24787_ hold2410/X hold1918/X _24817_/S vssd1 vssd1 vccd1 vccd1 _24788_/A sky130_fd_sc_hd__mux2_1
X_21999_ _22058_/A _21999_/B vssd1 vssd1 vccd1 vccd1 _21999_/Y sky130_fd_sc_hd__nand2_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _14585_/A hold95/X vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__nand2_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23738_ _23738_/A vssd1 vssd1 vccd1 vccd1 _25984_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _14525_/A hold191/X vssd1 vssd1 vccd1 vccd1 hold192/A sky130_fd_sc_hd__nand2_1
XFILLER_0_187_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23669_ _23669_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23670_/A sky130_fd_sc_hd__and2_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ _16210_/A _16214_/B vssd1 vssd1 vccd1 vccd1 _16210_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_153_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25408_ _26001_/CLK _25408_/D vssd1 vssd1 vccd1 vccd1 _25408_/Q sky130_fd_sc_hd__dfxtp_1
X_13422_ _13220_/A _14666_/A _13242_/X _19830_/A vssd1 vssd1 vccd1 vccd1 _13422_/X
+ sky130_fd_sc_hd__a22o_1
X_17190_ _17272_/A _17190_/B vssd1 vssd1 vccd1 vccd1 _17190_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_148_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16141_ _16135_/Y _16132_/Y _16156_/A vssd1 vssd1 vccd1 vccd1 _16150_/A sky130_fd_sc_hd__a21o_1
X_13353_ _13353_/A vssd1 vssd1 vccd1 vccd1 _19673_/A sky130_fd_sc_hd__clkbuf_8
X_25339_ _26298_/CLK hold271/X vssd1 vssd1 vccd1 vccd1 hold269/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16072_ _16084_/B _16073_/A vssd1 vssd1 vccd1 vccd1 _16072_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13284_ _26311_/Q _19518_/A vssd1 vssd1 vccd1 vccd1 _14599_/A sky130_fd_sc_hd__xor2_1
X_15023_ _15024_/B _15024_/A vssd1 vssd1 vccd1 vccd1 _15023_/X sky130_fd_sc_hd__or2_1
X_19900_ _19901_/B _19901_/A vssd1 vssd1 vccd1 vccd1 _19900_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19831_ _20672_/A _22539_/B _25638_/Q vssd1 vssd1 vccd1 vccd1 _20677_/C sky130_fd_sc_hd__nand3_1
X_19762_ _19763_/B _19763_/A vssd1 vssd1 vccd1 vccd1 _19762_/X sky130_fd_sc_hd__or2_1
X_16974_ _16974_/A _16974_/B vssd1 vssd1 vccd1 vccd1 _16974_/Y sky130_fd_sc_hd__nand2_1
X_18713_ _18955_/A _18713_/B _18894_/C vssd1 vssd1 vccd1 vccd1 _18714_/C sky130_fd_sc_hd__nand3_1
X_15925_ _15925_/A _15925_/B vssd1 vssd1 vccd1 vccd1 _15934_/A sky130_fd_sc_hd__nand2_1
X_19693_ _19691_/X _19692_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19693_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15856_ _15856_/A _15856_/B vssd1 vssd1 vccd1 vccd1 _15869_/A sky130_fd_sc_hd__nand2_1
X_18644_ _22348_/B _25630_/Q vssd1 vssd1 vccd1 vccd1 _18646_/A sky130_fd_sc_hd__nand2_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14807_ _14813_/B _22116_/A vssd1 vssd1 vccd1 vccd1 _22115_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_87_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15787_ _15787_/A _15823_/A vssd1 vssd1 vccd1 vccd1 _15789_/A sky130_fd_sc_hd__nand2_1
X_18575_ _18778_/A _18919_/A vssd1 vssd1 vccd1 vccd1 _18576_/B sky130_fd_sc_hd__xnor2_1
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999_ _26133_/Q _12907_/X _12998_/X vssd1 vssd1 vccd1 vccd1 _12999_/X sky130_fd_sc_hd__a21o_1
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14738_ _25842_/Q _13466_/A _14737_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14739_/A
+ sky130_fd_sc_hd__a22o_1
X_17526_ _17526_/A _17577_/A vssd1 vssd1 vccd1 vccd1 _17527_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17457_ _17624_/A _17457_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17457_/X sky130_fd_sc_hd__and3_1
X_14669_ _14669_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _14669_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16408_ _16473_/A hold966/X vssd1 vssd1 vccd1 vccd1 _16408_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17388_ _25618_/Q vssd1 vssd1 vccd1 vccd1 _21238_/B sky130_fd_sc_hd__inv_2
X_16339_ _16361_/A _16340_/A vssd1 vssd1 vccd1 vccd1 _16341_/A sky130_fd_sc_hd__or2_1
X_19127_ _19186_/A hold668/X vssd1 vssd1 vccd1 vccd1 hold669/A sky130_fd_sc_hd__nand2_1
XFILLER_0_172_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19058_ _19056_/Y _19057_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25705_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_164_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18009_ _18007_/X _17528_/X _18008_/X vssd1 vssd1 vccd1 vccd1 _18010_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_61_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21020_ _21018_/Y _21019_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _21020_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_168_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22971_ _23197_/A _22971_/B vssd1 vssd1 vccd1 vccd1 _22971_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24710_ hold2686/X hold2578/X _24740_/S vssd1 vssd1 vccd1 vccd1 _24711_/A sky130_fd_sc_hd__mux2_1
X_21922_ _22187_/A _23136_/A vssd1 vssd1 vccd1 vccd1 _21928_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_184_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25690_ _26324_/CLK _25690_/D vssd1 vssd1 vccd1 vccd1 _25690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24641_ _24641_/A vssd1 vssd1 vccd1 vccd1 _26276_/D sky130_fd_sc_hd__clkbuf_1
X_21853_ _22128_/A _23104_/A vssd1 vssd1 vccd1 vccd1 _21859_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20804_ _21416_/C _21692_/B vssd1 vssd1 vccd1 vccd1 _20806_/A sky130_fd_sc_hd__nand2_1
X_24572_ _26253_/Q hold2727/X _24587_/S vssd1 vssd1 vccd1 vccd1 _24572_/X sky130_fd_sc_hd__mux2_1
X_21784_ _21784_/A _21784_/B vssd1 vssd1 vccd1 vccd1 _21786_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_72_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26311_ _26313_/CLK _26311_/D vssd1 vssd1 vccd1 vccd1 _26311_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_93_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23523_ _24944_/S hold359/A _23522_/X vssd1 vssd1 vccd1 vccd1 _23523_/Y sky130_fd_sc_hd__o21ai_1
X_20735_ _21042_/A _20735_/B _20734_/X vssd1 vssd1 vccd1 vccd1 _20736_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_175_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26242_ _26244_/CLK _26242_/D vssd1 vssd1 vccd1 vccd1 _26242_/Q sky130_fd_sc_hd__dfxtp_2
X_23454_ _24922_/S hold239/A _23453_/X vssd1 vssd1 vccd1 vccd1 _23454_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_162_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20666_ _25855_/Q _20666_/B _20666_/C vssd1 vssd1 vccd1 vccd1 _20669_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_73_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22405_ _22561_/A _22405_/B vssd1 vssd1 vccd1 vccd1 _22405_/Y sky130_fd_sc_hd__nand2_1
X_26173_ _26175_/CLK _26173_/D vssd1 vssd1 vccd1 vccd1 _26173_/Q sky130_fd_sc_hd__dfxtp_1
X_20597_ _20597_/A _20597_/B vssd1 vssd1 vccd1 vccd1 _20601_/A sky130_fd_sc_hd__nand2_1
X_23385_ _24942_/S hold263/A _23384_/X vssd1 vssd1 vccd1 vccd1 _23385_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25124_ _25708_/CLK _25124_/D vssd1 vssd1 vccd1 vccd1 _25124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22336_ _22774_/B _22924_/A vssd1 vssd1 vccd1 vccd1 _22338_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25055_ _26142_/CLK _25055_/D vssd1 vssd1 vccd1 vccd1 _25055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22267_ _25819_/Q _22267_/B vssd1 vssd1 vccd1 vccd1 _22267_/Y sky130_fd_sc_hd__nor2_1
X_24006_ _24006_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24007_/A sky130_fd_sc_hd__and2_1
XFILLER_0_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21218_ _21218_/A _21218_/B vssd1 vssd1 vccd1 vccd1 _21659_/C sky130_fd_sc_hd__nand2_4
X_22198_ _22198_/A _23122_/A _22198_/C vssd1 vssd1 vccd1 vccd1 _22198_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_178_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21149_ _21148_/Y _20192_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21149_/X
+ sky130_fd_sc_hd__a211o_1
X_25957_ _26023_/CLK _25957_/D vssd1 vssd1 vccd1 vccd1 _25957_/Q sky130_fd_sc_hd__dfxtp_1
X_13971_ _26293_/Q _13801_/X _13793_/X _13970_/Y vssd1 vssd1 vccd1 vccd1 _13972_/B
+ sky130_fd_sc_hd__a22o_1
X_15710_ _16617_/A _15778_/B vssd1 vssd1 vccd1 vccd1 _16937_/A sky130_fd_sc_hd__nand2_2
X_24908_ _24908_/A _24959_/A vssd1 vssd1 vccd1 vccd1 _24908_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_38_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12922_ _26118_/Q _12907_/X _12921_/X vssd1 vssd1 vccd1 vccd1 _12922_/X sky130_fd_sc_hd__a21o_1
X_16690_ hold575/X vssd1 vssd1 vccd1 vccd1 _16692_/A sky130_fd_sc_hd__inv_2
XFILLER_0_88_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25888_ _26080_/CLK _25888_/D vssd1 vssd1 vccd1 vccd1 _25888_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_77_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15641_ _15641_/A _15641_/B vssd1 vssd1 vccd1 vccd1 _15693_/C sky130_fd_sc_hd__nor2_1
X_24839_ _15160_/A _15177_/B _24860_/S vssd1 vssd1 vccd1 vccd1 _24839_/X sky130_fd_sc_hd__mux2_1
X_12853_ _26105_/Q _12748_/X _12852_/X vssd1 vssd1 vccd1 vccd1 _12853_/X sky130_fd_sc_hd__a21o_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _21184_/B _19518_/A vssd1 vssd1 vccd1 vccd1 _18361_/B sky130_fd_sc_hd__nand2_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _15572_/A _15572_/B vssd1 vssd1 vccd1 vccd1 _15577_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_115_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _12726_/B _14310_/A _12752_/X _25589_/Q vssd1 vssd1 vccd1 vccd1 _12784_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _17311_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17311_/Y sky130_fd_sc_hd__nand2_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14523_ _14521_/Y hold321/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold322/A sky130_fd_sc_hd__a21oi_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18291_ _18494_/A _18637_/A vssd1 vssd1 vccd1 vccd1 _18292_/B sky130_fd_sc_hd__xnor2_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17393_/A _17242_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17242_/X sky130_fd_sc_hd__and3_1
X_14454_ _14452_/Y hold342/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold343/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13405_ hold995/X _13944_/A vssd1 vssd1 vccd1 vccd1 _13405_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17173_ _17441_/A _17173_/B vssd1 vssd1 vccd1 vccd1 _17173_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_4_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14385_ _14385_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14385_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16124_ _16124_/A _16124_/B vssd1 vssd1 vccd1 vccd1 _16134_/B sky130_fd_sc_hd__nand2_1
X_13336_ _26319_/Q _19630_/A vssd1 vssd1 vccd1 vccd1 _14623_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_12_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_5__f_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_5__f_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_161_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16055_ _16273_/C _16273_/B vssd1 vssd1 vccd1 vccd1 _16055_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_122_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13267_ _13220_/X _14589_/A _13242_/X _19473_/A vssd1 vssd1 vccd1 vccd1 _13267_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15006_ _15006_/A _15006_/B vssd1 vssd1 vccd1 vccd1 _15007_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13198_ _26169_/Q _13065_/X _13197_/X vssd1 vssd1 vccd1 vccd1 _13198_/X sky130_fd_sc_hd__a21o_1
X_19814_ _19813_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19815_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1709 _22638_/Y vssd1 vssd1 vccd1 vccd1 _25869_/D sky130_fd_sc_hd__dlygate4sd3_1
X_19745_ _20438_/A _22391_/B _25632_/Q vssd1 vssd1 vccd1 vccd1 _20443_/C sky130_fd_sc_hd__nand3_1
X_16957_ _16955_/Y _16956_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _16957_/Y sky130_fd_sc_hd__a21oi_1
X_15908_ _15908_/A _15908_/B vssd1 vssd1 vccd1 vccd1 _15921_/A sky130_fd_sc_hd__nand2_1
X_19676_ _19692_/B _19763_/B vssd1 vssd1 vccd1 vccd1 _19678_/A sky130_fd_sc_hd__xnor2_1
X_16888_ _16935_/A _16893_/B vssd1 vssd1 vccd1 vccd1 _16890_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_188_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18627_ _25885_/Q _22326_/A vssd1 vssd1 vccd1 vccd1 _18635_/A sky130_fd_sc_hd__or2_2
X_15839_ _15839_/A _15839_/B vssd1 vssd1 vccd1 vccd1 _15840_/A sky130_fd_sc_hd__nand2_1
X_18558_ _18555_/X _18269_/X _18557_/X vssd1 vssd1 vccd1 vccd1 _18559_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_118_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17509_ _17509_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17509_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_157_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18489_ _18955_/A _18489_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18490_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_74_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_13 _23496_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20520_ _20520_/A _25890_/Q vssd1 vssd1 vccd1 vccd1 _20526_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_24 _19017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_35 _26213_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_57 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20451_ _21546_/A _21249_/C vssd1 vssd1 vccd1 vccd1 _20452_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_133_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_68 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_79 _25837_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23170_ _23170_/A _23170_/B vssd1 vssd1 vccd1 vccd1 _23171_/A sky130_fd_sc_hd__xor2_1
X_20382_ _26286_/Q hold536/X vssd1 vssd1 vccd1 vccd1 _20382_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22121_ _18492_/A _25814_/Q _22119_/Y _22120_/Y vssd1 vssd1 vccd1 vccd1 _22122_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22052_ _18189_/B _25591_/Q _18191_/A vssd1 vssd1 vccd1 vccd1 _22053_/B sky130_fd_sc_hd__o21ai_2
X_21003_ _21003_/A _21003_/B vssd1 vssd1 vccd1 vccd1 _21529_/C sky130_fd_sc_hd__nand2_4
X_25811_ _25812_/CLK _25811_/D vssd1 vssd1 vccd1 vccd1 _25811_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_138_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25742_ _25745_/CLK _25742_/D vssd1 vssd1 vccd1 vccd1 _25742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22954_ _23197_/A _22954_/B vssd1 vssd1 vccd1 vccd1 _22954_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21905_ _18141_/A _25798_/Q _21903_/Y _21904_/Y vssd1 vssd1 vccd1 vccd1 _21906_/B
+ sky130_fd_sc_hd__a31o_1
X_25673_ _26303_/CLK _25673_/D vssd1 vssd1 vccd1 vccd1 _25673_/Q sky130_fd_sc_hd__dfxtp_1
X_22885_ _16851_/B _22421_/X _22879_/X _22880_/Y _22884_/X vssd1 vssd1 vccd1 vccd1
+ _22886_/A sky130_fd_sc_hd__a221o_1
X_24624_ hold2705/X hold2634/X _24664_/S vssd1 vssd1 vccd1 vccd1 _24625_/A sky130_fd_sc_hd__mux2_1
X_21836_ _18055_/A _25796_/Q _21834_/Y _21835_/Y vssd1 vssd1 vccd1 vccd1 _21837_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24555_ _24555_/A vssd1 vssd1 vccd1 vccd1 _26248_/D sky130_fd_sc_hd__clkbuf_1
X_21767_ _19317_/A _21766_/A _21766_/Y vssd1 vssd1 vccd1 vccd1 _21769_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23506_ _23503_/Y _23505_/Y _24946_/A vssd1 vssd1 vccd1 vccd1 _23506_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20718_ _20720_/B vssd1 vssd1 vccd1 vccd1 _20719_/B sky130_fd_sc_hd__inv_2
XFILLER_0_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24486_ hold2653/X hold2555/X _24510_/S vssd1 vssd1 vccd1 vccd1 _24487_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_135_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21698_ _26339_/Q hold431/X vssd1 vssd1 vccd1 vccd1 _21698_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_93_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26225_ _26226_/CLK _26225_/D vssd1 vssd1 vccd1 vccd1 _26225_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_163_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23437_ _24922_/S hold353/A _23436_/X vssd1 vssd1 vccd1 vccd1 _23437_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20649_ _21354_/B _21628_/B vssd1 vssd1 vccd1 vccd1 _20651_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_184_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14170_ _14170_/A vssd1 vssd1 vccd1 vccd1 _14170_/X sky130_fd_sc_hd__clkbuf_16
X_26156_ _26284_/CLK _26156_/D vssd1 vssd1 vccd1 vccd1 _26156_/Q sky130_fd_sc_hd__dfxtp_1
X_23368_ _23368_/A vssd1 vssd1 vccd1 vccd1 _25936_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13121_ _13049_/X _14512_/A _13067_/X _25653_/Q vssd1 vssd1 vccd1 vccd1 _13121_/X
+ sky130_fd_sc_hd__a22o_1
X_25107_ _26190_/CLK _25107_/D vssd1 vssd1 vccd1 vccd1 _25107_/Q sky130_fd_sc_hd__dfxtp_1
X_22319_ _22295_/X _22318_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _22319_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26087_ _26089_/CLK _26087_/D vssd1 vssd1 vccd1 vccd1 _26087_/Q sky130_fd_sc_hd__dfxtp_1
X_23299_ _23301_/A _23377_/B _23299_/C vssd1 vssd1 vccd1 vccd1 _23300_/A sky130_fd_sc_hd__and3_1
XFILLER_0_30_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25038_ _25135_/CLK _25038_/D vssd1 vssd1 vccd1 vccd1 _25038_/Q sky130_fd_sc_hd__dfxtp_1
X_13052_ _26143_/Q _12907_/X _13051_/X vssd1 vssd1 vccd1 vccd1 _13052_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17860_ _20434_/B _17860_/B vssd1 vssd1 vccd1 vccd1 _20428_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_100_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16811_ _16809_/X _16711_/X _16810_/Y _25876_/Q _14170_/X vssd1 vssd1 vccd1 vccd1
+ _16812_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17791_ _18098_/A vssd1 vssd1 vccd1 vccd1 _18611_/A sky130_fd_sc_hd__buf_12
Xclkbuf_4_13__f_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_95_clk/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19530_ _19529_/Y _19272_/X _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19531_/B
+ sky130_fd_sc_hd__a211o_1
X_16742_ _16742_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16742_/Y sky130_fd_sc_hd__nand2_1
X_13954_ _14061_/A _13954_/B vssd1 vssd1 vccd1 vccd1 _13954_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12905_ _17404_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12905_/X sky130_fd_sc_hd__or2_1
X_16673_ _16698_/A hold689/X vssd1 vssd1 vccd1 vccd1 hold690/A sky130_fd_sc_hd__nand2_1
X_19461_ _19478_/B _19551_/B vssd1 vssd1 vccd1 vccd1 _19463_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_194_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _26119_/CLK sky130_fd_sc_hd__clkbuf_16
X_13885_ _13941_/A _13885_/B vssd1 vssd1 vccd1 vccd1 _13885_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_186_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18412_ _18617_/A _18758_/A vssd1 vssd1 vccd1 vccd1 _18413_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15624_ _15624_/A vssd1 vssd1 vccd1 vccd1 _16904_/A sky130_fd_sc_hd__inv_2
XFILLER_0_154_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12836_ _12726_/B _14340_/A _12752_/X _25599_/Q vssd1 vssd1 vccd1 vccd1 _12836_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19392_ _19393_/B _19393_/A vssd1 vssd1 vccd1 vccd1 _19392_/X sky130_fd_sc_hd__or2_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15555_ _15551_/A _15504_/Y _15554_/Y vssd1 vssd1 vccd1 vccd1 _15555_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_139_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18343_ _18445_/A _18347_/B vssd1 vssd1 vccd1 vccd1 _18345_/A sky130_fd_sc_hd__nand2_1
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12767_ _12746_/X _12765_/X _14910_/B _12766_/X vssd1 vssd1 vccd1 vccd1 hold989/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _14506_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14506_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_189_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18274_ _18641_/A _19206_/A vssd1 vssd1 vccd1 vccd1 _18274_/Y sky130_fd_sc_hd__nand2_1
X_15486_ _15486_/A vssd1 vssd1 vccd1 vccd1 _15495_/B sky130_fd_sc_hd__inv_2
XFILLER_0_126_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12698_ _12698_/A vssd1 vssd1 vccd1 vccd1 _24991_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17225_ _17520_/A _17600_/A vssd1 vssd1 vccd1 vccd1 _17226_/B sky130_fd_sc_hd__xnor2_1
X_14437_ _14437_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14437_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17156_ _25633_/Q vssd1 vssd1 vccd1 vccd1 _20479_/B sky130_fd_sc_hd__inv_2
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14368_ _14404_/A hold83/X vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold806 hold806/A vssd1 vssd1 vccd1 vccd1 hold806/X sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ _16107_/A vssd1 vssd1 vccd1 vccd1 _16107_/Y sky130_fd_sc_hd__inv_2
Xhold817 hold817/A vssd1 vssd1 vccd1 vccd1 hold817/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 hold828/A vssd1 vssd1 vccd1 vccd1 hold828/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13319_ _26188_/Q _13239_/X _13318_/X vssd1 vssd1 vccd1 vccd1 _13319_/X sky130_fd_sc_hd__a21o_1
X_17087_ _19206_/A _17087_/B vssd1 vssd1 vccd1 vccd1 _17448_/A sky130_fd_sc_hd__xor2_4
Xhold839 hold839/A vssd1 vssd1 vccd1 vccd1 hold839/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_110_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14299_ _14344_/A hold182/X vssd1 vssd1 vccd1 vccd1 hold183/A sky130_fd_sc_hd__nand2_1
X_16038_ _16038_/A _16038_/B vssd1 vssd1 vccd1 vccd1 _16039_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2207 _14959_/Y vssd1 vssd1 vccd1 vccd1 hold2207/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2218 _26099_/Q vssd1 vssd1 vccd1 vccd1 hold2218/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2229 _12652_/X vssd1 vssd1 vccd1 vccd1 _12653_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1506 _13264_/X vssd1 vssd1 vccd1 vccd1 _25096_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1517 _25643_/Q vssd1 vssd1 vccd1 vccd1 _17642_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17989_ _18529_/A _17989_/B _18529_/C vssd1 vssd1 vccd1 vccd1 _17990_/C sky130_fd_sc_hd__nand3_1
Xhold1528 _19383_/Y vssd1 vssd1 vccd1 vccd1 _25728_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1539 _25725_/Q vssd1 vssd1 vccd1 vccd1 _19339_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19728_ _19725_/Y _19728_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19728_/X sky130_fd_sc_hd__and3b_1
X_19659_ _19659_/A _20200_/B vssd1 vssd1 vccd1 vccd1 _19659_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_185_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _25745_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22670_ _22670_/A _22670_/B vssd1 vssd1 vccd1 vccd1 _22671_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_176_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21621_ _21621_/A _21621_/B vssd1 vssd1 vccd1 vccd1 _21622_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_176_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xascon_wrapper_19 vssd1 vssd1 vccd1 vccd1 io_oeb[5] ascon_wrapper_19/LO sky130_fd_sc_hd__conb_1
XFILLER_0_117_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24340_ _24340_/A vssd1 vssd1 vccd1 vccd1 _26178_/D sky130_fd_sc_hd__clkbuf_1
X_21552_ _26330_/Q hold783/X vssd1 vssd1 vccd1 vccd1 _21552_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_28_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20503_ _20503_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _20503_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_62_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24271_ _24271_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24272_/A sky130_fd_sc_hd__and2_1
XFILLER_0_145_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21483_ _21483_/A _21483_/B _21483_/C vssd1 vssd1 vccd1 vccd1 _21484_/B sky130_fd_sc_hd__nand3_1
X_26010_ _26012_/CLK _26010_/D vssd1 vssd1 vccd1 vccd1 _26010_/Q sky130_fd_sc_hd__dfxtp_1
X_23222_ _23222_/A _24863_/S vssd1 vssd1 vccd1 vccd1 _23253_/C sky130_fd_sc_hd__nand2_1
X_20434_ _20434_/A _20434_/B vssd1 vssd1 vccd1 vccd1 _20436_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23153_ _23153_/A _23153_/B vssd1 vssd1 vccd1 vccd1 _23154_/B sky130_fd_sc_hd__nand2_1
X_20365_ _22954_/B vssd1 vssd1 vccd1 vccd1 _22353_/B sky130_fd_sc_hd__inv_2
XFILLER_0_113_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22104_ _22601_/A _22791_/B vssd1 vssd1 vccd1 vccd1 _22110_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_140_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23084_ _23075_/Y _23083_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _23084_/X sky130_fd_sc_hd__a21o_1
X_20296_ _20298_/A _20298_/B vssd1 vssd1 vccd1 vccd1 _20297_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_140_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22035_ _22653_/A _22035_/B vssd1 vssd1 vccd1 vccd1 _22035_/X sky130_fd_sc_hd__or2_1
Xhold2730 _26313_/Q vssd1 vssd1 vccd1 vccd1 hold2730/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2741 _25258_/Q vssd1 vssd1 vccd1 vccd1 _12483_/A sky130_fd_sc_hd__buf_1
Xhold2752 _25509_/Q vssd1 vssd1 vccd1 vccd1 hold863/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23986_ hold2466/X hold2418/X _24001_/S vssd1 vssd1 vccd1 vccd1 _23987_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25725_ _25729_/CLK _25725_/D vssd1 vssd1 vccd1 vccd1 _25725_/Q sky130_fd_sc_hd__dfxtp_1
X_22937_ _22937_/A _22937_/B vssd1 vssd1 vccd1 vccd1 _22937_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_176_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _25785_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_151_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25656_ _25797_/CLK _25656_/D vssd1 vssd1 vccd1 vccd1 _25656_/Q sky130_fd_sc_hd__dfxtp_2
X_13670_ _18327_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13670_/Y sky130_fd_sc_hd__nor2_1
X_22868_ _22868_/A _23001_/B _22868_/C vssd1 vssd1 vccd1 vccd1 _22868_/X sky130_fd_sc_hd__and3_1
XFILLER_0_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ _12621_/A vssd1 vssd1 vccd1 vccd1 _12645_/B sky130_fd_sc_hd__clkinvlp_2
X_24607_ _24607_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24608_/A sky130_fd_sc_hd__and2_1
XFILLER_0_183_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21819_ _22103_/A _23088_/A vssd1 vssd1 vccd1 vccd1 _21825_/B sky130_fd_sc_hd__nand2_1
X_25587_ _25587_/CLK _25587_/D vssd1 vssd1 vccd1 vccd1 _25587_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22799_ _22799_/A _22799_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22801_/A sky130_fd_sc_hd__or3_1
XFILLER_0_149_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15340_ _15340_/A vssd1 vssd1 vccd1 vccd1 _16796_/A sky130_fd_sc_hd__inv_2
XFILLER_0_183_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24538_ hold2657/X _26243_/Q _24587_/S vssd1 vssd1 vccd1 vccd1 _24538_/X sky130_fd_sc_hd__mux2_1
X_12552_ _25904_/Q _25903_/Q vssd1 vssd1 vccd1 vccd1 _17748_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15271_ _15272_/B _15271_/B vssd1 vssd1 vccd1 vccd1 _15271_/X sky130_fd_sc_hd__and2_1
XFILLER_0_184_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12483_ _12483_/A vssd1 vssd1 vccd1 vccd1 _15773_/S sky130_fd_sc_hd__buf_12
X_24469_ _24469_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24470_/A sky130_fd_sc_hd__and2_1
XFILLER_0_164_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17010_ _23199_/A vssd1 vssd1 vccd1 vccd1 _21791_/A sky130_fd_sc_hd__clkbuf_16
X_26208_ _26208_/CLK _26208_/D vssd1 vssd1 vccd1 vccd1 _26208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14222_ _14264_/A _14222_/B vssd1 vssd1 vccd1 vccd1 _14222_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_34_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26139_ _26139_/CLK _26139_/D vssd1 vssd1 vccd1 vccd1 _26139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14153_ _26322_/Q _13988_/X _13981_/X _14152_/Y vssd1 vssd1 vccd1 vccd1 _14154_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_100_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _25925_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_132_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13104_ _26281_/Q _25650_/Q vssd1 vssd1 vccd1 vccd1 _14503_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_42_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14084_ _18368_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14084_/Y sky130_fd_sc_hd__nor2_1
X_18961_ _19026_/A _18961_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18961_/X sky130_fd_sc_hd__and3_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17912_ _19052_/A _18413_/A vssd1 vssd1 vccd1 vccd1 _17913_/B sky130_fd_sc_hd__xnor2_4
X_13035_ _12891_/X _14461_/A _12909_/X _25637_/Q vssd1 vssd1 vccd1 vccd1 _13035_/X
+ sky130_fd_sc_hd__a22o_1
X_18892_ _18892_/A _25834_/Q _18892_/C vssd1 vssd1 vccd1 vccd1 _20835_/B sky130_fd_sc_hd__nand3_2
X_17843_ _18612_/A _25728_/Q _18083_/C vssd1 vssd1 vccd1 vccd1 _17844_/C sky130_fd_sc_hd__nand3_1
X_17774_ _17781_/A _17774_/B _17830_/A vssd1 vssd1 vccd1 vccd1 _17775_/C sky130_fd_sc_hd__nand3_4
X_14986_ _14986_/A _14998_/A vssd1 vssd1 vccd1 vccd1 _14986_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19513_ _19511_/Y _19512_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19513_/Y sky130_fd_sc_hd__a21oi_1
X_16725_ _16726_/B _16726_/A vssd1 vssd1 vccd1 vccd1 _16725_/X sky130_fd_sc_hd__or2_1
XFILLER_0_88_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13937_ _14000_/A hold485/X vssd1 vssd1 vccd1 vccd1 hold486/A sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_167_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _26287_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_135_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19444_ _19444_/A _21048_/B vssd1 vssd1 vccd1 vccd1 _19444_/Y sky130_fd_sc_hd__nor2_1
X_16656_ _16656_/A _16669_/A vssd1 vssd1 vccd1 vccd1 _16659_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13868_ _13880_/A hold722/X vssd1 vssd1 vccd1 vccd1 hold723/A sky130_fd_sc_hd__nand2_1
X_15607_ _15579_/X _15612_/A _15590_/B vssd1 vssd1 vccd1 vccd1 _15609_/A sky130_fd_sc_hd__a21o_1
X_12819_ _12726_/B _14331_/A _12752_/X _25596_/Q vssd1 vssd1 vccd1 vccd1 _12819_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19375_ _20908_/A _19373_/Y _20913_/C vssd1 vssd1 vccd1 vccd1 _19463_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_186_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16587_ _16587_/A _16587_/B vssd1 vssd1 vccd1 vccd1 _16588_/B sky130_fd_sc_hd__and2_1
XFILLER_0_146_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13799_ hold734/X _13797_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold735/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18326_ _18951_/A _25742_/Q vssd1 vssd1 vccd1 vccd1 _18328_/A sky130_fd_sc_hd__nand2_1
X_15538_ _26029_/Q _25965_/Q _15773_/S vssd1 vssd1 vccd1 vccd1 _15539_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_151_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15469_ _15467_/A _15446_/B _15468_/Y vssd1 vssd1 vccd1 vccd1 _15469_/Y sky130_fd_sc_hd__o21ai_1
X_18257_ _18257_/A _18257_/B vssd1 vssd1 vccd1 vccd1 _21772_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_167_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17208_ _19331_/A _17208_/B vssd1 vssd1 vccd1 vccd1 _17513_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18188_ _18190_/A _18190_/C vssd1 vssd1 vccd1 vccd1 _18189_/A sky130_fd_sc_hd__nand2_1
Xhold603 hold603/A vssd1 vssd1 vccd1 vccd1 hold603/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17139_ _17137_/Y _17138_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _17139_/Y sky130_fd_sc_hd__a21oi_1
Xhold614 hold614/A vssd1 vssd1 vccd1 vccd1 hold614/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold625 hold625/A vssd1 vssd1 vccd1 vccd1 hold625/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold636 hold636/A vssd1 vssd1 vccd1 vccd1 hold636/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 hold647/A vssd1 vssd1 vccd1 vccd1 hold647/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 hold658/A vssd1 vssd1 vccd1 vccd1 hold658/X sky130_fd_sc_hd__dlygate4sd3_1
X_20150_ _20150_/A _20949_/C vssd1 vssd1 vccd1 vccd1 _20152_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold669 hold669/A vssd1 vssd1 vccd1 vccd1 hold669/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20081_ _20080_/Y _21228_/A _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20081_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2004 _26146_/Q vssd1 vssd1 vccd1 vccd1 hold2004/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2015 _12640_/X vssd1 vssd1 vccd1 vccd1 _12641_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2026 _23742_/X vssd1 vssd1 vccd1 vccd1 _23743_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2037 _26171_/Q vssd1 vssd1 vccd1 vccd1 hold2037/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2048 _26037_/Q vssd1 vssd1 vccd1 vccd1 hold2048/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1303 _13043_/X vssd1 vssd1 vccd1 vccd1 _25058_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1314 _25556_/Q vssd1 vssd1 vccd1 vccd1 _16820_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2059 _25989_/Q vssd1 vssd1 vccd1 vccd1 _14770_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1325 _25802_/Q vssd1 vssd1 vccd1 vccd1 _21045_/B sky130_fd_sc_hd__clkbuf_2
Xhold1336 _20623_/Y vssd1 vssd1 vccd1 vccd1 _25789_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23840_ _23840_/A vssd1 vssd1 vccd1 vccd1 _26017_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1347 _25020_/Q vssd1 vssd1 vccd1 vccd1 _17269_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1358 _13226_/X vssd1 vssd1 vccd1 vccd1 _25090_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1369 _25410_/Q vssd1 vssd1 vccd1 vccd1 _14891_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23771_ _23771_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23772_/A sky130_fd_sc_hd__and2_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_158_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _26164_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20983_ _20983_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _20989_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_170_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25510_ _25510_/CLK hold959/X vssd1 vssd1 vccd1 vccd1 hold958/A sky130_fd_sc_hd__dfxtp_1
X_22722_ _22723_/B _22723_/A vssd1 vssd1 vccd1 vccd1 _22724_/A sky130_fd_sc_hd__or2_1
XFILLER_0_79_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25441_ _25501_/CLK _25441_/D vssd1 vssd1 vccd1 vccd1 _25441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22653_ _22653_/A _22653_/B vssd1 vssd1 vccd1 vccd1 _22653_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21604_ _21604_/A _21604_/B vssd1 vssd1 vccd1 vccd1 _21605_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25372_ _26193_/CLK hold34/X vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__dfxtp_1
X_22584_ _22584_/A _22900_/B vssd1 vssd1 vccd1 vccd1 _22584_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_69_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24323_ hold2384/X _26173_/Q _24356_/S vssd1 vssd1 vccd1 vccd1 _24323_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_161_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21535_ _26329_/Q _19130_/X hold827/X vssd1 vssd1 vccd1 vccd1 _21538_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24254_ _24254_/A vssd1 vssd1 vccd1 vccd1 _26150_/D sky130_fd_sc_hd__clkbuf_1
X_21466_ _21466_/A _21515_/A vssd1 vssd1 vccd1 vccd1 _21467_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_69_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23205_ _23212_/A _23205_/B vssd1 vssd1 vccd1 vccd1 _23206_/A sky130_fd_sc_hd__nand2_1
X_20417_ _20417_/A _21144_/B _20417_/C vssd1 vssd1 vccd1 vccd1 _20418_/B sky130_fd_sc_hd__nand3_1
X_24185_ _24185_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24186_/A sky130_fd_sc_hd__and2_1
XFILLER_0_120_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21397_ _21395_/Y _21396_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21397_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23136_ _23136_/A _23136_/B vssd1 vssd1 vccd1 vccd1 _23137_/B sky130_fd_sc_hd__nand2_1
X_20348_ _20346_/Y _20347_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _20348_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23067_ _23067_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _23067_/Y sky130_fd_sc_hd__nand2_1
X_20279_ _20281_/B vssd1 vssd1 vccd1 vccd1 _20280_/B sky130_fd_sc_hd__inv_2
XFILLER_0_179_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22018_ _19546_/A _22017_/A _22017_/Y vssd1 vssd1 vccd1 vccd1 _22020_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_175_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2560 _24501_/X vssd1 vssd1 vccd1 vccd1 _24502_/A sky130_fd_sc_hd__dlygate4sd3_1
X_14840_ _14900_/A hold955/X vssd1 vssd1 vccd1 vccd1 _14840_/Y sky130_fd_sc_hd__nand2_1
Xhold2571 _26232_/Q vssd1 vssd1 vccd1 vccd1 hold2571/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2582 _26250_/Q vssd1 vssd1 vccd1 vccd1 hold2582/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2593 _24458_/X vssd1 vssd1 vccd1 vccd1 _24459_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1870 _25855_/Q vssd1 vssd1 vccd1 vccd1 _22290_/B sky130_fd_sc_hd__dlygate4sd3_1
X_14771_ _14777_/B _22002_/A vssd1 vssd1 vccd1 vccd1 _22001_/B sky130_fd_sc_hd__xnor2_2
Xhold1881 _22000_/Y vssd1 vssd1 vccd1 vccd1 _25845_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23969_ _23969_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23970_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_149_clk clkbuf_4_11__f_clk/X vssd1 vssd1 vccd1 vccd1 _26308_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1892 _24332_/X vssd1 vssd1 vccd1 vccd1 _24333_/A sky130_fd_sc_hd__dlygate4sd3_1
X_16510_ _16510_/A hold940/X _16691_/B vssd1 vssd1 vccd1 vccd1 _16511_/B sky130_fd_sc_hd__and3_1
X_13722_ _13823_/A _13722_/B vssd1 vssd1 vccd1 vccd1 _13722_/Y sky130_fd_sc_hd__nand2_1
X_25708_ _25708_/CLK _25708_/D vssd1 vssd1 vccd1 vccd1 _25708_/Q sky130_fd_sc_hd__dfxtp_4
X_17490_ _17488_/Y _17489_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _17490_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_168_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16441_ _16441_/A _16441_/B vssd1 vssd1 vccd1 vccd1 _16442_/B sky130_fd_sc_hd__nor2_1
X_13653_ _26242_/Q _13612_/X _13605_/X _13652_/Y vssd1 vssd1 vccd1 vccd1 _13654_/B
+ sky130_fd_sc_hd__a22o_1
X_25639_ _26252_/CLK _25639_/D vssd1 vssd1 vccd1 vccd1 _25639_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12604_ _12643_/B _12610_/A vssd1 vssd1 vccd1 vccd1 _12606_/A sky130_fd_sc_hd__or2_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16372_ _16370_/Y _16372_/B vssd1 vssd1 vccd1 vccd1 _16378_/B sky130_fd_sc_hd__and2b_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19160_ _20174_/B _20174_/A vssd1 vssd1 vccd1 vccd1 _20175_/A sky130_fd_sc_hd__or2_1
XFILLER_0_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13584_ hold465/X _13583_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold466/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ _15326_/A _15324_/A vssd1 vssd1 vccd1 vccd1 _15323_/X sky130_fd_sc_hd__or2_1
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ input7/X vssd1 vssd1 vccd1 vccd1 _21099_/A sky130_fd_sc_hd__buf_12
XFILLER_0_171_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12535_ _12535_/A _15839_/B vssd1 vssd1 vccd1 vccd1 _15795_/A sky130_fd_sc_hd__nand2_8
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19091_ _19089_/A _19088_/Y _20024_/A vssd1 vssd1 vccd1 vccd1 _19990_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15254_ _16771_/B vssd1 vssd1 vccd1 vccd1 _22656_/B sky130_fd_sc_hd__inv_2
XFILLER_0_124_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18042_ _25860_/Q _21834_/A vssd1 vssd1 vccd1 vccd1 _18055_/A sky130_fd_sc_hd__or2_2
XFILLER_0_163_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14205_ hold784/X _14204_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold785/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15185_ _15185_/A _15185_/B vssd1 vssd1 vccd1 vccd1 _15271_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_105_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14136_ _14180_/A _14136_/B vssd1 vssd1 vccd1 vccd1 _14136_/Y sky130_fd_sc_hd__nand2_1
X_19993_ _26276_/Q _19483_/A hold725/X vssd1 vssd1 vccd1 vccd1 _19994_/C sky130_fd_sc_hd__a21o_1
X_14067_ _26308_/Q _13988_/X _13981_/X _14066_/Y vssd1 vssd1 vccd1 vccd1 _14068_/B
+ sky130_fd_sc_hd__a22o_1
X_18944_ _18986_/A _19673_/A vssd1 vssd1 vccd1 vccd1 _18944_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13018_ _14260_/A vssd1 vssd1 vccd1 vccd1 _13018_/X sky130_fd_sc_hd__clkbuf_8
X_18875_ _20797_/B _22617_/A vssd1 vssd1 vccd1 vccd1 _20790_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_20_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17826_ _21784_/A _25583_/Q vssd1 vssd1 vccd1 vccd1 _17828_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17757_ _17875_/B _17757_/B vssd1 vssd1 vccd1 vccd1 _17924_/A sky130_fd_sc_hd__nand2_1
X_14969_ _15033_/A _14982_/B vssd1 vssd1 vccd1 vccd1 _14969_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16708_ _22680_/A vssd1 vssd1 vccd1 vccd1 _16980_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_159_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17688_ _17688_/A _17688_/B vssd1 vssd1 vccd1 vccd1 _17693_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_147_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19427_ _26235_/Q hold641/X vssd1 vssd1 vccd1 vccd1 _19427_/Y sky130_fd_sc_hd__nand2_1
X_16639_ hold920/X _16640_/A vssd1 vssd1 vccd1 vccd1 _16639_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_58_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19358_ _19355_/Y _19358_/B _19980_/B vssd1 vssd1 vccd1 vccd1 _19358_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_88_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18309_ _21109_/C _21846_/A vssd1 vssd1 vccd1 vccd1 _21101_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19289_ _19289_/A _20702_/B vssd1 vssd1 vccd1 vccd1 _19289_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_73_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21320_ _21678_/B _21369_/A vssd1 vssd1 vccd1 vccd1 _21322_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_170_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold400 hold400/A vssd1 vssd1 vccd1 vccd1 hold400/X sky130_fd_sc_hd__dlygate4sd3_1
X_21251_ _21675_/C _21630_/B vssd1 vssd1 vccd1 vccd1 _21252_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_170_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold411 hold411/A vssd1 vssd1 vccd1 vccd1 hold411/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold422 hold422/A vssd1 vssd1 vccd1 vccd1 hold422/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold433 hold433/A vssd1 vssd1 vccd1 vccd1 hold433/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20202_ _20202_/A _25882_/Q vssd1 vssd1 vccd1 vccd1 _20208_/A sky130_fd_sc_hd__nand2_1
Xhold444 hold444/A vssd1 vssd1 vccd1 vccd1 hold444/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 hold455/A vssd1 vssd1 vccd1 vccd1 hold455/X sky130_fd_sc_hd__dlygate4sd3_1
X_21182_ _21180_/Y _21181_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21182_/Y sky130_fd_sc_hd__a21oi_1
Xhold466 hold466/A vssd1 vssd1 vccd1 vccd1 hold466/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold477 hold477/A vssd1 vssd1 vccd1 vccd1 hold477/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold488 hold488/A vssd1 vssd1 vccd1 vccd1 hold488/X sky130_fd_sc_hd__dlygate4sd3_1
X_20133_ _20135_/B _20135_/C vssd1 vssd1 vccd1 vccd1 _20134_/A sky130_fd_sc_hd__nand2_1
X_25990_ _25991_/CLK _25990_/D vssd1 vssd1 vccd1 vccd1 _25990_/Q sky130_fd_sc_hd__dfxtp_1
Xhold499 hold499/A vssd1 vssd1 vccd1 vccd1 hold499/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24941_ _24946_/A _24941_/B vssd1 vssd1 vccd1 vccd1 _24941_/Y sky130_fd_sc_hd__nor2_1
X_20064_ _21692_/A _21386_/A vssd1 vssd1 vccd1 vccd1 _20072_/A sky130_fd_sc_hd__nand2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1100 _16901_/Y vssd1 vssd1 vccd1 vccd1 _25568_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 _25541_/Q vssd1 vssd1 vccd1 vccd1 _16715_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 _13457_/X vssd1 vssd1 vccd1 vccd1 _25128_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24872_ _15996_/B _16011_/A _24956_/S vssd1 vssd1 vccd1 vccd1 _24873_/A sky130_fd_sc_hd__mux2_1
Xhold1133 _25012_/Q vssd1 vssd1 vccd1 vccd1 _17161_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1144 _12797_/X vssd1 vssd1 vccd1 vccd1 _25011_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 _25562_/Q vssd1 vssd1 vccd1 vccd1 _16858_/B sky130_fd_sc_hd__buf_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23823_ _23823_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23824_/A sky130_fd_sc_hd__and2_1
Xhold1166 _13232_/X vssd1 vssd1 vccd1 vccd1 _25091_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1177 _25746_/Q vssd1 vssd1 vccd1 vccd1 _19638_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1188 _12906_/X vssd1 vssd1 vccd1 vccd1 _25032_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1199 _25743_/Q vssd1 vssd1 vccd1 vccd1 _19596_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23754_ _14770_/B _25990_/Q _23754_/S vssd1 vssd1 vccd1 vccd1 _23754_/X sky130_fd_sc_hd__mux2_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20966_ _20969_/A _20969_/C vssd1 vssd1 vccd1 vccd1 _20967_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_166_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22705_ _22705_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22705_/Y sky130_fd_sc_hd__nand2_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23685_ _23685_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23686_/A sky130_fd_sc_hd__and2_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20897_ _20897_/A _21416_/C _20897_/C vssd1 vssd1 vccd1 vccd1 _20898_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_76_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25424_ _25491_/CLK _25424_/D vssd1 vssd1 vccd1 vccd1 _25424_/Q sky130_fd_sc_hd__dfxtp_1
X_22636_ _22627_/Y _22635_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22636_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_166_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25355_ _26308_/CLK hold211/X vssd1 vssd1 vccd1 vccd1 hold209/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22567_ _19844_/A _22566_/A _22566_/Y vssd1 vssd1 vccd1 vccd1 _22569_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24306_ _24306_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24307_/A sky130_fd_sc_hd__and2_1
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21518_ _21518_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21523_/A sky130_fd_sc_hd__nand2_1
X_25286_ _26240_/CLK hold85/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfxtp_1
X_22498_ _22498_/A _22498_/B vssd1 vssd1 vccd1 vccd1 _22499_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_17_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24237_ hold2249/X _26145_/Q _24279_/S vssd1 vssd1 vccd1 vccd1 _24237_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21449_ _21449_/A _21498_/A vssd1 vssd1 vccd1 vccd1 _21451_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24168_ _24168_/A vssd1 vssd1 vccd1 vccd1 _26122_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23119_ _23119_/A _23119_/B vssd1 vssd1 vccd1 vccd1 _23121_/A sky130_fd_sc_hd__nand2_1
X_24099_ _24560_/A vssd1 vssd1 vccd1 vccd1 _24188_/B sky130_fd_sc_hd__buf_8
XFILLER_0_101_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16990_ _20099_/B _25879_/Q _25815_/Q vssd1 vssd1 vccd1 vccd1 _16991_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_101_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15941_ _15941_/A _15941_/B vssd1 vssd1 vccd1 vccd1 _15942_/A sky130_fd_sc_hd__and2_1
X_18660_ _18660_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18660_/Y sky130_fd_sc_hd__nand2_1
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ _15874_/B _15874_/A vssd1 vssd1 vccd1 vccd1 _15875_/A sky130_fd_sc_hd__or2_1
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2390 _26056_/Q vssd1 vssd1 vccd1 vccd1 hold2390/X sky130_fd_sc_hd__dlygate4sd3_1
X_17611_ _17611_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _17611_/Y sky130_fd_sc_hd__nand2_1
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14823_ _14821_/Y _14822_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14823_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18591_ _18612_/A _18591_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18592_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_188_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ _17542_/A _17542_/B vssd1 vssd1 vccd1 vccd1 _17542_/X sky130_fd_sc_hd__xor2_2
X_14754_ _21933_/B _16711_/A vssd1 vssd1 vccd1 vccd1 _14755_/A sky130_fd_sc_hd__nand2_1
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13705_ _13760_/A hold377/X vssd1 vssd1 vccd1 vccd1 hold378/A sky130_fd_sc_hd__nand2_1
X_14685_ _14688_/A hold317/X vssd1 vssd1 vccd1 vccd1 hold318/A sky130_fd_sc_hd__nand2_1
X_17473_ _17473_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17473_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19212_ _19210_/X _19211_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19212_/Y sky130_fd_sc_hd__a21oi_1
X_16424_ _16676_/A _16424_/B vssd1 vssd1 vccd1 vccd1 _16426_/A sky130_fd_sc_hd__nor2_1
X_13636_ _13642_/A hold835/X vssd1 vssd1 vccd1 vccd1 _13636_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19143_ _19972_/B _19234_/A vssd1 vssd1 vccd1 vccd1 _19145_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_54_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16355_ hold950/X vssd1 vssd1 vccd1 vccd1 _16358_/B sky130_fd_sc_hd__inv_2
X_13567_ _13642_/A hold849/X vssd1 vssd1 vccd1 vccd1 _13567_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_109_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15306_ _15306_/A _15306_/B vssd1 vssd1 vccd1 vccd1 _15326_/B sky130_fd_sc_hd__nand2_1
X_12518_ _23245_/A _12533_/A vssd1 vssd1 vccd1 vccd1 _12518_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16286_ _16297_/B _16286_/B vssd1 vssd1 vccd1 vccd1 _16309_/A sky130_fd_sc_hd__nand2_1
X_19074_ _19074_/A _19074_/B vssd1 vssd1 vccd1 vccd1 _19074_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_48_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13498_ _13522_/A hold530/X vssd1 vssd1 vccd1 vccd1 hold531/A sky130_fd_sc_hd__nand2_1
XFILLER_0_124_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18025_ _19244_/A vssd1 vssd1 vccd1 vccd1 _22219_/B sky130_fd_sc_hd__inv_2
XFILLER_0_41_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15237_ _15235_/Y _15236_/Y _15090_/X vssd1 vssd1 vccd1 vccd1 hold886/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_164_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15168_ _15168_/A vssd1 vssd1 vccd1 vccd1 _25438_/D sky130_fd_sc_hd__clkbuf_1
X_14119_ _25814_/Q vssd1 vssd1 vccd1 vccd1 _18490_/B sky130_fd_sc_hd__inv_2
X_15099_ _15100_/B _15100_/A vssd1 vssd1 vccd1 vccd1 _15101_/A sky130_fd_sc_hd__or2_1
XFILLER_0_10_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19976_ _19974_/Y _19975_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _19976_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18927_ _25708_/Q vssd1 vssd1 vccd1 vccd1 _22692_/B sky130_fd_sc_hd__inv_2
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18858_ _18858_/A _18858_/B vssd1 vssd1 vccd1 vccd1 _18858_/X sky130_fd_sc_hd__xor2_1
X_17809_ _18611_/A _17813_/B vssd1 vssd1 vccd1 vccd1 _17811_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18789_ _18951_/A _18793_/B vssd1 vssd1 vccd1 vccd1 _18791_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20820_ _20820_/A _25859_/Q vssd1 vssd1 vccd1 vccd1 _20825_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_82_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20751_ _20751_/A _22590_/B vssd1 vssd1 vccd1 vccd1 _20752_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_65_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23470_ hold191/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23470_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_175_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20682_ _20682_/A _20682_/B vssd1 vssd1 vccd1 vccd1 _21645_/B sky130_fd_sc_hd__nand2_8
XFILLER_0_46_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22421_ _22421_/A vssd1 vssd1 vccd1 vccd1 _22421_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25140_ _25785_/CLK hold511/X vssd1 vssd1 vccd1 vccd1 hold509/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22352_ _22353_/B _22353_/A vssd1 vssd1 vccd1 vccd1 _22354_/A sky130_fd_sc_hd__or2_1
XFILLER_0_116_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21303_ _21662_/B _21710_/B vssd1 vssd1 vccd1 vccd1 _21305_/A sky130_fd_sc_hd__nand2_1
X_25071_ _26284_/CLK _25071_/D vssd1 vssd1 vccd1 vccd1 _25071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22283_ _22283_/A _25855_/Q vssd1 vssd1 vccd1 vccd1 _22284_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_131_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24022_ _24022_/A vssd1 vssd1 vccd1 vccd1 _26075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold230 hold230/A vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
X_21234_ _21234_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21234_/Y sky130_fd_sc_hd__nand2_1
Xhold241 hold241/A vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 hold252/A vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 hold263/A vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 hold274/A vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 hold285/A vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__dlygate4sd3_1
X_21165_ _21165_/A _21165_/B vssd1 vssd1 vccd1 vccd1 _21630_/B sky130_fd_sc_hd__nand2_4
Xhold296 hold296/A vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20116_ _21007_/C vssd1 vssd1 vccd1 vccd1 _21010_/B sky130_fd_sc_hd__inv_2
XFILLER_0_176_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25973_ _26040_/CLK _25973_/D vssd1 vssd1 vccd1 vccd1 _25973_/Q sky130_fd_sc_hd__dfxtp_1
X_21096_ _21096_/A _21096_/B vssd1 vssd1 vccd1 vccd1 _21097_/A sky130_fd_sc_hd__nand2_1
X_24924_ _16501_/B _16508_/Y _24944_/S vssd1 vssd1 vccd1 vccd1 _24924_/X sky130_fd_sc_hd__mux2_1
X_20047_ _20047_/A _22697_/B vssd1 vssd1 vccd1 vccd1 _20051_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_99_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24855_ _24853_/X _24854_/X _24858_/S vssd1 vssd1 vccd1 vccd1 _24855_/X sky130_fd_sc_hd__mux2_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23806_ hold1967/X _26007_/Q _23831_/S vssd1 vssd1 vccd1 vccd1 _23806_/X sky130_fd_sc_hd__mux2_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24786_ _24786_/A vssd1 vssd1 vccd1 vccd1 _26323_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21998_ _21970_/X _21997_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _21998_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23737_ _23737_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23738_/A sky130_fd_sc_hd__and2_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20949_ _20949_/A _20949_/B _20949_/C vssd1 vssd1 vccd1 vccd1 _20953_/A sky130_fd_sc_hd__nand3_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_80_clk clkbuf_leaf_82_clk/A vssd1 vssd1 vccd1 vccd1 _25860_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _14590_/A vssd1 vssd1 vccd1 vccd1 _14525_/A sky130_fd_sc_hd__buf_8
X_23668_ hold2224/X _25962_/Q _23677_/S vssd1 vssd1 vccd1 vccd1 _23668_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13421_ _26333_/Q _19830_/A vssd1 vssd1 vccd1 vccd1 _14666_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_181_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25407_ _26001_/CLK _25407_/D vssd1 vssd1 vccd1 vccd1 _25407_/Q sky130_fd_sc_hd__dfxtp_1
X_22619_ _22620_/B _22620_/A vssd1 vssd1 vccd1 vccd1 _22621_/A sky130_fd_sc_hd__or2_1
XFILLER_0_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23599_ _23599_/A _23599_/B vssd1 vssd1 vccd1 vccd1 _23599_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_181_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16140_ _16150_/B _16140_/B vssd1 vssd1 vccd1 vccd1 _16156_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25338_ _26298_/CLK hold106/X vssd1 vssd1 vccd1 vccd1 hold104/A sky130_fd_sc_hd__dfxtp_1
X_13352_ _13315_/X _13350_/X _13300_/X _13351_/X vssd1 vssd1 vccd1 vccd1 _13352_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16071_ _16071_/A _16071_/B vssd1 vssd1 vccd1 vccd1 _16073_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_180_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25269_ _26096_/CLK hold259/X vssd1 vssd1 vccd1 vccd1 hold257/A sky130_fd_sc_hd__dfxtp_1
X_13283_ _13283_/A vssd1 vssd1 vccd1 vccd1 _19518_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_161_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15022_ _15019_/A _15014_/A _15034_/A vssd1 vssd1 vccd1 vccd1 _15024_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19830_ _19830_/A _20673_/B vssd1 vssd1 vccd1 vccd1 _19830_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_124_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19761_ _19779_/B _19849_/B vssd1 vssd1 vccd1 vccd1 _19763_/A sky130_fd_sc_hd__xnor2_1
X_16973_ _16974_/B _16974_/A vssd1 vssd1 vccd1 vccd1 _16973_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18712_ _18954_/A _25761_/Q vssd1 vssd1 vccd1 vccd1 _18714_/A sky130_fd_sc_hd__nand2_1
X_15924_ _15925_/B _15925_/A vssd1 vssd1 vccd1 vccd1 _15926_/A sky130_fd_sc_hd__or2_1
X_19692_ _19692_/A _19692_/B vssd1 vssd1 vccd1 vccd1 _19692_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_189_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18643_ _19715_/A vssd1 vssd1 vccd1 vccd1 _22348_/B sky130_fd_sc_hd__inv_2
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _15855_/A _15855_/B vssd1 vssd1 vccd1 vccd1 _15856_/B sky130_fd_sc_hd__nand2_1
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806_ _15839_/A _14806_/B vssd1 vssd1 vccd1 vccd1 _22116_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18574_ _18574_/A _20199_/A vssd1 vssd1 vccd1 vccd1 _18919_/A sky130_fd_sc_hd__xor2_4
X_15786_ _15786_/A _15786_/B vssd1 vssd1 vccd1 vccd1 _15823_/A sky130_fd_sc_hd__nor2_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12998_ _12891_/X _14440_/A _12909_/X _25630_/Q vssd1 vssd1 vccd1 vccd1 _12998_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17525_ _17523_/Y _17524_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _17525_/Y sky130_fd_sc_hd__a21oi_1
X_14737_ _25842_/Q _12527_/A _14931_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14737_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_clk _25759_/CLK vssd1 vssd1 vccd1 vccd1 _26084_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17456_ _17456_/A _17456_/B vssd1 vssd1 vccd1 vccd1 _17456_/X sky130_fd_sc_hd__xor2_1
X_14668_ _14666_/Y hold222/X _14646_/X vssd1 vssd1 vccd1 vccd1 hold223/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16407_ _16405_/X _16406_/Y _16231_/A vssd1 vssd1 vccd1 vccd1 _16407_/X sky130_fd_sc_hd__a21o_1
X_13619_ _25734_/Q vssd1 vssd1 vccd1 vccd1 _18138_/B sky130_fd_sc_hd__inv_2
X_17387_ _17385_/Y _17386_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _17387_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14599_ _14599_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14599_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_144_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19126_ _19126_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _19126_/Y sky130_fd_sc_hd__nand2_1
X_16338_ _16490_/A _16380_/B _16337_/X vssd1 vssd1 vccd1 vccd1 _16340_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_27_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19057_ _19186_/A _19057_/B vssd1 vssd1 vccd1 vccd1 _19057_/Y sky130_fd_sc_hd__nand2_1
X_16269_ _16269_/A _16269_/B vssd1 vssd1 vccd1 vccd1 _16269_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18008_ _18535_/A _18008_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _18008_/X sky130_fd_sc_hd__and3_1
XFILLER_0_61_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19959_ _19959_/A _19970_/A vssd1 vssd1 vccd1 vccd1 _19961_/A sky130_fd_sc_hd__xnor2_1
X_22970_ _22961_/Y _22969_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22970_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_184_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21921_ _22676_/A vssd1 vssd1 vccd1 vccd1 _22187_/A sky130_fd_sc_hd__inv_2
XFILLER_0_179_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24640_ _24640_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24641_/A sky130_fd_sc_hd__and2_1
X_21852_ _22626_/A vssd1 vssd1 vccd1 vccd1 _22128_/A sky130_fd_sc_hd__inv_2
XFILLER_0_117_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20803_ _20803_/A _20803_/B _21368_/C vssd1 vssd1 vccd1 vccd1 _20807_/A sky130_fd_sc_hd__nand3_1
X_24571_ _24571_/A vssd1 vssd1 vccd1 vccd1 _26253_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21783_ _25839_/Q _25775_/Q vssd1 vssd1 vccd1 vccd1 _21784_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_148_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_62_clk _25472_/CLK vssd1 vssd1 vccd1 vccd1 _25515_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23522_ hold92/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23522_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_72_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26310_ _26313_/CLK _26310_/D vssd1 vssd1 vccd1 vccd1 _26310_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_136_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20734_ _20733_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20734_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26241_ _26244_/CLK _26241_/D vssd1 vssd1 vccd1 vccd1 _26241_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_46_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23453_ hold170/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23453_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_19_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20665_ _20665_/A _25855_/Q vssd1 vssd1 vccd1 vccd1 _20669_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_151_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22404_ _22389_/X _22403_/Y _17229_/B vssd1 vssd1 vccd1 vccd1 _22404_/Y sky130_fd_sc_hd__o21ai_1
X_26172_ _26175_/CLK _26172_/D vssd1 vssd1 vccd1 vccd1 _26172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23384_ hold155/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23384_/X sky130_fd_sc_hd__or2b_1
X_20596_ _20596_/A _22488_/B vssd1 vssd1 vccd1 vccd1 _20597_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_150_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25123_ _26335_/CLK _25123_/D vssd1 vssd1 vccd1 vccd1 _25123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22335_ _22775_/A _22923_/A vssd1 vssd1 vccd1 vccd1 _22338_/A sky130_fd_sc_hd__nand2_1
X_25054_ _25636_/CLK _25054_/D vssd1 vssd1 vccd1 vccd1 _25054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22266_ _22266_/A _25883_/Q vssd1 vssd1 vccd1 vccd1 _22266_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_143_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24005_ _24560_/A vssd1 vssd1 vccd1 vccd1 _24096_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_0_131_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21217_ _21216_/B _21217_/B _21217_/C vssd1 vssd1 vccd1 vccd1 _21218_/B sky130_fd_sc_hd__nand3b_1
X_22197_ _22198_/A _22198_/C _23122_/A vssd1 vssd1 vccd1 vccd1 _22197_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21148_ _26309_/Q hold695/X vssd1 vssd1 vccd1 vccd1 _21148_/Y sky130_fd_sc_hd__nand2_1
X_25956_ _26021_/CLK _25956_/D vssd1 vssd1 vccd1 vccd1 _25956_/Q sky130_fd_sc_hd__dfxtp_1
X_13970_ _18087_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13970_/Y sky130_fd_sc_hd__nor2_1
X_21079_ _21081_/B _21081_/C vssd1 vssd1 vccd1 vccd1 _21080_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_189_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24907_ _24899_/X _24906_/X _24949_/S vssd1 vssd1 vccd1 vccd1 _24908_/A sky130_fd_sc_hd__mux2_1
X_12921_ _12891_/X _14391_/A _12909_/X _25615_/Q vssd1 vssd1 vccd1 vccd1 _12921_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25887_ _26084_/CLK _25887_/D vssd1 vssd1 vccd1 vccd1 _25887_/Q sky130_fd_sc_hd__dfxtp_2
X_15640_ _16911_/A _15640_/B vssd1 vssd1 vccd1 vccd1 _15641_/B sky130_fd_sc_hd__and2_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24838_ _15123_/A _15144_/B _24860_/S vssd1 vssd1 vccd1 vccd1 _24838_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12852_ _12726_/B _14352_/A _12752_/X _25602_/Q vssd1 vssd1 vccd1 vccd1 _12852_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15571_ _16883_/A _24864_/A vssd1 vssd1 vccd1 vccd1 _15572_/B sky130_fd_sc_hd__nand2_1
X_12783_ _26220_/Q _25589_/Q vssd1 vssd1 vccd1 vccd1 _14310_/A sky130_fd_sc_hd__xor2_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24769_ hold2532/X _26318_/Q _24817_/S vssd1 vssd1 vccd1 vccd1 _24769_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_53_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _26009_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17310_ _17308_/X _17241_/X _17309_/X vssd1 vssd1 vccd1 vccd1 _17311_/A sky130_fd_sc_hd__a21o_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14522_ _14525_/A hold320/X vssd1 vssd1 vccd1 vccd1 hold321/A sky130_fd_sc_hd__nand2_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ _18290_/A _21074_/A vssd1 vssd1 vccd1 vccd1 _18637_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17241_ _22704_/A vssd1 vssd1 vccd1 vccd1 _17241_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_127_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14453_ _14465_/A hold341/X vssd1 vssd1 vccd1 vccd1 hold342/A sky130_fd_sc_hd__nand2_1
XFILLER_0_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13404_ _26202_/Q _13239_/X _13403_/X vssd1 vssd1 vccd1 vccd1 _13404_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_37_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17172_ _17492_/A _17570_/A vssd1 vssd1 vccd1 vccd1 _17173_/B sky130_fd_sc_hd__xnor2_1
X_14384_ _14382_/Y hold165/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold166/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16123_ _16123_/A _16123_/B vssd1 vssd1 vccd1 vccd1 _16124_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_153_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13335_ _13335_/A vssd1 vssd1 vccd1 vccd1 _19630_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16054_ _16056_/A _16054_/B _16054_/C vssd1 vssd1 vccd1 vccd1 _16273_/C sky130_fd_sc_hd__and3_1
X_13266_ _26308_/Q _19473_/A vssd1 vssd1 vccd1 vccd1 _14589_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_110_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15005_ _22144_/B _15778_/B _15006_/B vssd1 vssd1 vccd1 vccd1 _15005_/X sky130_fd_sc_hd__a21o_1
X_13197_ _13049_/X _14554_/A _13067_/X _19317_/A vssd1 vssd1 vccd1 vccd1 _13197_/X
+ sky130_fd_sc_hd__a22o_1
X_19813_ _26262_/Q hold713/X vssd1 vssd1 vccd1 vccd1 _19813_/Y sky130_fd_sc_hd__nand2_1
X_19744_ _19744_/A _20439_/B vssd1 vssd1 vccd1 vccd1 _19744_/Y sky130_fd_sc_hd__nor2_1
X_16956_ _16977_/A _16956_/B vssd1 vssd1 vccd1 vccd1 _16956_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_21_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15907_ _15907_/A _15907_/B vssd1 vssd1 vccd1 vccd1 _15908_/B sky130_fd_sc_hd__nand2_1
X_19675_ _20235_/A _19673_/Y _20240_/C vssd1 vssd1 vccd1 vccd1 _19763_/B sky130_fd_sc_hd__o21a_2
X_16887_ _16885_/Y _16886_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16887_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18626_ _18626_/A _18626_/B vssd1 vssd1 vccd1 vccd1 _22326_/A sky130_fd_sc_hd__nand2_1
X_15838_ hold506/X vssd1 vssd1 vccd1 vccd1 _15844_/B sky130_fd_sc_hd__inv_2
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18557_ _19026_/A _18557_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18557_/X sky130_fd_sc_hd__and3_1
X_15769_ _15787_/A _15786_/B vssd1 vssd1 vccd1 vccd1 _15769_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_188_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_clk _25472_/CLK vssd1 vssd1 vccd1 vccd1 _25573_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17508_ _17506_/X _17241_/X _17507_/X vssd1 vssd1 vccd1 vccd1 _17509_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_74_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18488_ _18954_/A _25750_/Q vssd1 vssd1 vccd1 vccd1 _18490_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_157_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17439_ _17437_/Y _17438_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _17439_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_14 _23496_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 _18718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_36 _26213_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_47 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_58 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20450_ _21547_/A vssd1 vssd1 vccd1 vccd1 _21546_/A sky130_fd_sc_hd__inv_2
XANTENNA_69 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19109_ _19109_/A _21789_/A _19109_/C vssd1 vssd1 vccd1 vccd1 _19109_/X sky130_fd_sc_hd__and3_1
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20381_ _26286_/Q _20078_/X hold536/X vssd1 vssd1 vccd1 vccd1 _20384_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22120_ _25814_/Q _22120_/B vssd1 vssd1 vccd1 vccd1 _22120_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_140_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22051_ _22051_/A _22051_/B vssd1 vssd1 vccd1 vccd1 _22053_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_11_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21002_ _21002_/A _21002_/B _21002_/C vssd1 vssd1 vccd1 vccd1 _21003_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25810_ _25812_/CLK _25810_/D vssd1 vssd1 vccd1 vccd1 _25810_/Q sky130_fd_sc_hd__dfxtp_2
X_22953_ _22944_/Y _22952_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22953_/X sky130_fd_sc_hd__a21o_1
X_25741_ _25745_/CLK hold982/X vssd1 vssd1 vccd1 vccd1 hold981/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21904_ _25798_/Q _21904_/B vssd1 vssd1 vccd1 vccd1 _21904_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_97_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22884_ _22884_/A _23001_/B _22884_/C vssd1 vssd1 vccd1 vccd1 _22884_/X sky130_fd_sc_hd__and3_1
X_25672_ _26302_/CLK _25672_/D vssd1 vssd1 vccd1 vccd1 _25672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21835_ _25796_/Q _21835_/B vssd1 vssd1 vccd1 vccd1 _21835_/Y sky130_fd_sc_hd__nor2_1
X_24623_ _24623_/A vssd1 vssd1 vccd1 vccd1 _26270_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_clk _25184_/CLK vssd1 vssd1 vccd1 vccd1 _26275_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_183_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24554_ _24554_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24555_/A sky130_fd_sc_hd__and2_1
XFILLER_0_78_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21766_ _21766_/A _21766_/B vssd1 vssd1 vccd1 vccd1 _21766_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_148_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20717_ _20720_/A _20720_/C vssd1 vssd1 vccd1 vccd1 _20719_/A sky130_fd_sc_hd__nand2_1
X_23505_ _24944_/S hold227/A _23504_/X vssd1 vssd1 vccd1 vccd1 _23505_/Y sky130_fd_sc_hd__o21ai_1
X_24485_ _24485_/A vssd1 vssd1 vccd1 vccd1 _26225_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21697_ _26339_/Q _19130_/X hold431/X vssd1 vssd1 vccd1 vccd1 _21700_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26224_ _26234_/CLK _26224_/D vssd1 vssd1 vccd1 vccd1 _26224_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_34_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23436_ hold284/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23436_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_68_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20648_ _20648_/A _20648_/B _21305_/B vssd1 vssd1 vccd1 vccd1 _20652_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_123_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26155_ _26284_/CLK _26155_/D vssd1 vssd1 vccd1 vccd1 _26155_/Q sky130_fd_sc_hd__dfxtp_1
X_23367_ _23372_/A _23377_/B _23367_/C vssd1 vssd1 vccd1 vccd1 _23367_/X sky130_fd_sc_hd__and3_1
X_20579_ _20578_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20579_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_150_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ _26284_/Q _25653_/Q vssd1 vssd1 vccd1 vccd1 _14512_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22318_ _22316_/X _22317_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _22318_/Y sky130_fd_sc_hd__a21oi_2
X_25106_ _26325_/CLK _25106_/D vssd1 vssd1 vccd1 vccd1 _25106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26086_ _26112_/CLK _26086_/D vssd1 vssd1 vccd1 vccd1 _26086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23298_ _23298_/A _23298_/B vssd1 vssd1 vccd1 vccd1 _23299_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25037_ _26121_/CLK _25037_/D vssd1 vssd1 vccd1 vccd1 _25037_/Q sky130_fd_sc_hd__dfxtp_1
X_13051_ _13049_/X _14473_/A _12909_/X _25640_/Q vssd1 vssd1 vccd1 vccd1 _13051_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22249_ _18089_/A _25790_/Q _22247_/Y _22248_/Y vssd1 vssd1 vccd1 vccd1 _22250_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16810_ _16810_/A _16810_/B vssd1 vssd1 vccd1 vccd1 _16810_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_100_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17790_ _18100_/A _17794_/A vssd1 vssd1 vccd1 vccd1 _18098_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16741_ _16739_/X _16711_/X _16740_/Y _25866_/Q _14170_/X vssd1 vssd1 vccd1 vccd1
+ _16742_/A sky130_fd_sc_hd__a32o_1
X_25939_ _25939_/CLK hold478/X vssd1 vssd1 vccd1 vccd1 hold476/A sky130_fd_sc_hd__dfxtp_1
X_13953_ _26290_/Q _13801_/X _13793_/X _13952_/Y vssd1 vssd1 vccd1 vccd1 _13954_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12904_ _26115_/Q _12748_/X _12903_/X vssd1 vssd1 vccd1 vccd1 _12904_/X sky130_fd_sc_hd__a21o_1
X_19460_ _21074_/A _19458_/Y _21078_/C vssd1 vssd1 vccd1 vccd1 _19551_/B sky130_fd_sc_hd__o21a_2
X_16672_ _16672_/A _16697_/B vssd1 vssd1 vccd1 vccd1 _16672_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13884_ _26279_/Q _13801_/X _13793_/X _13883_/Y vssd1 vssd1 vccd1 vccd1 _13885_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18411_ _18411_/A _21237_/A vssd1 vssd1 vccd1 vccd1 _18758_/A sky130_fd_sc_hd__xor2_4
X_15623_ hold946/X vssd1 vssd1 vccd1 vccd1 _15625_/A sky130_fd_sc_hd__inv_2
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19391_ _19407_/B _19478_/B vssd1 vssd1 vccd1 vccd1 _19393_/A sky130_fd_sc_hd__xnor2_1
X_12835_ _26230_/Q _25599_/Q vssd1 vssd1 vccd1 vccd1 _14340_/A sky130_fd_sc_hd__xor2_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _25752_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18342_ _25871_/Q _21912_/A vssd1 vssd1 vccd1 vccd1 _18350_/A sky130_fd_sc_hd__or2_2
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _15550_/B _15516_/B _15531_/B vssd1 vssd1 vccd1 vccd1 _15554_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12766_ hold988/X _14264_/A vssd1 vssd1 vccd1 vccd1 _12766_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _14503_/Y hold66/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18273_ _19199_/A vssd1 vssd1 vccd1 vccd1 _18641_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15485_ _15483_/Y _15484_/Y _15464_/X vssd1 vssd1 vccd1 vccd1 hold917/A sky130_fd_sc_hd__a21oi_1
X_12697_ _12699_/A _24836_/B _12697_/C vssd1 vssd1 vccd1 vccd1 _12697_/X sky130_fd_sc_hd__and3_1
XFILLER_0_140_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17224_ _19830_/A _17224_/B vssd1 vssd1 vccd1 vccd1 _17600_/A sky130_fd_sc_hd__xor2_4
X_14436_ _14434_/Y hold303/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold304/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_182_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17155_ _19275_/A _17155_/B vssd1 vssd1 vccd1 vccd1 _17485_/A sky130_fd_sc_hd__xor2_4
X_14367_ _14367_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14367_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold807 hold807/A vssd1 vssd1 vccd1 vccd1 hold807/X sky130_fd_sc_hd__dlygate4sd3_1
X_16106_ _16106_/A vssd1 vssd1 vccd1 vccd1 _16106_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_141_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold818 hold818/A vssd1 vssd1 vccd1 vccd1 hold818/X sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ _13220_/X _14614_/A _13242_/X _19588_/A vssd1 vssd1 vccd1 vccd1 _13318_/X
+ sky130_fd_sc_hd__a22o_1
Xhold829 hold829/A vssd1 vssd1 vccd1 vccd1 hold829/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_17086_ _20468_/B _25850_/Q _25786_/Q vssd1 vssd1 vccd1 vccd1 _17087_/B sky130_fd_sc_hd__mux2_2
X_14298_ _14298_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14298_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_150_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16037_ _16038_/B _16038_/A vssd1 vssd1 vccd1 vccd1 _16039_/A sky130_fd_sc_hd__or2_1
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13249_ _13220_/X _14578_/A _13242_/X _19430_/A vssd1 vssd1 vccd1 vccd1 _13249_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2208 _14960_/Y vssd1 vssd1 vccd1 vccd1 _25419_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2219 _24098_/X vssd1 vssd1 vccd1 vccd1 _24100_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1507 _25895_/Q vssd1 vssd1 vccd1 vccd1 _23101_/B sky130_fd_sc_hd__buf_1
XFILLER_0_23_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17988_ _18528_/A _25724_/Q vssd1 vssd1 vccd1 vccd1 _17990_/A sky130_fd_sc_hd__nand2_1
Xhold1518 _17643_/Y vssd1 vssd1 vccd1 vccd1 _25643_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1529 _25820_/Q vssd1 vssd1 vccd1 vccd1 _21444_/B sky130_fd_sc_hd__dlygate4sd3_1
X_19727_ _19726_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19728_/B
+ sky130_fd_sc_hd__a211o_1
X_16939_ _16939_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16939_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19658_ _19655_/Y _19658_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19658_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_189_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18609_ _18793_/A _25756_/Q _18891_/C vssd1 vssd1 vccd1 vccd1 _18610_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19589_ _20010_/A _22095_/B _25621_/Q vssd1 vssd1 vccd1 vccd1 _20014_/C sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_17_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _25712_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21620_ _21636_/A _21620_/B _21619_/X vssd1 vssd1 vccd1 vccd1 _21621_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_90_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21551_ _26330_/Q _19130_/X hold783/X vssd1 vssd1 vccd1 vccd1 _21554_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_173_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20502_ _20502_/A _20502_/B vssd1 vssd1 vccd1 vccd1 _20503_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_145_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24270_ hold2201/X hold2182/X _24279_/S vssd1 vssd1 vccd1 vccd1 _24271_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_172_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21482_ _21482_/A _21531_/A vssd1 vssd1 vccd1 vccd1 _21483_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_173_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23221_ _23221_/A vssd1 vssd1 vccd1 vccd1 _25908_/D sky130_fd_sc_hd__clkbuf_1
X_20433_ _20435_/B _20435_/C vssd1 vssd1 vccd1 vccd1 _20434_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23152_ _23152_/A _23152_/B vssd1 vssd1 vccd1 vccd1 _23153_/B sky130_fd_sc_hd__nand2_1
X_20364_ _20364_/A _25886_/Q vssd1 vssd1 vccd1 vccd1 _20370_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22103_ _22103_/A _22792_/A vssd1 vssd1 vccd1 vccd1 _22110_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_113_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23083_ _23083_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _23083_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_140_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20295_ _21144_/B _21482_/A vssd1 vssd1 vccd1 vccd1 _20298_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_80_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22034_ _22032_/Y _22033_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _22034_/Y sky130_fd_sc_hd__a21oi_1
Xhold2720 _26274_/Q vssd1 vssd1 vccd1 vccd1 hold2720/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2731 _24757_/X vssd1 vssd1 vccd1 vccd1 _24758_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2742 _26311_/Q vssd1 vssd1 vccd1 vccd1 hold2742/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2753 _25647_/Q vssd1 vssd1 vccd1 vccd1 hold2753/X sky130_fd_sc_hd__dlygate4sd3_1
X_23985_ _23985_/A vssd1 vssd1 vccd1 vccd1 _26063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25724_ _25791_/CLK _25724_/D vssd1 vssd1 vccd1 vccd1 _25724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22936_ _22927_/Y _22935_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22936_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_79_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25655_ _26289_/CLK _25655_/D vssd1 vssd1 vccd1 vccd1 _25655_/Q sky130_fd_sc_hd__dfxtp_2
X_22867_ _22866_/A _22849_/X _22866_/B vssd1 vssd1 vccd1 vccd1 _22868_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12620_ _12620_/A vssd1 vssd1 vccd1 vccd1 _24977_/D sky130_fd_sc_hd__clkbuf_1
X_24606_ hold2615/X _26265_/Q _24664_/S vssd1 vssd1 vccd1 vccd1 _24606_/X sky130_fd_sc_hd__mux2_1
X_21818_ _22601_/A vssd1 vssd1 vccd1 vccd1 _22103_/A sky130_fd_sc_hd__inv_2
XFILLER_0_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22798_ _26060_/Q vssd1 vssd1 vccd1 vccd1 _22799_/A sky130_fd_sc_hd__inv_2
X_25586_ _25587_/CLK _25586_/D vssd1 vssd1 vccd1 vccd1 _25586_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_167_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ _14267_/A _25903_/Q vssd1 vssd1 vccd1 vccd1 _12551_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_176_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24537_ _24537_/A vssd1 vssd1 vccd1 vccd1 _26242_/D sky130_fd_sc_hd__clkbuf_1
X_21749_ _21749_/A _21749_/B vssd1 vssd1 vccd1 vccd1 _21751_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_109_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15270_ _15270_/A _15270_/B vssd1 vssd1 vccd1 vccd1 _15277_/A sky130_fd_sc_hd__nand2_1
X_12482_ _12482_/A vssd1 vssd1 vccd1 vccd1 _14277_/A sky130_fd_sc_hd__inv_2
XFILLER_0_19_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24468_ _24560_/A vssd1 vssd1 vccd1 vccd1 _24557_/B sky130_fd_sc_hd__buf_8
XFILLER_0_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26207_ _26207_/CLK _26207_/D vssd1 vssd1 vccd1 vccd1 _26207_/Q sky130_fd_sc_hd__dfxtp_1
X_14221_ _26333_/Q _13518_/B _14170_/X _14220_/Y vssd1 vssd1 vccd1 vccd1 _14222_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23419_ _23412_/X _23418_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _23419_/X sky130_fd_sc_hd__mux2_1
X_24399_ _24399_/A vssd1 vssd1 vccd1 vccd1 _26197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14152_ _18592_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14152_/Y sky130_fd_sc_hd__nor2_1
X_26138_ _26139_/CLK _26138_/D vssd1 vssd1 vccd1 vccd1 _26138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13103_ _13018_/X _13101_/X _13096_/X _13102_/X vssd1 vssd1 vccd1 vccd1 _13103_/X
+ sky130_fd_sc_hd__o211a_1
X_14083_ _25808_/Q vssd1 vssd1 vccd1 vccd1 _18368_/B sky130_fd_sc_hd__inv_2
X_18960_ _18960_/A _18960_/B vssd1 vssd1 vccd1 vccd1 _18960_/X sky130_fd_sc_hd__xor2_1
X_26069_ _26069_/CLK _26069_/D vssd1 vssd1 vccd1 vccd1 _26069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17911_ _17911_/A _20740_/A vssd1 vssd1 vccd1 vccd1 _18413_/A sky130_fd_sc_hd__xor2_4
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ _26268_/Q _25637_/Q vssd1 vssd1 vccd1 vccd1 _14461_/A sky130_fd_sc_hd__xor2_2
X_18891_ _18952_/A _25770_/Q _18891_/C vssd1 vssd1 vccd1 vccd1 _18892_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_119_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17842_ _18611_/A _17846_/B vssd1 vssd1 vccd1 vccd1 _17844_/A sky130_fd_sc_hd__nand2_1
X_17773_ _17773_/A _17773_/B vssd1 vssd1 vccd1 vccd1 _18118_/B sky130_fd_sc_hd__nand2_4
X_14985_ _14998_/A _14986_/A vssd1 vssd1 vccd1 vccd1 _14985_/X sky130_fd_sc_hd__or2_1
XFILLER_0_135_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19512_ _19723_/A _19512_/B vssd1 vssd1 vccd1 vccd1 _19512_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_92_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16724_ _16980_/A _16729_/B vssd1 vssd1 vccd1 vccd1 _16726_/B sky130_fd_sc_hd__nand2_1
X_13936_ hold687/X _13935_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold688/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19443_ _19440_/Y _19443_/B _19980_/B vssd1 vssd1 vccd1 vccd1 _19443_/X sky130_fd_sc_hd__and3b_1
X_16655_ _16655_/A _16655_/B vssd1 vssd1 vccd1 vccd1 _16669_/A sky130_fd_sc_hd__nor2_1
X_13867_ hold726/X _13866_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold727/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15606_ _15612_/B vssd1 vssd1 vccd1 vccd1 _15609_/B sky130_fd_sc_hd__inv_2
XFILLER_0_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12818_ _26227_/Q _25596_/Q vssd1 vssd1 vccd1 vccd1 _14331_/A sky130_fd_sc_hd__xor2_2
X_19374_ _20908_/A _21904_/B _25606_/Q vssd1 vssd1 vccd1 vccd1 _20913_/C sky130_fd_sc_hd__nand3_1
X_16586_ _16587_/B _16587_/A vssd1 vssd1 vccd1 vccd1 _16588_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ _14345_/A vssd1 vssd1 vccd1 vccd1 _13798_/X sky130_fd_sc_hd__buf_6
X_18325_ _18325_/A _21154_/B _18325_/C vssd1 vssd1 vccd1 vccd1 _21136_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_155_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15537_ _25565_/Q vssd1 vssd1 vccd1 vccd1 _22948_/B sky130_fd_sc_hd__inv_2
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12749_ _26214_/Q _25583_/Q vssd1 vssd1 vccd1 vccd1 _14292_/A sky130_fd_sc_hd__xor2_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18256_ _21048_/B _19444_/A vssd1 vssd1 vccd1 vccd1 _18257_/B sky130_fd_sc_hd__nand2_1
X_15468_ _15466_/A _15442_/B _15459_/A vssd1 vssd1 vccd1 vccd1 _15468_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17207_ _20818_/B _25859_/Q _25795_/Q vssd1 vssd1 vccd1 vccd1 _17208_/B sky130_fd_sc_hd__mux2_2
X_14419_ _14419_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14419_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_181_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18187_ _18529_/A hold891/A _18529_/C vssd1 vssd1 vccd1 vccd1 _18190_/C sky130_fd_sc_hd__nand3_1
X_15399_ _22812_/B _15812_/B vssd1 vssd1 vccd1 vccd1 _15400_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17138_ _17272_/A _17138_/B vssd1 vssd1 vccd1 vccd1 _17138_/Y sky130_fd_sc_hd__nand2_1
Xhold604 hold604/A vssd1 vssd1 vccd1 vccd1 hold604/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold615 hold615/A vssd1 vssd1 vccd1 vccd1 hold615/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 hold626/A vssd1 vssd1 vccd1 vccd1 hold626/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold637 hold637/A vssd1 vssd1 vccd1 vccd1 hold637/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 hold648/A vssd1 vssd1 vccd1 vccd1 hold648/X sky130_fd_sc_hd__dlygate4sd3_1
X_17069_ _25593_/Q vssd1 vssd1 vccd1 vccd1 _20429_/B sky130_fd_sc_hd__inv_2
XFILLER_0_40_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold659 hold659/A vssd1 vssd1 vccd1 vccd1 hold659/X sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_6_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _26135_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20080_ _26278_/Q hold602/X vssd1 vssd1 vccd1 vccd1 _20080_/Y sky130_fd_sc_hd__nand2_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2005 _24243_/X vssd1 vssd1 vccd1 vccd1 _24244_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2016 _26181_/Q vssd1 vssd1 vccd1 vccd1 hold2016/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2027 _25581_/Q vssd1 vssd1 vccd1 vccd1 _12496_/A sky130_fd_sc_hd__buf_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2038 _24320_/X vssd1 vssd1 vccd1 vccd1 _24321_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1304 _25801_/Q vssd1 vssd1 vccd1 vccd1 _21019_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2049 _25979_/Q vssd1 vssd1 vccd1 vccd1 hold2049/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1315 _16821_/Y vssd1 vssd1 vccd1 vccd1 _25556_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1326 _21046_/Y vssd1 vssd1 vccd1 vccd1 _25802_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1337 _25554_/Q vssd1 vssd1 vccd1 vccd1 _16806_/B sky130_fd_sc_hd__clkbuf_2
Xhold1348 _12845_/X vssd1 vssd1 vccd1 vccd1 _25020_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1359 _25094_/Q vssd1 vssd1 vccd1 vccd1 _18597_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23770_ hold2346/X _14824_/B _23831_/S vssd1 vssd1 vccd1 vccd1 _23771_/A sky130_fd_sc_hd__mux2_1
X_20982_ _20982_/A _20982_/B vssd1 vssd1 vccd1 vccd1 _20983_/A sky130_fd_sc_hd__nand2_1
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22721_ _25709_/Q _22720_/A _22720_/Y vssd1 vssd1 vccd1 vccd1 _22723_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_189_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25440_ _25501_/CLK hold928/X vssd1 vssd1 vccd1 vccd1 hold927/A sky130_fd_sc_hd__dfxtp_1
X_22652_ _22652_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _22652_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21603_ _21636_/A _21603_/B _21602_/X vssd1 vssd1 vccd1 vccd1 _21604_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_34_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22583_ _16750_/B _22421_/X _22577_/X _22578_/Y _22582_/X vssd1 vssd1 vccd1 vccd1
+ _22584_/A sky130_fd_sc_hd__a221o_1
X_25371_ _26193_/CLK hold451/X vssd1 vssd1 vccd1 vccd1 hold449/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24322_ _24322_/A vssd1 vssd1 vccd1 vccd1 _26172_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21534_ _21534_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21539_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24253_ _24253_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24254_/A sky130_fd_sc_hd__and2_1
XFILLER_0_69_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21465_ _21465_/A _21514_/A vssd1 vssd1 vccd1 vccd1 _21467_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23204_ _23204_/A vssd1 vssd1 vccd1 vccd1 _25903_/D sky130_fd_sc_hd__inv_2
XFILLER_0_71_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20416_ _21222_/C _21531_/A vssd1 vssd1 vccd1 vccd1 _20417_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24184_ _26127_/Q hold2159/X _24203_/S vssd1 vssd1 vccd1 vccd1 _24184_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21396_ _21573_/A _21396_/B vssd1 vssd1 vccd1 vccd1 _21396_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_102_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23135_ _23135_/A _23135_/B vssd1 vssd1 vccd1 vccd1 _23137_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_114_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20347_ _20660_/A _20347_/B vssd1 vssd1 vccd1 vccd1 _20347_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23066_ _16926_/B _22421_/A _23060_/X _23061_/Y _23065_/X vssd1 vssd1 vccd1 vccd1
+ _23067_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20278_ _20281_/A _20281_/C vssd1 vssd1 vccd1 vccd1 _20280_/A sky130_fd_sc_hd__nand2_1
X_22017_ _22017_/A _22017_/B vssd1 vssd1 vccd1 vccd1 _22017_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_179_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2550 _24983_/Q vssd1 vssd1 vccd1 vccd1 _12656_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2561 _26334_/Q vssd1 vssd1 vccd1 vccd1 hold2561/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2572 _24507_/X vssd1 vssd1 vccd1 vccd1 _24508_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2583 _24563_/X vssd1 vssd1 vccd1 vccd1 _24564_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2594 _26301_/Q vssd1 vssd1 vccd1 vccd1 hold2594/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1860 _26193_/Q vssd1 vssd1 vccd1 vccd1 hold1860/X sky130_fd_sc_hd__dlygate4sd3_1
X_14770_ _15839_/A _14770_/B vssd1 vssd1 vccd1 vccd1 _22002_/A sky130_fd_sc_hd__nand2_1
Xhold1871 _22291_/Y vssd1 vssd1 vccd1 vccd1 _25855_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23968_ hold2357/X _26058_/Q _24001_/S vssd1 vssd1 vccd1 vccd1 _23968_/X sky130_fd_sc_hd__mux2_1
Xhold1882 _25849_/Q vssd1 vssd1 vccd1 vccd1 _22113_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1893 _25852_/Q vssd1 vssd1 vccd1 vccd1 _22201_/B sky130_fd_sc_hd__dlygate4sd3_1
X_25707_ _25708_/CLK _25707_/D vssd1 vssd1 vccd1 vccd1 _25707_/Q sky130_fd_sc_hd__dfxtp_4
X_13721_ _26253_/Q _13612_/X _13605_/X _13720_/Y vssd1 vssd1 vccd1 vccd1 _13722_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22919_ _22910_/Y _22918_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22919_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23899_ _23899_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23900_/A sky130_fd_sc_hd__and2_1
XFILLER_0_168_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16440_ _16439_/X _16440_/B vssd1 vssd1 vccd1 vccd1 _16440_/X sky130_fd_sc_hd__and2b_1
X_13652_ _18263_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13652_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_67_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25638_ _26142_/CLK _25638_/D vssd1 vssd1 vccd1 vccd1 _25638_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_184_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12603_ _12603_/A vssd1 vssd1 vccd1 vccd1 _24973_/D sky130_fd_sc_hd__clkbuf_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _16371_/A hold914/X vssd1 vssd1 vccd1 vccd1 _16372_/B sky130_fd_sc_hd__nand2_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25569_ _26069_/CLK _25569_/D vssd1 vssd1 vccd1 vccd1 _25569_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ _13583_/A _13583_/B vssd1 vssd1 vccd1 vccd1 _13583_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_137_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18110_ _18252_/A _18110_/B vssd1 vssd1 vccd1 vccd1 _18110_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_82_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15322_ _15311_/A _15306_/B _15306_/A vssd1 vssd1 vccd1 vccd1 _15324_/A sky130_fd_sc_hd__a21bo_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _23629_/B _23199_/C _12726_/B _12533_/X hold6/X vssd1 vssd1 vccd1 vccd1 hold7/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19090_ _20023_/B _20023_/A vssd1 vssd1 vccd1 vccd1 _20024_/A sky130_fd_sc_hd__or2_1
XFILLER_0_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18041_ _18041_/A _18041_/B vssd1 vssd1 vccd1 vccd1 _21834_/A sky130_fd_sc_hd__nand2_1
X_15253_ hold2552/X _15252_/Y _15090_/X vssd1 vssd1 vccd1 vccd1 _15253_/Y sky130_fd_sc_hd__a21oi_1
X_14204_ _14264_/A _14204_/B vssd1 vssd1 vccd1 vccd1 _14204_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15184_ _15184_/A _15184_/B vssd1 vssd1 vccd1 vccd1 _15185_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14135_ _26319_/Q _13988_/X _13981_/X _14134_/Y vssd1 vssd1 vccd1 vccd1 _14136_/B
+ sky130_fd_sc_hd__a22o_1
X_19992_ _19991_/Y _21228_/A _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _19994_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14066_ _18308_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14066_/Y sky130_fd_sc_hd__nor2_1
X_18943_ _18943_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18943_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13017_ _12930_/X _13015_/X _13005_/X _13016_/X vssd1 vssd1 vccd1 vccd1 _13017_/X
+ sky130_fd_sc_hd__o211a_1
X_18874_ _18874_/A _18874_/B _18874_/C vssd1 vssd1 vccd1 vccd1 _22617_/A sky130_fd_sc_hd__nand3_2
X_17825_ _25647_/Q vssd1 vssd1 vccd1 vccd1 _21784_/A sky130_fd_sc_hd__inv_2
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17756_ _17874_/B _17874_/A vssd1 vssd1 vccd1 vccd1 _17875_/B sky130_fd_sc_hd__nand2_1
X_14968_ _14982_/B _15033_/A vssd1 vssd1 vccd1 vccd1 _14968_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16707_ _16701_/Y _16706_/Y _16594_/X vssd1 vssd1 vccd1 vccd1 _16707_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13919_ _14000_/A hold389/X vssd1 vssd1 vccd1 vccd1 hold390/A sky130_fd_sc_hd__nand2_1
XFILLER_0_89_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17687_ _17717_/A _17750_/B _17692_/C vssd1 vssd1 vccd1 vccd1 _17690_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_159_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14899_ _14899_/A _14899_/B vssd1 vssd1 vccd1 vccd1 _14899_/Y sky130_fd_sc_hd__nand2_1
X_19426_ _26235_/Q _12537_/B hold641/X vssd1 vssd1 vccd1 vccd1 _19426_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16638_ _16676_/A _16638_/B vssd1 vssd1 vccd1 vccd1 _16640_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19357_ _19356_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19358_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16569_ _16567_/X _16568_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 hold911/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18308_ _18308_/A _18308_/B _18308_/C vssd1 vssd1 vccd1 vccd1 _21846_/A sky130_fd_sc_hd__nand3_2
X_19288_ _19285_/Y _19288_/B _19980_/B vssd1 vssd1 vccd1 vccd1 _19288_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_5_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18239_ _18445_/A _18243_/B vssd1 vssd1 vccd1 vccd1 _18241_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21250_ _21678_/B _21627_/C vssd1 vssd1 vccd1 vccd1 _21252_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold401 hold401/A vssd1 vssd1 vccd1 vccd1 hold401/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 hold412/A vssd1 vssd1 vccd1 vccd1 hold412/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold423 hold423/A vssd1 vssd1 vccd1 vccd1 hold423/X sky130_fd_sc_hd__dlygate4sd3_1
X_20201_ _20204_/A _20204_/C vssd1 vssd1 vccd1 vccd1 _20202_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_130_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold434 hold434/A vssd1 vssd1 vccd1 vccd1 hold434/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 hold445/A vssd1 vssd1 vccd1 vccd1 hold445/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21181_ _21235_/A _21181_/B vssd1 vssd1 vccd1 vccd1 _21181_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold456 hold456/A vssd1 vssd1 vccd1 vccd1 hold456/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold467 hold467/A vssd1 vssd1 vccd1 vccd1 hold467/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold478 hold478/A vssd1 vssd1 vccd1 vccd1 hold478/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20132_ _20132_/A _20132_/B vssd1 vssd1 vccd1 vccd1 _20135_/B sky130_fd_sc_hd__nand2_1
Xhold489 hold489/A vssd1 vssd1 vccd1 vccd1 hold489/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24940_ hold950/A hold914/A _24940_/S vssd1 vssd1 vccd1 vccd1 _24941_/B sky130_fd_sc_hd__mux2_1
X_20063_ _20063_/A _20063_/B vssd1 vssd1 vccd1 vccd1 _21386_/A sky130_fd_sc_hd__nand2_4
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 _25046_/Q vssd1 vssd1 vccd1 vccd1 _17514_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1112 _16716_/Y vssd1 vssd1 vccd1 vccd1 _25541_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1123 _25555_/Q vssd1 vssd1 vccd1 vccd1 _16813_/B sky130_fd_sc_hd__buf_1
X_24871_ _25916_/Q _24871_/B vssd1 vssd1 vccd1 vccd1 _24959_/B sky130_fd_sc_hd__nor2_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1134 _12802_/X vssd1 vssd1 vccd1 vccd1 _25012_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 _25547_/Q vssd1 vssd1 vccd1 vccd1 _16757_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1156 _16859_/Y vssd1 vssd1 vccd1 vccd1 _25562_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23822_ hold2032/X _26012_/Q _23831_/S vssd1 vssd1 vccd1 vccd1 _23822_/X sky130_fd_sc_hd__mux2_1
Xhold1167 _25407_/Q vssd1 vssd1 vccd1 vccd1 _14860_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1178 _19639_/Y vssd1 vssd1 vccd1 vccd1 _25746_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 _25575_/Q vssd1 vssd1 vccd1 vccd1 _16949_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23753_ _23753_/A vssd1 vssd1 vccd1 vccd1 _25989_/D sky130_fd_sc_hd__clkbuf_1
X_20965_ _20965_/A _20965_/B vssd1 vssd1 vccd1 vccd1 _20969_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22704_ _22704_/A vssd1 vssd1 vccd1 vccd1 _23027_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_178_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23684_ hold2085/X hold1974/X _23754_/S vssd1 vssd1 vccd1 vccd1 _23685_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20896_ _21693_/A _21467_/B vssd1 vssd1 vccd1 vccd1 _20897_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_177_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25423_ _25425_/CLK _25423_/D vssd1 vssd1 vccd1 vccd1 _25423_/Q sky130_fd_sc_hd__dfxtp_1
X_22635_ _22635_/A _22900_/B vssd1 vssd1 vccd1 vccd1 _22635_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_64_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22566_ _22566_/A _22566_/B vssd1 vssd1 vccd1 vccd1 _22566_/Y sky130_fd_sc_hd__nand2_1
X_25354_ _26308_/CLK hold94/X vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24305_ hold2058/X hold1920/X _24356_/S vssd1 vssd1 vccd1 vccd1 _24306_/A sky130_fd_sc_hd__mux2_1
X_21517_ _21517_/A _21517_/B vssd1 vssd1 vccd1 vccd1 _21518_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_145_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22497_ _22890_/B _23040_/B vssd1 vssd1 vccd1 vccd1 _22498_/B sky130_fd_sc_hd__nand2_1
X_25285_ _26235_/CLK hold397/X vssd1 vssd1 vccd1 vccd1 hold395/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24236_ _24236_/A vssd1 vssd1 vccd1 vccd1 _26144_/D sky130_fd_sc_hd__clkbuf_1
X_21448_ _21448_/A _21448_/B _21448_/C vssd1 vssd1 vccd1 vccd1 _21452_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_160_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24167_ _24167_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24168_/A sky130_fd_sc_hd__and2_1
XFILLER_0_47_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21379_ _21379_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21379_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_101_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23118_ _23116_/X _23117_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _23118_/Y sky130_fd_sc_hd__a21oi_1
X_24098_ hold2218/X _26100_/Q _24126_/S vssd1 vssd1 vccd1 vccd1 _24098_/X sky130_fd_sc_hd__mux2_1
Xhold990 hold990/A vssd1 vssd1 vccd1 vccd1 hold990/X sky130_fd_sc_hd__dlygate4sd3_1
X_15940_ _15940_/A _15940_/B vssd1 vssd1 vccd1 vccd1 _15941_/A sky130_fd_sc_hd__nor2_1
X_23049_ _23049_/A _23193_/B _23049_/C vssd1 vssd1 vccd1 vccd1 _23049_/X sky130_fd_sc_hd__and3_1
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15871_ _16274_/A _15895_/B _15870_/Y vssd1 vssd1 vccd1 vccd1 _15874_/A sky130_fd_sc_hd__a21o_1
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2380 _26235_/Q vssd1 vssd1 vccd1 vccd1 hold2380/X sky130_fd_sc_hd__dlygate4sd3_1
X_17610_ _17608_/X _17528_/X _17609_/X vssd1 vssd1 vccd1 vccd1 _17611_/A sky130_fd_sc_hd__a21o_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14822_ _14900_/A _14822_/B vssd1 vssd1 vccd1 vccd1 _14822_/Y sky130_fd_sc_hd__nand2_1
Xhold2391 _26134_/Q vssd1 vssd1 vccd1 vccd1 hold2391/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ _18611_/A _25755_/Q vssd1 vssd1 vccd1 vccd1 _18592_/A sky130_fd_sc_hd__nand2_1
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1690 _25874_/Q vssd1 vssd1 vccd1 vccd1 _22756_/B sky130_fd_sc_hd__buf_1
X_17541_ _17541_/A _17593_/A vssd1 vssd1 vccd1 vccd1 _17542_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _14759_/B _21934_/A vssd1 vssd1 vccd1 vccd1 _21933_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_169_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13704_ hold573/X _13703_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold574/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17472_ _17470_/X _17241_/X _17471_/X vssd1 vssd1 vccd1 vccd1 _17473_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14684_ _14684_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _14684_/Y sky130_fd_sc_hd__nand2_1
X_19211_ _19211_/A _19211_/B vssd1 vssd1 vccd1 vccd1 _19211_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_67_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16423_ _16421_/Y _16422_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 hold895/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_168_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ _13630_/Y _13634_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold842/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19142_ _20309_/A _18151_/B _20314_/C vssd1 vssd1 vccd1 vccd1 _19234_/A sky130_fd_sc_hd__o21ai_4
X_16354_ _16352_/X _16353_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 hold969/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13566_ hold561/X _13565_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold562/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15305_ _15305_/A _15305_/B vssd1 vssd1 vccd1 vccd1 _15306_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12517_ _24050_/A input2/X vssd1 vssd1 vccd1 vccd1 _12533_/A sky130_fd_sc_hd__and2b_2
XFILLER_0_124_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19073_ _19073_/A _19073_/B vssd1 vssd1 vccd1 vccd1 _19074_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16285_ _16285_/A _16285_/B vssd1 vssd1 vccd1 vccd1 _16286_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_180_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13497_ _13492_/Y _13496_/Y _12558_/B vssd1 vssd1 vccd1 vccd1 hold767/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18024_ _18024_/A _19177_/A vssd1 vssd1 vccd1 vccd1 _19053_/A sky130_fd_sc_hd__xnor2_4
X_15236_ _15956_/A hold885/X vssd1 vssd1 vccd1 vccd1 _15236_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_152_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15167_ _15167_/A _23629_/B vssd1 vssd1 vccd1 vccd1 _15168_/A sky130_fd_sc_hd__and2_1
XFILLER_0_125_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14118_ _14118_/A hold821/X vssd1 vssd1 vccd1 vccd1 _14118_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15098_ _16146_/B _15543_/B vssd1 vssd1 vccd1 vccd1 _15100_/A sky130_fd_sc_hd__nand2b_1
X_19975_ _19975_/A _19975_/B vssd1 vssd1 vccd1 vccd1 _19975_/Y sky130_fd_sc_hd__nand2_1
X_18926_ _25708_/Q _20044_/B vssd1 vssd1 vccd1 vccd1 _18929_/A sky130_fd_sc_hd__nor2_1
X_14049_ _14061_/A _14049_/B vssd1 vssd1 vccd1 vccd1 _14049_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_157_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18857_ _18996_/A _19045_/A vssd1 vssd1 vccd1 vccd1 _18858_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17808_ _25855_/Q _22277_/A vssd1 vssd1 vccd1 vccd1 _17816_/A sky130_fd_sc_hd__or2_2
X_18788_ _25893_/Q _22512_/A vssd1 vssd1 vccd1 vccd1 _18796_/A sky130_fd_sc_hd__or2_2
XFILLER_0_171_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17739_ _17709_/A _17709_/C _17738_/Y vssd1 vssd1 vccd1 vccd1 _17740_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20750_ _21403_/B vssd1 vssd1 vccd1 vccd1 _21400_/C sky130_fd_sc_hd__inv_2
XFILLER_0_175_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19409_ _19401_/X _19408_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19409_/Y sky130_fd_sc_hd__o21ai_1
X_20681_ _20681_/A _20681_/B _20681_/C vssd1 vssd1 vccd1 vccd1 _20682_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_119_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22420_ _22420_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _22420_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22351_ _19715_/A _22350_/A _22350_/Y vssd1 vssd1 vccd1 vccd1 _22353_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21302_ _21302_/A _21302_/B _21302_/C vssd1 vssd1 vccd1 vccd1 _21306_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_116_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25070_ _26154_/CLK _25070_/D vssd1 vssd1 vccd1 vccd1 _25070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22282_ _25855_/Q _22283_/A vssd1 vssd1 vccd1 vccd1 _22284_/A sky130_fd_sc_hd__or2_1
XFILLER_0_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24021_ _24021_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24022_/A sky130_fd_sc_hd__and2_1
XFILLER_0_14_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold220 hold220/A vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
X_21233_ _21233_/A _21233_/B vssd1 vssd1 vccd1 vccd1 _21234_/A sky130_fd_sc_hd__nand2_1
Xhold231 hold231/A vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 hold242/A vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 hold253/A vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 hold264/A vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21164_ _21164_/A _21164_/B _21164_/C vssd1 vssd1 vccd1 vccd1 _21165_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_106_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold275 hold275/A vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 hold286/A vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 hold297/A vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__dlygate4sd3_1
X_20115_ _20115_/A _20115_/B vssd1 vssd1 vccd1 vccd1 _21007_/C sky130_fd_sc_hd__xor2_4
X_25972_ _26040_/CLK _25972_/D vssd1 vssd1 vccd1 vccd1 _25972_/Q sky130_fd_sc_hd__dfxtp_1
X_21095_ _21636_/A _21095_/B _21094_/X vssd1 vssd1 vccd1 vccd1 _21096_/B sky130_fd_sc_hd__or3b_1
X_24923_ _24957_/S _24923_/B vssd1 vssd1 vccd1 vccd1 _24923_/Y sky130_fd_sc_hd__nor2_1
X_20046_ _25900_/Q vssd1 vssd1 vccd1 vccd1 _22697_/B sky130_fd_sc_hd__inv_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24854_ _15441_/A _15458_/B _24860_/S vssd1 vssd1 vccd1 vccd1 _24854_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23805_ _23805_/A vssd1 vssd1 vccd1 vccd1 _26006_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24785_ _24785_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24786_/A sky130_fd_sc_hd__and2_1
X_21997_ _21995_/X _21996_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _21997_/Y sky130_fd_sc_hd__a21oi_2
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23736_ _14714_/B _25984_/Q _23754_/S vssd1 vssd1 vccd1 vccd1 _23736_/X sky130_fd_sc_hd__mux2_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20948_ _21500_/B _21451_/B vssd1 vssd1 vccd1 vccd1 _20949_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_166_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23667_ _23667_/A vssd1 vssd1 vccd1 vccd1 _25961_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20879_ _20879_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _20879_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_181_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25406_ _25999_/CLK _25406_/D vssd1 vssd1 vccd1 vccd1 _25406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13420_ _13420_/A vssd1 vssd1 vccd1 vccd1 _19830_/A sky130_fd_sc_hd__buf_6
XFILLER_0_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22618_ _25705_/Q _22617_/A _22617_/Y vssd1 vssd1 vccd1 vccd1 _22620_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23598_ _23598_/A _23598_/B vssd1 vssd1 vccd1 vccd1 _23599_/A sky130_fd_sc_hd__or2_1
XFILLER_0_64_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25337_ _26171_/CLK hold229/X vssd1 vssd1 vccd1 vccd1 hold227/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13351_ _18920_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13351_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22549_ _22549_/A _22549_/B vssd1 vssd1 vccd1 vccd1 _22550_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16070_ _16070_/A _16070_/B vssd1 vssd1 vccd1 vccd1 _16084_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_23_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25268_ _26221_/CLK hold142/X vssd1 vssd1 vccd1 vccd1 hold140/A sky130_fd_sc_hd__dfxtp_1
X_13282_ _13207_/X _13280_/X _13192_/X _13281_/X vssd1 vssd1 vccd1 vccd1 _13282_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15021_ _15021_/A _15021_/B vssd1 vssd1 vccd1 vccd1 _15034_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_60_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24219_ hold2234/X hold1961/X _24279_/S vssd1 vssd1 vccd1 vccd1 _24220_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_121_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25199_ _26281_/CLK hold613/X vssd1 vssd1 vccd1 vccd1 hold611/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16972_ _22145_/B _16977_/B vssd1 vssd1 vccd1 vccd1 _16974_/B sky130_fd_sc_hd__nand2_1
X_19760_ _20478_/A _19758_/Y _20483_/C vssd1 vssd1 vccd1 vccd1 _19849_/B sky130_fd_sc_hd__o21a_1
X_15923_ _15900_/A _15941_/B _15922_/Y vssd1 vssd1 vccd1 vccd1 _15925_/A sky130_fd_sc_hd__a21o_1
X_18711_ _18711_/A _25825_/Q _18711_/C vssd1 vssd1 vccd1 vccd1 _20487_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19691_ _19692_/B _19692_/A vssd1 vssd1 vccd1 vccd1 _19691_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_212_clk _26093_/CLK vssd1 vssd1 vccd1 vccd1 _26219_/CLK sky130_fd_sc_hd__clkbuf_16
X_18642_ _18640_/Y _18641_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25676_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_189_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _15855_/B _15855_/A vssd1 vssd1 vccd1 vccd1 _15856_/A sky130_fd_sc_hd__or2_1
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14805_ _14803_/Y _14804_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14805_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ _20208_/B _22239_/A vssd1 vssd1 vccd1 vccd1 _20199_/A sky130_fd_sc_hd__nand2_2
X_15785_ _15783_/X hold1383/X _15464_/X vssd1 vssd1 vccd1 vccd1 _15785_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12997_ _26261_/Q _25630_/Q vssd1 vssd1 vccd1 vccd1 _14440_/A sky130_fd_sc_hd__xor2_2
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17524_ _17605_/A _17524_/B vssd1 vssd1 vccd1 vccd1 _17524_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_87_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14736_ _14736_/A vssd1 vssd1 vccd1 vccd1 _14931_/A sky130_fd_sc_hd__inv_2
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17455_ _17505_/A _17622_/B vssd1 vssd1 vccd1 vccd1 _17456_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14667_ _14688_/A hold221/X vssd1 vssd1 vccd1 vccd1 hold222/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16406_ _16406_/A _16416_/A vssd1 vssd1 vccd1 vccd1 _16406_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_131_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13618_ _13642_/A hold491/X vssd1 vssd1 vccd1 vccd1 hold492/A sky130_fd_sc_hd__nand2_1
XFILLER_0_172_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17386_ _17467_/A _17386_/B vssd1 vssd1 vccd1 vccd1 _17386_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_55_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14598_ _14596_/Y hold159/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold160/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19125_ _19120_/X _18879_/X _19124_/X vssd1 vssd1 vccd1 vccd1 _19126_/A sky130_fd_sc_hd__a21o_1
X_16337_ _16310_/X _16334_/B _16319_/A _16336_/Y vssd1 vssd1 vccd1 vccd1 _16337_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13549_ _25723_/Q vssd1 vssd1 vccd1 vccd1 _17944_/B sky130_fd_sc_hd__inv_2
XFILLER_0_55_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19056_ _19056_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _19056_/Y sky130_fd_sc_hd__nand2_1
X_16268_ _16266_/Y _16267_/Y _16076_/X vssd1 vssd1 vccd1 vccd1 _16268_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18007_ _18997_/A _18007_/B vssd1 vssd1 vccd1 vccd1 _18007_/X sky130_fd_sc_hd__xor2_4
X_15219_ hold2650/X _15218_/Y _15090_/X vssd1 vssd1 vccd1 vccd1 _15219_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16199_ _16208_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16199_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_112_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19958_ _19958_/A _19980_/B _19958_/C vssd1 vssd1 vccd1 vccd1 _19958_/X sky130_fd_sc_hd__and3_1
X_18909_ _25899_/Q _22664_/A vssd1 vssd1 vccd1 vccd1 _18917_/A sky130_fd_sc_hd__or2_2
X_19889_ _19887_/X _19888_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19889_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_203_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _26109_/CLK sky130_fd_sc_hd__clkbuf_16
X_21920_ _23135_/A _22676_/A vssd1 vssd1 vccd1 vccd1 _21928_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21851_ _23103_/A _22626_/A vssd1 vssd1 vccd1 vccd1 _21859_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20802_ _21692_/B _21419_/B vssd1 vssd1 vccd1 vccd1 _20803_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_148_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21782_ _22073_/A _23072_/A vssd1 vssd1 vccd1 vccd1 _21788_/B sky130_fd_sc_hd__nand2_1
X_24570_ _24570_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24571_/A sky130_fd_sc_hd__and2_1
XFILLER_0_38_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23521_ _24944_/S hold209/A _23520_/X vssd1 vssd1 vccd1 vccd1 _23521_/Y sky130_fd_sc_hd__o21ai_1
X_20733_ _26295_/Q hold718/X vssd1 vssd1 vccd1 vccd1 _20733_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_92_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26240_ _26240_/CLK _26240_/D vssd1 vssd1 vccd1 vccd1 _26240_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_175_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20664_ _20666_/B _20666_/C vssd1 vssd1 vccd1 vccd1 _20665_/A sky130_fd_sc_hd__nand2_1
X_23452_ _24922_/S hold302/A _23451_/X vssd1 vssd1 vccd1 vccd1 _23452_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_163_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22403_ _22401_/X _22402_/Y _22900_/B vssd1 vssd1 vccd1 vccd1 _22403_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23383_ _23391_/A vssd1 vssd1 vccd1 vccd1 _24942_/S sky130_fd_sc_hd__buf_12
X_26171_ _26171_/CLK _26171_/D vssd1 vssd1 vccd1 vccd1 _26171_/Q sky130_fd_sc_hd__dfxtp_1
X_20595_ _21335_/C vssd1 vssd1 vccd1 vccd1 _21338_/B sky130_fd_sc_hd__inv_2
XFILLER_0_34_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25122_ _26335_/CLK _25122_/D vssd1 vssd1 vccd1 vccd1 _25122_/Q sky130_fd_sc_hd__dfxtp_1
X_22334_ _22924_/A vssd1 vssd1 vccd1 vccd1 _22923_/A sky130_fd_sc_hd__inv_2
XFILLER_0_147_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22265_ _22265_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _22265_/X sky130_fd_sc_hd__and2_1
XFILLER_0_131_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25053_ _26139_/CLK _25053_/D vssd1 vssd1 vccd1 vccd1 _25053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24004_ hold2449/X hold2430/X _24047_/S vssd1 vssd1 vccd1 vccd1 _24006_/A sky130_fd_sc_hd__mux2_1
X_21216_ _21216_/A _21216_/B vssd1 vssd1 vccd1 vccd1 _21218_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22196_ _22196_/A _22196_/B vssd1 vssd1 vccd1 vccd1 _23122_/A sky130_fd_sc_hd__nand2_8
X_21147_ _26309_/Q _20731_/X hold695/X vssd1 vssd1 vccd1 vccd1 _21150_/B sky130_fd_sc_hd__a21oi_1
X_25955_ _26021_/CLK _25955_/D vssd1 vssd1 vccd1 vccd1 _25955_/Q sky130_fd_sc_hd__dfxtp_1
X_21078_ _25868_/Q _21078_/B _21078_/C vssd1 vssd1 vccd1 vccd1 _21081_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_77_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24906_ _24902_/X _24905_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _24906_/X sky130_fd_sc_hd__mux2_1
X_12920_ _26246_/Q _25615_/Q vssd1 vssd1 vccd1 vccd1 _14391_/A sky130_fd_sc_hd__xor2_1
X_20029_ _21676_/A _21369_/A vssd1 vssd1 vccd1 vccd1 _20031_/A sky130_fd_sc_hd__nand2_1
X_25886_ _26080_/CLK _25886_/D vssd1 vssd1 vccd1 vccd1 _25886_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24837_ _24837_/A vssd1 vssd1 vccd1 vccd1 _26340_/D sky130_fd_sc_hd__clkbuf_1
X_12851_ _26233_/Q _25602_/Q vssd1 vssd1 vccd1 vccd1 _14352_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_68_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15570_ _24864_/A _16883_/A vssd1 vssd1 vccd1 vccd1 _15572_/A sky130_fd_sc_hd__or2_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12782_ _12746_/X _12780_/X _14910_/B _12781_/X vssd1 vssd1 vccd1 vccd1 _12782_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24768_ _24768_/A vssd1 vssd1 vccd1 vccd1 _26317_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14521_ _14521_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14521_/Y sky130_fd_sc_hd__nand2_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23719_ _23719_/A vssd1 vssd1 vccd1 vccd1 _25978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24699_ _24699_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24700_/A sky130_fd_sc_hd__and2_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17240_ _21716_/A vssd1 vssd1 vccd1 vccd1 _22704_/A sky130_fd_sc_hd__buf_8
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _14452_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14452_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13403_ _13220_/X _14657_/A _13242_/X _19788_/A vssd1 vssd1 vccd1 vccd1 _13403_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17171_ _19774_/A _17171_/B vssd1 vssd1 vccd1 vccd1 _17570_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_24_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14383_ _14404_/A hold164/X vssd1 vssd1 vccd1 vccd1 hold165/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16122_ _16123_/B _16123_/A vssd1 vssd1 vccd1 vccd1 _16124_/A sky130_fd_sc_hd__or2_1
XFILLER_0_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13334_ _13315_/X _13332_/X _13300_/X _13333_/X vssd1 vssd1 vccd1 vccd1 _13334_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16053_ _16053_/A _16053_/B vssd1 vssd1 vccd1 vccd1 _16056_/A sky130_fd_sc_hd__and2_1
XFILLER_0_150_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13265_ _13265_/A vssd1 vssd1 vccd1 vccd1 _19473_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_150_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15004_ _15002_/X hold2297/X _14928_/X vssd1 vssd1 vccd1 vccd1 _15004_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13196_ _26297_/Q _19317_/A vssd1 vssd1 vccd1 vccd1 _14554_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_138_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19812_ _26262_/Q _19134_/X hold713/X vssd1 vssd1 vccd1 vccd1 _19812_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19743_ _19740_/Y _19743_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19743_/X sky130_fd_sc_hd__and3b_1
X_16955_ _16955_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16955_/Y sky130_fd_sc_hd__nand2_1
X_15906_ _15907_/B _15907_/A vssd1 vssd1 vccd1 vccd1 _15908_/A sky130_fd_sc_hd__or2_1
X_16886_ _16977_/A _16886_/B vssd1 vssd1 vccd1 vccd1 _16886_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19674_ _20235_/A _22267_/B _25627_/Q vssd1 vssd1 vccd1 vccd1 _20240_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_95_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15837_ _16274_/A vssd1 vssd1 vccd1 vccd1 _15846_/B sky130_fd_sc_hd__inv_2
X_18625_ _20322_/B _19701_/A vssd1 vssd1 vccd1 vccd1 _18626_/B sky130_fd_sc_hd__nand2_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15768_ _15786_/B _15787_/A vssd1 vssd1 vccd1 vccd1 _15768_/X sky130_fd_sc_hd__or2_1
X_18556_ _19082_/A vssd1 vssd1 vccd1 vccd1 _19026_/A sky130_fd_sc_hd__clkbuf_8
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14719_ _25840_/Q _13466_/A _14718_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14720_/A
+ sky130_fd_sc_hd__a22o_1
X_17507_ _17624_/A _17507_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17507_/X sky130_fd_sc_hd__and3_1
XFILLER_0_129_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18487_ _18487_/A _25814_/Q _18487_/C vssd1 vssd1 vccd1 vccd1 _20062_/C sky130_fd_sc_hd__nand3_2
X_15699_ _15560_/A _15825_/A _15829_/A vssd1 vssd1 vccd1 vccd1 _15701_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_118_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17438_ _17467_/A _17438_/B vssd1 vssd1 vccd1 vccd1 _17438_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_15 _23602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_26 _18878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_37 _25912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_48 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17369_ _21184_/B _25872_/Q _25808_/Q vssd1 vssd1 vccd1 vccd1 _17370_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_103_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_59 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19108_ _26213_/Q _19483_/A hold452/X vssd1 vssd1 vccd1 vccd1 _19109_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_103_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20380_ _20380_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20385_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19039_ _19039_/A _19039_/B vssd1 vssd1 vccd1 vccd1 _19039_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_141_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22050_ _25847_/Q _25783_/Q vssd1 vssd1 vccd1 vccd1 _22051_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21001_ _21001_/A _21001_/B vssd1 vssd1 vccd1 vccd1 _21003_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25740_ _25740_/CLK _25740_/D vssd1 vssd1 vccd1 vccd1 _25740_/Q sky130_fd_sc_hd__dfxtp_1
X_22952_ _22952_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _22952_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21903_ _21903_/A _25862_/Q vssd1 vssd1 vccd1 vccd1 _21903_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25671_ _26302_/CLK _25671_/D vssd1 vssd1 vccd1 vccd1 _25671_/Q sky130_fd_sc_hd__dfxtp_1
X_22883_ _22882_/A _22849_/X _22882_/B vssd1 vssd1 vccd1 vccd1 _22884_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24622_ _24622_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24623_/A sky130_fd_sc_hd__and2_1
X_21834_ _21834_/A _25860_/Q vssd1 vssd1 vccd1 vccd1 _21834_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_38_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24553_ hold2689/X hold2688/X _24587_/S vssd1 vssd1 vccd1 vccd1 _24554_/A sky130_fd_sc_hd__mux2_1
X_21765_ _17960_/A _25794_/Q _21763_/Y _21764_/Y vssd1 vssd1 vccd1 vccd1 _21766_/B
+ sky130_fd_sc_hd__a31o_1
X_23504_ hold104/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23504_/X sky130_fd_sc_hd__or2b_1
X_20716_ _20716_/A _22569_/B _20716_/C vssd1 vssd1 vccd1 vccd1 _20720_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_108_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24484_ _24484_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24485_/A sky130_fd_sc_hd__and2_1
X_21696_ _21696_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _21701_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_110_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26223_ _26232_/CLK _26223_/D vssd1 vssd1 vccd1 vccd1 _26223_/Q sky130_fd_sc_hd__dfxtp_2
X_23435_ _24945_/S vssd1 vssd1 vccd1 vccd1 _24922_/S sky130_fd_sc_hd__buf_12
XFILLER_0_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20647_ _21628_/B _21351_/C vssd1 vssd1 vccd1 vccd1 _20648_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_34_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26154_ _26154_/CLK _26154_/D vssd1 vssd1 vccd1 vccd1 _26154_/Q sky130_fd_sc_hd__dfxtp_1
X_23366_ _23366_/A _23366_/B vssd1 vssd1 vccd1 vccd1 _23366_/Y sky130_fd_sc_hd__nand2_1
X_20578_ _26291_/Q hold777/X vssd1 vssd1 vccd1 vccd1 _20578_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25105_ _26190_/CLK _25105_/D vssd1 vssd1 vccd1 vccd1 _25105_/Q sky130_fd_sc_hd__dfxtp_1
X_22317_ _22317_/A _22317_/B _23186_/A vssd1 vssd1 vccd1 vccd1 _22317_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_81_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26085_ _26249_/CLK _26085_/D vssd1 vssd1 vccd1 vccd1 _26085_/Q sky130_fd_sc_hd__dfxtp_1
X_23297_ _23303_/A vssd1 vssd1 vccd1 vccd1 _23301_/A sky130_fd_sc_hd__inv_2
XFILLER_0_131_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25036_ _26119_/CLK _25036_/D vssd1 vssd1 vccd1 vccd1 _25036_/Q sky130_fd_sc_hd__dfxtp_1
X_13050_ _26271_/Q _25640_/Q vssd1 vssd1 vccd1 vccd1 _14473_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_131_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22248_ _25790_/Q _22248_/B vssd1 vssd1 vccd1 vccd1 _22248_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_178_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22179_ _25816_/Q _22179_/B vssd1 vssd1 vccd1 vccd1 _22179_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_121_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16740_ _16740_/A _16740_/B vssd1 vssd1 vccd1 vccd1 _16740_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25938_ _25938_/CLK _25938_/D vssd1 vssd1 vccd1 vccd1 _25938_/Q sky130_fd_sc_hd__dfxtp_1
X_13952_ _17945_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13952_/Y sky130_fd_sc_hd__nor2_1
X_12903_ _12891_/X _14382_/A _12752_/X _25612_/Q vssd1 vssd1 vccd1 vccd1 _12903_/X
+ sky130_fd_sc_hd__a22o_1
X_16671_ _16680_/A _16671_/B vssd1 vssd1 vccd1 vccd1 _16672_/A sky130_fd_sc_hd__xnor2_1
X_25869_ _25876_/CLK _25869_/D vssd1 vssd1 vccd1 vccd1 _25869_/Q sky130_fd_sc_hd__dfxtp_2
X_13883_ _17881_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13883_/Y sky130_fd_sc_hd__nor2_1
X_15622_ hold946/X _15624_/A vssd1 vssd1 vccd1 vccd1 _15626_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_159_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18410_ _21243_/B _22017_/A vssd1 vssd1 vccd1 vccd1 _21237_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_159_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12834_ _12746_/X _12832_/X _12827_/X _12833_/X vssd1 vssd1 vccd1 vccd1 _12834_/X
+ sky130_fd_sc_hd__o211a_1
X_19390_ _20935_/A _19388_/Y _20940_/C vssd1 vssd1 vccd1 vccd1 _19478_/B sky130_fd_sc_hd__o21a_2
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18341_ _18341_/A _18341_/B vssd1 vssd1 vccd1 vccd1 _21912_/A sky130_fd_sc_hd__nand2_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _15553_/A _15822_/A vssd1 vssd1 vccd1 vccd1 _15557_/A sky130_fd_sc_hd__nand2_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12765_ _26088_/Q _12748_/X _12764_/X vssd1 vssd1 vccd1 vccd1 _12765_/X sky130_fd_sc_hd__a21o_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _14525_/A hold65/X vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__nand2_1
XFILLER_0_139_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18272_ _18272_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18272_/Y sky130_fd_sc_hd__nand2_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _15956_/A hold916/X vssd1 vssd1 vccd1 vccd1 _15484_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12696_/A _12713_/A vssd1 vssd1 vccd1 vccd1 _12696_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17223_ _20673_/B _25894_/Q _25830_/Q vssd1 vssd1 vccd1 vccd1 _17224_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14435_ _14465_/A hold302/X vssd1 vssd1 vccd1 vccd1 hold303/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17154_ _20663_/B _25855_/Q _20699_/B vssd1 vssd1 vccd1 vccd1 _17155_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14366_ _14364_/Y hold396/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold397/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16105_ _16160_/A _16158_/B vssd1 vssd1 vccd1 vccd1 _16133_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13317_ _26316_/Q _19588_/A vssd1 vssd1 vccd1 vccd1 _14614_/A sky130_fd_sc_hd__xor2_1
Xhold808 hold808/A vssd1 vssd1 vccd1 vccd1 hold808/X sky130_fd_sc_hd__dlygate4sd3_1
X_17085_ _25594_/Q vssd1 vssd1 vccd1 vccd1 _20468_/B sky130_fd_sc_hd__inv_2
Xhold819 hold819/A vssd1 vssd1 vccd1 vccd1 hold819/X sky130_fd_sc_hd__dlygate4sd3_1
X_14297_ _14295_/Y hold102/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold103/A sky130_fd_sc_hd__a21oi_1
X_16036_ _22203_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _16038_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13248_ _26305_/Q _19430_/A vssd1 vssd1 vccd1 vccd1 _14578_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_149_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13179_ _26166_/Q _13065_/X _13178_/X vssd1 vssd1 vccd1 vccd1 _13179_/X sky130_fd_sc_hd__a21o_1
Xhold2209 _26169_/Q vssd1 vssd1 vccd1 vccd1 hold2209/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1508 _23102_/Y vssd1 vssd1 vccd1 vccd1 _25895_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17987_ _17987_/A _25788_/Q _17987_/C vssd1 vssd1 vccd1 vccd1 _20553_/B sky130_fd_sc_hd__nand3_1
Xhold1519 _25759_/Q vssd1 vssd1 vccd1 vccd1 _19824_/B sky130_fd_sc_hd__dlygate4sd3_1
X_19726_ _26256_/Q hold365/X vssd1 vssd1 vccd1 vccd1 _19726_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_165_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16938_ _16936_/X _16711_/X _16937_/Y _25895_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16939_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19657_ _19656_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19658_/B
+ sky130_fd_sc_hd__a211o_1
X_16869_ _16869_/A _16869_/B vssd1 vssd1 vccd1 vccd1 _16869_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18608_ _18792_/A _18612_/B vssd1 vssd1 vccd1 vccd1 _18610_/A sky130_fd_sc_hd__nand2_1
X_19588_ _19588_/A _20011_/B vssd1 vssd1 vccd1 vccd1 _19588_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18539_ _21099_/A vssd1 vssd1 vccd1 vccd1 _18539_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21550_ _21550_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21555_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20501_ _21042_/A _20501_/B _20500_/X vssd1 vssd1 vccd1 vccd1 _20502_/B sky130_fd_sc_hd__or3b_1
X_21481_ _21481_/A _21530_/A vssd1 vssd1 vccd1 vccd1 _21483_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23220_ _23220_/A _24836_/B _23227_/A vssd1 vssd1 vccd1 vccd1 _23221_/A sky130_fd_sc_hd__and3_1
XFILLER_0_160_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20432_ _25849_/Q _20432_/B _20432_/C vssd1 vssd1 vccd1 vccd1 _20435_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_67_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23151_ _23151_/A _23151_/B vssd1 vssd1 vccd1 vccd1 _23153_/A sky130_fd_sc_hd__nand2_1
X_20363_ _20366_/A _20366_/C vssd1 vssd1 vccd1 vccd1 _20364_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22102_ _22791_/B vssd1 vssd1 vccd1 vccd1 _22792_/A sky130_fd_sc_hd__inv_2
XFILLER_0_114_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23082_ _16933_/B _22421_/A _23076_/X _23077_/Y _23081_/X vssd1 vssd1 vccd1 vccd1
+ _23083_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_28_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20294_ _21141_/C vssd1 vssd1 vccd1 vccd1 _21144_/B sky130_fd_sc_hd__inv_2
XFILLER_0_80_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22033_ _22058_/A _22033_/B vssd1 vssd1 vccd1 vccd1 _22033_/Y sky130_fd_sc_hd__nand2_1
Xhold2710 _25460_/Q vssd1 vssd1 vccd1 vccd1 _15546_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2721 _24973_/Q vssd1 vssd1 vccd1 vccd1 _12599_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2732 _26244_/Q vssd1 vssd1 vccd1 vccd1 hold2732/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2743 _24751_/X vssd1 vssd1 vccd1 vccd1 _24752_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2754 _25653_/Q vssd1 vssd1 vccd1 vccd1 hold2754/X sky130_fd_sc_hd__dlygate4sd3_1
X_23984_ _23984_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23985_/A sky130_fd_sc_hd__and2_1
XFILLER_0_138_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25723_ _25729_/CLK _25723_/D vssd1 vssd1 vccd1 vccd1 _25723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22935_ _22935_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _22935_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25654_ _26248_/CLK _25654_/D vssd1 vssd1 vccd1 vccd1 _25654_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_167_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22866_ _22866_/A _22866_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22868_/A sky130_fd_sc_hd__or3_1
XFILLER_0_74_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24605_ _24605_/A vssd1 vssd1 vccd1 vccd1 _26264_/D sky130_fd_sc_hd__clkbuf_1
X_21817_ _23087_/A _22601_/A vssd1 vssd1 vccd1 vccd1 _21825_/A sky130_fd_sc_hd__nand2_1
X_25585_ _26121_/CLK _25585_/D vssd1 vssd1 vccd1 vccd1 _25585_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_183_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22797_ _15384_/B _22680_/X _14273_/X vssd1 vssd1 vccd1 vccd1 _22797_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24536_ _24536_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24537_/A sky130_fd_sc_hd__and2_1
X_12550_ _17707_/B _17742_/A _17674_/A vssd1 vssd1 vccd1 vccd1 _12550_/Y sky130_fd_sc_hd__o21ai_1
X_21748_ _25838_/Q _25774_/Q vssd1 vssd1 vccd1 vccd1 _21749_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_148_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24467_ hold2584/X _26220_/Q _24510_/S vssd1 vssd1 vccd1 vccd1 _24467_/X sky130_fd_sc_hd__mux2_1
X_21679_ _21679_/A _21679_/B vssd1 vssd1 vccd1 vccd1 _21680_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_163_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26206_ _26207_/CLK _26206_/D vssd1 vssd1 vccd1 vccd1 _26206_/Q sky130_fd_sc_hd__dfxtp_1
X_14220_ _18814_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14220_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_151_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23418_ _23414_/Y _23417_/Y _24858_/S vssd1 vssd1 vccd1 vccd1 _23418_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_34_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24398_ _24398_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24399_/A sky130_fd_sc_hd__and2_1
XFILLER_0_61_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26137_ _26139_/CLK _26137_/D vssd1 vssd1 vccd1 vccd1 _26137_/Q sky130_fd_sc_hd__dfxtp_1
X_14151_ _25819_/Q vssd1 vssd1 vccd1 vccd1 _18592_/B sky130_fd_sc_hd__inv_2
X_23349_ _23349_/A vssd1 vssd1 vccd1 vccd1 _25932_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13102_ _17963_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13102_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26068_ _26069_/CLK _26068_/D vssd1 vssd1 vccd1 vccd1 _26068_/Q sky130_fd_sc_hd__dfxtp_1
X_14082_ _14118_/A hold789/X vssd1 vssd1 vccd1 vccd1 _14082_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_104_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17910_ _20747_/B _21731_/A vssd1 vssd1 vccd1 vccd1 _20740_/A sky130_fd_sc_hd__nand2_2
X_25019_ _26109_/CLK _25019_/D vssd1 vssd1 vccd1 vccd1 _25019_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ _13018_/X _13031_/X _13005_/X _13032_/X vssd1 vssd1 vccd1 vccd1 _13033_/X
+ sky130_fd_sc_hd__o211a_1
X_18890_ _18951_/A _18894_/B vssd1 vssd1 vccd1 vccd1 _18892_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17841_ _25856_/Q _22307_/A vssd1 vssd1 vccd1 vccd1 _17849_/A sky130_fd_sc_hd__or2_2
XFILLER_0_121_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14984_ _15033_/A _15032_/B _14983_/Y vssd1 vssd1 vccd1 vccd1 _14986_/A sky130_fd_sc_hd__a21o_1
X_17772_ _17781_/A _17774_/B vssd1 vssd1 vccd1 vccd1 _17773_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_89_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19511_ _19503_/X _19510_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19511_/Y sky130_fd_sc_hd__o21ai_1
X_16723_ _16721_/Y _16722_/Y _16594_/X vssd1 vssd1 vccd1 vccd1 _16723_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13935_ _13941_/A _13935_/B vssd1 vssd1 vccd1 vccd1 _13935_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16654_ _16654_/A vssd1 vssd1 vccd1 vccd1 _16655_/B sky130_fd_sc_hd__inv_2
X_19442_ _19441_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19443_/B
+ sky130_fd_sc_hd__a211o_1
X_13866_ _13941_/A _13866_/B vssd1 vssd1 vccd1 vccd1 _13866_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_18_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15605_ _15605_/A _15605_/B vssd1 vssd1 vccd1 vccd1 _15612_/B sky130_fd_sc_hd__nor2_1
X_12817_ _12746_/X _12815_/X _14910_/B _12816_/X vssd1 vssd1 vccd1 vccd1 _12817_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16585_ _16585_/A _16691_/B vssd1 vssd1 vccd1 vccd1 _16587_/A sky130_fd_sc_hd__nand2_1
X_19373_ _19373_/A _20909_/B vssd1 vssd1 vccd1 vccd1 _19373_/Y sky130_fd_sc_hd__nor2_1
X_13797_ _13823_/A _13797_/B vssd1 vssd1 vccd1 vccd1 _13797_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_151_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15536_ hold2623/X _15535_/Y _15464_/X vssd1 vssd1 vccd1 vccd1 _15536_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18324_ _18446_/A _25742_/Q _18952_/C vssd1 vssd1 vccd1 vccd1 _18325_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_139_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _14262_/B vssd1 vssd1 vccd1 vccd1 _12748_/X sky130_fd_sc_hd__clkbuf_16
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18255_ _21773_/B _25611_/Q vssd1 vssd1 vccd1 vccd1 _18257_/A sky130_fd_sc_hd__nand2_1
X_15467_ _15467_/A _15467_/B vssd1 vssd1 vccd1 vccd1 _15552_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_115_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12679_ _12679_/A vssd1 vssd1 vccd1 vccd1 _12684_/A sky130_fd_sc_hd__inv_2
XFILLER_0_25_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17206_ _25603_/Q vssd1 vssd1 vccd1 vccd1 _20818_/B sky130_fd_sc_hd__inv_2
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14418_ _14416_/Y hold138/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold139/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18186_ _18528_/A _18186_/B vssd1 vssd1 vccd1 vccd1 _18190_/A sky130_fd_sc_hd__nand2_1
X_15398_ _22815_/B _15398_/B vssd1 vssd1 vccd1 vccd1 _22812_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_181_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17137_ _17137_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17137_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_13_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14349_ _14688_/A vssd1 vssd1 vccd1 vccd1 _14404_/A sky130_fd_sc_hd__clkbuf_8
Xhold605 hold605/A vssd1 vssd1 vccd1 vccd1 hold605/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold616 hold616/A vssd1 vssd1 vccd1 vccd1 hold616/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 hold627/A vssd1 vssd1 vccd1 vccd1 hold627/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold638 hold638/A vssd1 vssd1 vccd1 vccd1 hold638/X sky130_fd_sc_hd__dlygate4sd3_1
X_17068_ _25650_/Q _17068_/B vssd1 vssd1 vccd1 vccd1 _17638_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_100_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold649 hold649/A vssd1 vssd1 vccd1 vccd1 hold649/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16019_ _16017_/X _16018_/Y _15805_/X vssd1 vssd1 vccd1 vccd1 _16019_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2006 _25998_/Q vssd1 vssd1 vccd1 vccd1 _14851_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2017 _24350_/X vssd1 vssd1 vccd1 vccd1 _24351_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2028 _12498_/X vssd1 vssd1 vccd1 vccd1 _24998_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2039 _26022_/Q vssd1 vssd1 vccd1 vccd1 hold2039/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1305 _21020_/Y vssd1 vssd1 vccd1 vccd1 _25801_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1316 _25727_/Q vssd1 vssd1 vccd1 vccd1 _19367_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1327 _25088_/Q vssd1 vssd1 vccd1 vccd1 _18475_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1338 _16807_/Y vssd1 vssd1 vccd1 vccd1 _25554_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1349 _25762_/Q vssd1 vssd1 vccd1 vccd1 _19865_/B sky130_fd_sc_hd__dlygate4sd3_1
X_19709_ _19723_/A _19709_/B vssd1 vssd1 vccd1 vccd1 _19709_/Y sky130_fd_sc_hd__nand2_1
X_20981_ _20981_/A _20981_/B _20981_/C vssd1 vssd1 vccd1 vccd1 _20982_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_170_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22720_ _22720_/A _22720_/B vssd1 vssd1 vccd1 vccd1 _22720_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22651_ _22651_/A _22651_/B vssd1 vssd1 vccd1 vccd1 _22652_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_149_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21602_ _21601_/Y _21203_/X _20986_/A _20957_/A vssd1 vssd1 vccd1 vccd1 _21602_/X
+ sky130_fd_sc_hd__a211o_1
X_25370_ _26198_/CLK hold145/X vssd1 vssd1 vccd1 vccd1 hold143/A sky130_fd_sc_hd__dfxtp_1
X_22582_ _22582_/A _23001_/B _22582_/C vssd1 vssd1 vccd1 vccd1 _22582_/X sky130_fd_sc_hd__and3_1
XFILLER_0_91_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24321_ _24321_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24322_/A sky130_fd_sc_hd__and2_1
XFILLER_0_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21533_ _21533_/A _21533_/B vssd1 vssd1 vccd1 vccd1 _21534_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24252_ hold2245/X hold2237/X _24279_/S vssd1 vssd1 vccd1 vccd1 _24253_/A sky130_fd_sc_hd__mux2_1
X_21464_ _21464_/A _21464_/B _21464_/C vssd1 vssd1 vccd1 vccd1 _21468_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_44_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23203_ _23212_/A _23203_/B vssd1 vssd1 vccd1 vccd1 _23204_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_114_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20415_ _21225_/B _21530_/A vssd1 vssd1 vccd1 vccd1 _20417_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_161_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24183_ _24183_/A vssd1 vssd1 vccd1 vccd1 _26127_/D sky130_fd_sc_hd__clkbuf_1
X_21395_ _21395_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21395_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23134_ _23132_/X _23133_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _23134_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20346_ _20346_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _20346_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_141_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23065_ _23065_/A _23193_/B _23065_/C vssd1 vssd1 vccd1 vccd1 _23065_/X sky130_fd_sc_hd__and3_1
X_20277_ _20277_/A _22302_/B _20277_/C vssd1 vssd1 vccd1 vccd1 _20281_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22016_ _18411_/A _25810_/Q _22014_/Y _22015_/Y vssd1 vssd1 vccd1 vccd1 _22017_/B
+ sky130_fd_sc_hd__a31o_1
Xhold2540 _12696_/Y vssd1 vssd1 vccd1 vccd1 _12697_/C sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2551 _25443_/Q vssd1 vssd1 vccd1 vccd1 _15238_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2562 _24820_/X vssd1 vssd1 vccd1 vccd1 _24821_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2573 _26224_/Q vssd1 vssd1 vccd1 vccd1 hold2573/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2584 _26219_/Q vssd1 vssd1 vccd1 vccd1 hold2584/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1850 _25840_/Q vssd1 vssd1 vccd1 vccd1 _21828_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2595 _24719_/X vssd1 vssd1 vccd1 vccd1 _24720_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1861 _24388_/X vssd1 vssd1 vccd1 vccd1 _24389_/A sky130_fd_sc_hd__dlygate4sd3_1
X_23967_ _23967_/A vssd1 vssd1 vccd1 vccd1 _26057_/D sky130_fd_sc_hd__clkbuf_1
Xhold1872 _25846_/Q vssd1 vssd1 vccd1 vccd1 _22033_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1883 _22114_/Y vssd1 vssd1 vccd1 vccd1 _25849_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1894 _22202_/Y vssd1 vssd1 vccd1 vccd1 _25852_/D sky130_fd_sc_hd__dlygate4sd3_1
X_25706_ _26335_/CLK _25706_/D vssd1 vssd1 vccd1 vccd1 _25706_/Q sky130_fd_sc_hd__dfxtp_4
X_13720_ _18489_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13720_/Y sky130_fd_sc_hd__nor2_1
X_22918_ _22918_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _22918_/Y sky130_fd_sc_hd__nand2_1
X_23898_ hold2061/X hold2048/X _23907_/S vssd1 vssd1 vccd1 vccd1 _23899_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_169_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13651_ _25739_/Q vssd1 vssd1 vccd1 vccd1 _18263_/B sky130_fd_sc_hd__inv_2
X_25637_ _26151_/CLK _25637_/D vssd1 vssd1 vccd1 vccd1 _25637_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_169_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22849_ _23191_/C vssd1 vssd1 vccd1 vccd1 _22849_/X sky130_fd_sc_hd__buf_6
XFILLER_0_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12602_ _12610_/A _23377_/B _12602_/C vssd1 vssd1 vccd1 vccd1 _12603_/A sky130_fd_sc_hd__and3b_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ hold914/X _16371_/A vssd1 vssd1 vccd1 vccd1 _16370_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_149_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25568_ _25573_/CLK _25568_/D vssd1 vssd1 vccd1 vccd1 _25568_/Q sky130_fd_sc_hd__dfxtp_1
X_13582_ _26231_/Q _13426_/X _13468_/X _13581_/Y vssd1 vssd1 vccd1 vccd1 _13583_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15321_ _15321_/A _15321_/B vssd1 vssd1 vccd1 vccd1 _15326_/A sky130_fd_sc_hd__or2_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12533_ _12533_/A _24745_/A vssd1 vssd1 vccd1 vccd1 _12533_/X sky130_fd_sc_hd__and2_1
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24519_ _24519_/A vssd1 vssd1 vccd1 vccd1 _26236_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25499_ _26341_/CLK hold862/X vssd1 vssd1 vccd1 vccd1 hold861/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18040_ _20856_/B _19345_/A vssd1 vssd1 vccd1 vccd1 _18041_/B sky130_fd_sc_hd__nand2_1
X_15252_ _15252_/A _15252_/B vssd1 vssd1 vccd1 vccd1 _15252_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_109_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14203_ _26330_/Q _13518_/B _14170_/X _14202_/Y vssd1 vssd1 vccd1 vccd1 _14204_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15183_ _15181_/X hold2527/X _15090_/X vssd1 vssd1 vccd1 vccd1 _15183_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14134_ _18530_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14134_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_123_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19991_ _26276_/Q hold725/X vssd1 vssd1 vccd1 vccd1 _19991_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_162_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14065_ _25805_/Q vssd1 vssd1 vccd1 vccd1 _18308_/B sky130_fd_sc_hd__inv_2
X_18942_ _18940_/X _18879_/X _18941_/X vssd1 vssd1 vccd1 vccd1 _18943_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_24_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13016_ _17564_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13016_/X sky130_fd_sc_hd__or2_1
X_18873_ _18955_/A _18873_/B _18894_/C vssd1 vssd1 vccd1 vccd1 _18874_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_146_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17824_ _20067_/B _25647_/Q vssd1 vssd1 vccd1 vccd1 _17828_/A sky130_fd_sc_hd__nand2_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14967_ _14967_/A _14967_/B vssd1 vssd1 vccd1 vccd1 _15033_/A sky130_fd_sc_hd__nand2_2
X_17755_ _17711_/A _25902_/Q _17831_/B vssd1 vssd1 vccd1 vccd1 _17874_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_89_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16706_ _16857_/B _16706_/B vssd1 vssd1 vccd1 vccd1 _16706_/Y sky130_fd_sc_hd__nand2_1
X_13918_ hold737/X _13916_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold738/A sky130_fd_sc_hd__a21oi_1
X_14898_ _25860_/Q _13466_/A _14897_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14899_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17686_ _17686_/A _23208_/A vssd1 vssd1 vccd1 vccd1 _17692_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_77_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19425_ _19423_/Y _19424_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19425_/Y sky130_fd_sc_hd__a21oi_1
X_16637_ _16635_/Y _16636_/Y _16594_/X vssd1 vssd1 vccd1 vccd1 hold949/A sky130_fd_sc_hd__a21oi_1
X_13849_ hold781/X _13848_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold782/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19356_ _26230_/Q hold786/X vssd1 vssd1 vccd1 vccd1 _19356_/Y sky130_fd_sc_hd__nand2_1
X_16568_ _16698_/A hold910/X vssd1 vssd1 vccd1 vccd1 _16568_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18307_ _18952_/A _18307_/B _18952_/C vssd1 vssd1 vccd1 vccd1 _18308_/C sky130_fd_sc_hd__nand3_1
X_15519_ _15956_/A hold878/X vssd1 vssd1 vccd1 vccd1 _15519_/Y sky130_fd_sc_hd__nand2_1
X_16499_ _16501_/B _16501_/A vssd1 vssd1 vccd1 vccd1 _16500_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_127_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19287_ _19286_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19288_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_154_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18238_ _25866_/Q _21737_/A vssd1 vssd1 vccd1 vccd1 _18246_/A sky130_fd_sc_hd__or2_2
XFILLER_0_167_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18169_ _18446_/A _19481_/B _18952_/C vssd1 vssd1 vccd1 vccd1 _18170_/C sky130_fd_sc_hd__nand3_1
Xhold402 hold402/A vssd1 vssd1 vccd1 vccd1 hold402/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold413 hold413/A vssd1 vssd1 vccd1 vccd1 hold413/X sky130_fd_sc_hd__dlygate4sd3_1
X_20200_ _20200_/A _20200_/B vssd1 vssd1 vccd1 vccd1 _20204_/A sky130_fd_sc_hd__nand2_1
Xhold424 hold424/A vssd1 vssd1 vccd1 vccd1 hold424/X sky130_fd_sc_hd__dlygate4sd3_1
X_21180_ _21180_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21180_/Y sky130_fd_sc_hd__nand2_1
Xhold435 hold435/A vssd1 vssd1 vccd1 vccd1 hold435/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 hold446/A vssd1 vssd1 vccd1 vccd1 hold446/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_25_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold457 hold457/A vssd1 vssd1 vccd1 vccd1 hold457/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold468 hold468/A vssd1 vssd1 vccd1 vccd1 hold468/X sky130_fd_sc_hd__dlygate4sd3_1
X_20131_ _20131_/A _22179_/B vssd1 vssd1 vccd1 vccd1 _20132_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold479 hold479/A vssd1 vssd1 vccd1 vccd1 hold479/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20062_ _20062_/A _20062_/B _20062_/C vssd1 vssd1 vccd1 vccd1 _20063_/B sky130_fd_sc_hd__nand3_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 _12981_/X vssd1 vssd1 vccd1 vccd1 _25046_/D sky130_fd_sc_hd__dlygate4sd3_1
X_24870_ _24870_/A _24870_/B vssd1 vssd1 vccd1 vccd1 _24870_/Y sky130_fd_sc_hd__nand2_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 _25065_/Q vssd1 vssd1 vccd1 vccd1 _17653_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1124 _16814_/Y vssd1 vssd1 vccd1 vccd1 _25555_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1135 _25079_/Q vssd1 vssd1 vccd1 vccd1 _18293_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 _16758_/Y vssd1 vssd1 vccd1 vccd1 _25547_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23821_ _23821_/A vssd1 vssd1 vccd1 vccd1 _26011_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1157 _25721_/Q vssd1 vssd1 vccd1 vccd1 _19283_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1168 _14865_/Y vssd1 vssd1 vccd1 vccd1 _25407_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 _25557_/Q vssd1 vssd1 vccd1 vccd1 _16827_/B sky130_fd_sc_hd__buf_1
XFILLER_0_139_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23752_ _23752_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23753_/A sky130_fd_sc_hd__and2_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20964_ _20964_/A _21972_/B vssd1 vssd1 vccd1 vccd1 _20965_/A sky130_fd_sc_hd__nand2_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22703_ _22703_/A _22703_/B vssd1 vssd1 vccd1 vccd1 _22705_/A sky130_fd_sc_hd__xor2_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23683_ _23683_/A vssd1 vssd1 vccd1 vccd1 _25966_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20895_ _21692_/A _21464_/C vssd1 vssd1 vccd1 vccd1 _20897_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25422_ _25422_/CLK _25422_/D vssd1 vssd1 vccd1 vccd1 _25422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22634_ _16764_/B _22421_/X _22628_/X _22629_/Y _22633_/X vssd1 vssd1 vccd1 vccd1
+ _22635_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_137_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25353_ _26308_/CLK hold361/X vssd1 vssd1 vccd1 vccd1 hold359/A sky130_fd_sc_hd__dfxtp_1
X_22565_ _18836_/A _25831_/Q _22563_/Y _22564_/Y vssd1 vssd1 vccd1 vccd1 _22566_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24304_ _24304_/A vssd1 vssd1 vccd1 vccd1 _26166_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21516_ _21516_/A _21516_/B _21516_/C vssd1 vssd1 vccd1 vccd1 _21517_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_91_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25284_ _26235_/CLK hold52/X vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22496_ _22496_/A _23039_/A vssd1 vssd1 vccd1 vccd1 _22498_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24235_ _24235_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24236_/A sky130_fd_sc_hd__and2_1
XFILLER_0_134_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21447_ _21498_/A _21450_/A vssd1 vssd1 vccd1 vccd1 _21448_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_160_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24166_ hold2046/X _26122_/Q _24203_/S vssd1 vssd1 vccd1 vccd1 _24166_/X sky130_fd_sc_hd__mux2_1
X_21378_ _21378_/A _21378_/B vssd1 vssd1 vccd1 vccd1 _21379_/A sky130_fd_sc_hd__nand2_1
X_23117_ _23197_/A _23117_/B vssd1 vssd1 vccd1 vccd1 _23117_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_102_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20329_ _20329_/A _20329_/B vssd1 vssd1 vccd1 vccd1 _20331_/A sky130_fd_sc_hd__nand2_1
X_24097_ _24097_/A vssd1 vssd1 vccd1 vccd1 _26099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold980 hold980/A vssd1 vssd1 vccd1 vccd1 hold980/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 hold991/A vssd1 vssd1 vccd1 vccd1 hold991/X sky130_fd_sc_hd__dlygate4sd3_1
X_23048_ _23047_/A _22849_/X _23047_/B vssd1 vssd1 vccd1 vccd1 _23049_/C sky130_fd_sc_hd__o21ai_1
X_15870_ _15857_/B _15869_/A _15856_/A vssd1 vssd1 vccd1 vccd1 _15870_/Y sky130_fd_sc_hd__o21ai_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2370 _12613_/Y vssd1 vssd1 vccd1 vccd1 _12618_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14821_ _14821_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14821_/Y sky130_fd_sc_hd__nand2_1
Xhold2381 _25671_/Q vssd1 vssd1 vccd1 vccd1 _13227_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2392 _26182_/Q vssd1 vssd1 vccd1 vccd1 hold2392/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24999_ _25860_/CLK hold7/X vssd1 vssd1 vccd1 vccd1 _24999_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1680 _22839_/Y vssd1 vssd1 vccd1 vccd1 _25879_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ _15839_/A _14752_/B vssd1 vssd1 vccd1 vccd1 _21934_/A sky130_fd_sc_hd__nand2_1
Xhold1691 _22757_/Y vssd1 vssd1 vccd1 vccd1 _25874_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17540_ _17538_/Y _17539_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _17540_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _13703_/A _13703_/B vssd1 vssd1 vccd1 vccd1 _13703_/Y sky130_fd_sc_hd__nand2_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17471_ _17624_/A _17471_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17471_/X sky130_fd_sc_hd__and3_1
XFILLER_0_86_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14683_ _14681_/Y hold147/X _14646_/X vssd1 vssd1 vccd1 vccd1 hold148/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19210_ _19211_/B _19211_/A vssd1 vssd1 vccd1 vccd1 _19210_/X sky130_fd_sc_hd__or2_1
X_16422_ _16473_/A hold894/X vssd1 vssd1 vccd1 vccd1 _16422_/Y sky130_fd_sc_hd__nand2_1
X_13634_ _13703_/A _13634_/B vssd1 vssd1 vccd1 vccd1 _13634_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_168_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16353_ _16473_/A hold968/X vssd1 vssd1 vccd1 vccd1 _16353_/Y sky130_fd_sc_hd__nand2_1
X_19141_ _20309_/A _22026_/A _25590_/Q vssd1 vssd1 vccd1 vccd1 _20314_/C sky130_fd_sc_hd__nand3_2
X_13565_ _13583_/A _13565_/B vssd1 vssd1 vccd1 vccd1 _13565_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_137_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15304_ _15305_/B _15305_/A vssd1 vssd1 vccd1 vccd1 _15306_/A sky130_fd_sc_hd__or2_1
XFILLER_0_171_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12516_ _24050_/B _12503_/A _12515_/X vssd1 vssd1 vccd1 vccd1 _24050_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_137_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19072_ _19070_/Y _19071_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25707_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16284_ _16284_/A vssd1 vssd1 vccd1 vccd1 _16297_/B sky130_fd_sc_hd__inv_2
XFILLER_0_136_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13496_ _13583_/A _13496_/B vssd1 vssd1 vccd1 vccd1 _13496_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15235_ _15221_/X _15266_/B _15234_/Y vssd1 vssd1 vccd1 vccd1 _15235_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18023_ _20216_/B _18023_/B vssd1 vssd1 vccd1 vccd1 _19177_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_164_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15166_ _15184_/B _15166_/B vssd1 vssd1 vccd1 vccd1 _15167_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_22_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14117_ hold588/X _14116_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold589/A sky130_fd_sc_hd__a21oi_1
X_15097_ _22425_/B _15810_/B vssd1 vssd1 vccd1 vccd1 _16146_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19974_ _19969_/X _19973_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19974_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14048_ _26305_/Q _13988_/X _13981_/X _14047_/Y vssd1 vssd1 vccd1 vccd1 _14049_/B
+ sky130_fd_sc_hd__a22o_1
X_18925_ _18922_/Y _18923_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25690_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18856_ _18856_/A _20751_/A vssd1 vssd1 vccd1 vccd1 _19045_/A sky130_fd_sc_hd__xor2_4
X_17807_ _17807_/A _17807_/B vssd1 vssd1 vccd1 vccd1 _22277_/A sky130_fd_sc_hd__nand2_1
X_18787_ _18787_/A _18787_/B vssd1 vssd1 vccd1 vccd1 _22512_/A sky130_fd_sc_hd__nand2_1
X_15999_ _15999_/A _15999_/B vssd1 vssd1 vccd1 vccd1 _16054_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_179_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17738_ _17738_/A vssd1 vssd1 vccd1 vccd1 _17738_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17669_ _25656_/Q vssd1 vssd1 vccd1 vccd1 _22076_/B sky130_fd_sc_hd__inv_2
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19408_ _19406_/X _19407_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19408_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20680_ _20680_/A _20680_/B vssd1 vssd1 vccd1 vccd1 _20682_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_174_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19339_ _19452_/A _19339_/B vssd1 vssd1 vccd1 vccd1 _19339_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22350_ _22350_/A _22350_/B vssd1 vssd1 vccd1 vccd1 _22350_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_171_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21301_ _21710_/B _21659_/C vssd1 vssd1 vccd1 vccd1 _21302_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22281_ _19275_/A _22280_/A _22280_/Y vssd1 vssd1 vccd1 vccd1 _22283_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24020_ hold2420/X _26075_/Q _24047_/S vssd1 vssd1 vccd1 vccd1 _24020_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold210 hold210/A vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
X_21232_ _21636_/A _21232_/B _21231_/X vssd1 vssd1 vccd1 vccd1 _21233_/B sky130_fd_sc_hd__or3b_1
Xhold221 hold221/A vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold232 hold232/A vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 hold243/A vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold254 hold254/A vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 hold265/A vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
X_21163_ _21163_/A _21163_/B vssd1 vssd1 vccd1 vccd1 _21165_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_180_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold276 hold276/A vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 hold287/A vssd1 vssd1 vccd1 vccd1 hold287/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold298 hold298/A vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
X_20114_ _20114_/A _20114_/B vssd1 vssd1 vccd1 vccd1 _20115_/B sky130_fd_sc_hd__xor2_2
X_25971_ _26041_/CLK _25971_/D vssd1 vssd1 vccd1 vccd1 _25971_/Q sky130_fd_sc_hd__dfxtp_1
X_21094_ _21093_/Y _20192_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21094_/X
+ sky130_fd_sc_hd__a211o_1
X_24922_ hold904/A hold910/A _24922_/S vssd1 vssd1 vccd1 vccd1 _24923_/B sky130_fd_sc_hd__mux2_1
X_20045_ _20048_/A _20048_/C vssd1 vssd1 vccd1 vccd1 _20047_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_176_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24853_ _15403_/B _15425_/B _24860_/S vssd1 vssd1 vccd1 vccd1 _24853_/X sky130_fd_sc_hd__mux2_1
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23804_ _23804_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23805_/A sky130_fd_sc_hd__and2_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24784_ hold2676/X hold2410/X _24817_/S vssd1 vssd1 vccd1 vccd1 _24785_/A sky130_fd_sc_hd__mux2_1
X_21996_ _21996_/A _21996_/B _23010_/A vssd1 vssd1 vccd1 vccd1 _21996_/Y sky130_fd_sc_hd__nand3_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23735_ _23735_/A vssd1 vssd1 vccd1 vccd1 _25983_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ _21497_/C vssd1 vssd1 vccd1 vccd1 _21500_/B sky130_fd_sc_hd__inv_2
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23666_ _23666_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23667_/A sky130_fd_sc_hd__and2_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20878_ _20878_/A _20878_/B vssd1 vssd1 vccd1 vccd1 _20879_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_138_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25405_ _25999_/CLK _25405_/D vssd1 vssd1 vccd1 vccd1 _25405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22617_ _22617_/A _22617_/B vssd1 vssd1 vccd1 vccd1 _22617_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_119_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23597_ _23597_/A _24967_/Q _23597_/C vssd1 vssd1 vccd1 vccd1 _23598_/B sky130_fd_sc_hd__and3_1
XFILLER_0_14_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25336_ _25797_/CLK hold133/X vssd1 vssd1 vccd1 vccd1 hold131/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13350_ _26193_/Q _13239_/X _13349_/X vssd1 vssd1 vccd1 vccd1 _13350_/X sky130_fd_sc_hd__a21o_1
X_22548_ _22923_/A _23072_/B vssd1 vssd1 vccd1 vccd1 _22549_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_84_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25267_ _26221_/CLK hold280/X vssd1 vssd1 vccd1 vccd1 hold278/A sky130_fd_sc_hd__dfxtp_1
X_13281_ _18699_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13281_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22479_ _22479_/A _22479_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22481_/A sky130_fd_sc_hd__or3_1
XFILLER_0_122_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15020_ _15018_/X _15019_/Y _14928_/X vssd1 vssd1 vccd1 vccd1 _25426_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24218_ _24218_/A vssd1 vssd1 vccd1 vccd1 _26138_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25198_ _25779_/CLK hold559/X vssd1 vssd1 vccd1 vccd1 hold557/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24149_ _24149_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24150_/A sky130_fd_sc_hd__and2_1
XFILLER_0_130_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16971_ _16969_/Y _16970_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _16971_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18710_ _18793_/A _25761_/Q _18891_/C vssd1 vssd1 vccd1 vccd1 _18711_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15922_ _15909_/B _15921_/A _15908_/A vssd1 vssd1 vccd1 vccd1 _15922_/Y sky130_fd_sc_hd__o21ai_1
X_19690_ _19706_/B _19779_/B vssd1 vssd1 vccd1 vccd1 _19692_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18641_ _18641_/A _19458_/A vssd1 vssd1 vccd1 vccd1 _18641_/Y sky130_fd_sc_hd__nand2_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15853_ _21759_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _15855_/A sky130_fd_sc_hd__nand2_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14804_ _14900_/A _14804_/B vssd1 vssd1 vccd1 vccd1 _14804_/Y sky130_fd_sc_hd__nand2_1
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18572_ _18572_/A _18572_/B _18572_/C vssd1 vssd1 vccd1 vccd1 _22239_/A sky130_fd_sc_hd__nand3_2
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15784_ _15784_/A _15786_/A vssd1 vssd1 vccd1 vccd1 _15784_/Y sky130_fd_sc_hd__nand2_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ _12930_/X _12994_/X _12917_/X _12995_/X vssd1 vssd1 vccd1 vccd1 _12996_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ _17523_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17523_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_157_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14735_ _21864_/B _15778_/B vssd1 vssd1 vccd1 vccd1 _14736_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_143_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14666_ _14666_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _14666_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ _17452_/Y _17453_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _17454_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16405_ _16416_/A _16406_/A vssd1 vssd1 vccd1 vccd1 _16405_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13617_ hold600/X _13616_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold601/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17385_ _17385_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17385_/Y sky130_fd_sc_hd__nand2_1
X_14597_ _14645_/A hold158/X vssd1 vssd1 vccd1 vccd1 hold159/A sky130_fd_sc_hd__nand2_1
XFILLER_0_184_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19124_ _19124_/A _19994_/B _19124_/C vssd1 vssd1 vccd1 vccd1 _19124_/X sky130_fd_sc_hd__and3_1
X_16336_ _16336_/A _16336_/B vssd1 vssd1 vccd1 vccd1 _16336_/Y sky130_fd_sc_hd__nor2_1
X_13548_ _13642_/A hold581/X vssd1 vssd1 vccd1 vccd1 hold582/A sky130_fd_sc_hd__nand2_1
XFILLER_0_153_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16267_ _16473_/A hold999/X vssd1 vssd1 vccd1 vccd1 _16267_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19055_ _19053_/X _18879_/X _19054_/X vssd1 vssd1 vccd1 vccd1 _19056_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_152_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13479_ hold498/X _13478_/Y _12558_/B vssd1 vssd1 vccd1 vccd1 hold499/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15218_ _15218_/A _15218_/B vssd1 vssd1 vccd1 vccd1 _15218_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_140_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18006_ _19066_/A _18454_/A vssd1 vssd1 vccd1 vccd1 _18007_/B sky130_fd_sc_hd__xnor2_2
X_16198_ _16190_/Y _16188_/Y _16214_/A vssd1 vssd1 vccd1 vccd1 _16208_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15149_ _15149_/A _15149_/B vssd1 vssd1 vccd1 vccd1 _15149_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_2_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19957_ _26273_/Q _19134_/X hold780/X vssd1 vssd1 vccd1 vccd1 _19958_/C sky130_fd_sc_hd__a21o_1
X_18908_ _18908_/A _18908_/B vssd1 vssd1 vccd1 vccd1 _22664_/A sky130_fd_sc_hd__or2_1
X_19888_ _19888_/A _19888_/B vssd1 vssd1 vccd1 vccd1 _19888_/Y sky130_fd_sc_hd__nand2_1
X_18839_ _19026_/A _18839_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18839_/X sky130_fd_sc_hd__and3_1
XFILLER_0_179_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21850_ _21850_/A _21850_/B vssd1 vssd1 vccd1 vccd1 _22626_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_78_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20801_ _21693_/B vssd1 vssd1 vccd1 vccd1 _21692_/B sky130_fd_sc_hd__inv_2
XFILLER_0_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21781_ _22575_/A vssd1 vssd1 vccd1 vccd1 _22073_/A sky130_fd_sc_hd__inv_2
XFILLER_0_78_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23520_ hold185/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23520_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_147_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20732_ _26295_/Q _20731_/X hold718/X vssd1 vssd1 vccd1 vccd1 _20735_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23451_ hold122/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23451_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_147_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20663_ _20663_/A _20663_/B vssd1 vssd1 vccd1 vccd1 _20666_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_133_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22402_ _22402_/A _23103_/A _22402_/C vssd1 vssd1 vccd1 vccd1 _22402_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_46_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26170_ _26171_/CLK _26170_/D vssd1 vssd1 vccd1 vccd1 _26170_/Q sky130_fd_sc_hd__dfxtp_1
X_23382_ _24863_/S vssd1 vssd1 vccd1 vccd1 _23391_/A sky130_fd_sc_hd__buf_12
X_20594_ _20594_/A _20594_/B vssd1 vssd1 vccd1 vccd1 _21335_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25121_ _26330_/CLK _25121_/D vssd1 vssd1 vccd1 vccd1 _25121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22333_ _22333_/A _22333_/B vssd1 vssd1 vccd1 vccd1 _22924_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_143_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25052_ _26135_/CLK _25052_/D vssd1 vssd1 vccd1 vccd1 _25052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22264_ _22262_/X _15839_/B _22263_/Y _14852_/A _21725_/X vssd1 vssd1 vccd1 vccd1
+ _22265_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24003_ _24003_/A vssd1 vssd1 vccd1 vccd1 _26069_/D sky130_fd_sc_hd__clkbuf_1
X_21215_ _21217_/B _21217_/C vssd1 vssd1 vccd1 vccd1 _21216_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_143_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22195_ _22195_/A _22195_/B vssd1 vssd1 vccd1 vccd1 _22196_/B sky130_fd_sc_hd__nand2_2
X_21146_ _21146_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _21151_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25954_ _26021_/CLK _25954_/D vssd1 vssd1 vccd1 vccd1 _25954_/Q sky130_fd_sc_hd__dfxtp_1
X_21077_ _21077_/A _25868_/Q vssd1 vssd1 vccd1 vccd1 _21081_/B sky130_fd_sc_hd__nand2_1
X_24905_ _24903_/X _24904_/X _24946_/A vssd1 vssd1 vccd1 vccd1 _24905_/X sky130_fd_sc_hd__mux2_1
X_20028_ _20028_/A _20028_/B _20952_/B vssd1 vssd1 vccd1 vccd1 _20032_/A sky130_fd_sc_hd__nand3_1
X_25885_ _25901_/CLK _25885_/D vssd1 vssd1 vccd1 vccd1 _25885_/Q sky130_fd_sc_hd__dfxtp_2
X_12850_ _12840_/X _12848_/X _12827_/X _12849_/X vssd1 vssd1 vccd1 vccd1 _12850_/X
+ sky130_fd_sc_hd__o211a_1
X_24836_ _24836_/A _24836_/B vssd1 vssd1 vccd1 vccd1 _24837_/A sky130_fd_sc_hd__and2_1
XFILLER_0_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _17109_/B _14264_/A vssd1 vssd1 vccd1 vccd1 _12781_/X sky130_fd_sc_hd__or2_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24767_ _24767_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24768_/A sky130_fd_sc_hd__and2_1
X_21979_ _23168_/A vssd1 vssd1 vccd1 vccd1 _23167_/A sky130_fd_sc_hd__inv_2
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14520_ _14518_/Y hold9/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__a21oi_1
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23718_ _23718_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23719_/A sky130_fd_sc_hd__and2_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24698_ hold2613/X hold2602/X _24740_/S vssd1 vssd1 vccd1 vccd1 _24699_/A sky130_fd_sc_hd__mux2_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14449_/Y hold57/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23649_ _23649_/A vssd1 vssd1 vccd1 vccd1 _25955_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13402_ _26330_/Q _19788_/A vssd1 vssd1 vccd1 vccd1 _14657_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_25_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17170_ _20518_/B _25890_/Q _25826_/Q vssd1 vssd1 vccd1 vccd1 _17171_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_107_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14382_ _14382_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14382_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_187_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16121_ _22365_/B _16691_/B vssd1 vssd1 vccd1 vccd1 _16123_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25319_ _26252_/CLK hold196/X vssd1 vssd1 vccd1 vccd1 hold194/A sky130_fd_sc_hd__dfxtp_1
X_13333_ _18859_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13333_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_130_clk clkbuf_leaf_82_clk/A vssd1 vssd1 vccd1 vccd1 _26339_/CLK sky130_fd_sc_hd__clkbuf_16
X_26299_ _26299_/CLK _26299_/D vssd1 vssd1 vccd1 vccd1 _26299_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16052_ _16052_/A _16052_/B vssd1 vssd1 vccd1 vccd1 _16053_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13264_ _13207_/X _13262_/X _13192_/X _13263_/X vssd1 vssd1 vccd1 vccd1 _13264_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15003_ _15003_/A _15015_/B vssd1 vssd1 vccd1 vccd1 _15003_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13195_ _13195_/A vssd1 vssd1 vccd1 vccd1 _19317_/A sky130_fd_sc_hd__buf_4
X_19811_ _19809_/Y _19810_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19811_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19742_ _19741_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19743_/B
+ sky130_fd_sc_hd__a211o_1
X_16954_ _16952_/X _16711_/A _16953_/Y _25897_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16955_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_47_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15905_ _21899_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _15907_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_189_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19673_ _19673_/A _20236_/B vssd1 vssd1 vccd1 vccd1 _19673_/Y sky130_fd_sc_hd__nor2_1
X_16885_ _16885_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16885_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_197_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _26244_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_154_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18624_ _22327_/B _25629_/Q vssd1 vssd1 vccd1 vccd1 _18626_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_189_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15836_ _15836_/A _15836_/B vssd1 vssd1 vccd1 vccd1 _16274_/A sky130_fd_sc_hd__nand2_4
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18555_ _18555_/A _18555_/B vssd1 vssd1 vccd1 vccd1 _18555_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_188_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15767_ _15701_/A _15824_/B _15766_/Y vssd1 vssd1 vccd1 vccd1 _15787_/A sky130_fd_sc_hd__a21o_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12979_ _14064_/A vssd1 vssd1 vccd1 vccd1 _13133_/B sky130_fd_sc_hd__buf_8
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17506_ _17506_/A _17506_/B vssd1 vssd1 vccd1 vccd1 _17506_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_75_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14718_ _25840_/Q _12527_/A _14913_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14718_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18486_ _18793_/A _19695_/B _18891_/C vssd1 vssd1 vccd1 vccd1 _18487_/C sky130_fd_sc_hd__nand3_1
X_15698_ _15698_/A _15698_/B vssd1 vssd1 vccd1 vccd1 _15829_/A sky130_fd_sc_hd__nand2_1
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17437_ _17437_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17437_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14649_ _14688_/A hold287/X vssd1 vssd1 vccd1 vccd1 hold288/A sky130_fd_sc_hd__nand2_1
XFILLER_0_117_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_16 _23602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_27 _18966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_38 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_49 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17368_ _25616_/Q vssd1 vssd1 vccd1 vccd1 _21184_/B sky130_fd_sc_hd__inv_2
XFILLER_0_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19107_ _22786_/A vssd1 vssd1 vccd1 vccd1 _21789_/A sky130_fd_sc_hd__clkbuf_16
X_16319_ _16319_/A vssd1 vssd1 vccd1 vccd1 _16321_/A sky130_fd_sc_hd__inv_2
XFILLER_0_127_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_121_clk clkbuf_4_14__f_clk/X vssd1 vssd1 vccd1 vccd1 _26198_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17299_ _17467_/A _17299_/B vssd1 vssd1 vccd1 vccd1 _17299_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19038_ _19038_/A _19038_/B vssd1 vssd1 vccd1 vccd1 _19039_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21000_ _21002_/B vssd1 vssd1 vccd1 vccd1 _21001_/B sky130_fd_sc_hd__inv_2
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22951_ _16879_/B _22421_/X _22945_/X _22946_/Y _22950_/X vssd1 vssd1 vccd1 vccd1
+ _22952_/A sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_188_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _25743_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21902_ _21902_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _21902_/X sky130_fd_sc_hd__and2_1
X_25670_ _26303_/CLK _25670_/D vssd1 vssd1 vccd1 vccd1 _25670_/Q sky130_fd_sc_hd__dfxtp_1
X_22882_ _22882_/A _22882_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22884_/A sky130_fd_sc_hd__or3_1
XFILLER_0_78_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24621_ hold2608/X _26270_/Q _24664_/S vssd1 vssd1 vccd1 vccd1 _24621_/X sky130_fd_sc_hd__mux2_1
X_21833_ _21833_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _21833_/X sky130_fd_sc_hd__and2_1
X_24552_ _24552_/A vssd1 vssd1 vccd1 vccd1 _26247_/D sky130_fd_sc_hd__clkbuf_1
X_21764_ _25794_/Q _21764_/B vssd1 vssd1 vccd1 vccd1 _21764_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_66_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23503_ _24940_/S hold269/A _23502_/X vssd1 vssd1 vccd1 vccd1 _23503_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_136_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20715_ _23101_/B vssd1 vssd1 vccd1 vccd1 _22569_/B sky130_fd_sc_hd__inv_2
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24483_ hold2573/X _26225_/Q _24510_/S vssd1 vssd1 vccd1 vccd1 _24483_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_92_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21695_ _21695_/A _21695_/B vssd1 vssd1 vccd1 vccd1 _21696_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26222_ _26232_/CLK _26222_/D vssd1 vssd1 vccd1 vccd1 _26222_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_184_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23434_ _24956_/S hold251/A _23433_/X vssd1 vssd1 vccd1 vccd1 _23434_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20646_ _21629_/B vssd1 vssd1 vccd1 vccd1 _21628_/B sky130_fd_sc_hd__inv_4
XFILLER_0_116_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26153_ _26154_/CLK _26153_/D vssd1 vssd1 vccd1 vccd1 _26153_/Q sky130_fd_sc_hd__dfxtp_1
X_23365_ _23365_/A vssd1 vssd1 vccd1 vccd1 _23372_/A sky130_fd_sc_hd__inv_2
XFILLER_0_144_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_112_clk clkbuf_4_14__f_clk/X vssd1 vssd1 vccd1 vccd1 _26208_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_132_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20577_ _26291_/Q _20078_/X hold777/X vssd1 vssd1 vccd1 vccd1 _20580_/B sky130_fd_sc_hd__a21oi_1
X_25104_ _26190_/CLK _25104_/D vssd1 vssd1 vccd1 vccd1 _25104_/Q sky130_fd_sc_hd__dfxtp_1
X_22316_ _22317_/A _22317_/B _23186_/A vssd1 vssd1 vccd1 vccd1 _22316_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26084_ _26084_/CLK _26084_/D vssd1 vssd1 vccd1 vccd1 _26084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23296_ _23298_/B _23298_/A vssd1 vssd1 vccd1 vccd1 _23303_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_132_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25035_ _26119_/CLK _25035_/D vssd1 vssd1 vccd1 vccd1 _25035_/Q sky130_fd_sc_hd__dfxtp_1
X_22247_ _22247_/A _25854_/Q vssd1 vssd1 vccd1 vccd1 _22247_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_108_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22178_ _22178_/A _25880_/Q vssd1 vssd1 vccd1 vccd1 _22178_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_178_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21129_ _21129_/A _21129_/B vssd1 vssd1 vccd1 vccd1 _21132_/B sky130_fd_sc_hd__nand2_1
X_25937_ _25939_/CLK _25937_/D vssd1 vssd1 vccd1 vccd1 _25937_/Q sky130_fd_sc_hd__dfxtp_1
X_13951_ _25787_/Q vssd1 vssd1 vccd1 vccd1 _17945_/B sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_179_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _25783_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12902_ _26243_/Q _25612_/Q vssd1 vssd1 vccd1 vccd1 _14382_/A sky130_fd_sc_hd__xor2_1
X_16670_ _16670_/A _16670_/B vssd1 vssd1 vccd1 vccd1 _16671_/B sky130_fd_sc_hd__nand2_1
X_13882_ _14120_/A vssd1 vssd1 vccd1 vccd1 _13996_/B sky130_fd_sc_hd__buf_8
X_25868_ _26046_/CLK _25868_/D vssd1 vssd1 vccd1 vccd1 _25868_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_69_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15621_ _15621_/A _16548_/B vssd1 vssd1 vccd1 vccd1 _15624_/A sky130_fd_sc_hd__nor2_1
X_12833_ _17242_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12833_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24819_ _24819_/A vssd1 vssd1 vccd1 vccd1 _26334_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25799_ _25803_/CLK _25799_/D vssd1 vssd1 vccd1 vccd1 _25799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18340_ _21157_/B _19504_/A vssd1 vssd1 vccd1 vccd1 _18341_/B sky130_fd_sc_hd__nand2_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _15552_/A _15552_/B vssd1 vssd1 vccd1 vccd1 _15822_/A sky130_fd_sc_hd__and2_1
X_12764_ _12726_/B _14298_/A _12752_/X _25585_/Q vssd1 vssd1 vccd1 vccd1 _12764_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14503_ _14503_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14503_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15483_ _15470_/X _15502_/B _15482_/Y vssd1 vssd1 vccd1 vccd1 _15483_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18271_ _18268_/X _18269_/X _18270_/X vssd1 vssd1 vccd1 vccd1 _18272_/A sky130_fd_sc_hd__a21o_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _12713_/A _12696_/A vssd1 vssd1 vccd1 vccd1 _12699_/A sky130_fd_sc_hd__or2_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17222_ _25638_/Q vssd1 vssd1 vccd1 vccd1 _20673_/B sky130_fd_sc_hd__inv_2
X_14434_ _14434_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14434_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_108_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14365_ _14404_/A hold395/X vssd1 vssd1 vccd1 vccd1 hold396/A sky130_fd_sc_hd__nand2_1
X_17153_ _25599_/Q vssd1 vssd1 vccd1 vccd1 _20663_/B sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_103_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _25938_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16104_ _16104_/A _16106_/A vssd1 vssd1 vccd1 vccd1 _16158_/B sky130_fd_sc_hd__and2_1
XFILLER_0_12_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13316_ _13316_/A vssd1 vssd1 vccd1 vccd1 _19588_/A sky130_fd_sc_hd__clkbuf_8
X_17084_ _19176_/A _17084_/B vssd1 vssd1 vccd1 vccd1 _17645_/A sky130_fd_sc_hd__xor2_4
Xhold809 hold809/A vssd1 vssd1 vccd1 vccd1 hold809/X sky130_fd_sc_hd__dlygate4sd3_1
X_14296_ _14344_/A hold101/X vssd1 vssd1 vccd1 vccd1 hold102/A sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16035_ hold704/X vssd1 vssd1 vccd1 vccd1 _16038_/B sky130_fd_sc_hd__inv_2
XFILLER_0_150_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13247_ _13247_/A vssd1 vssd1 vccd1 vccd1 _19430_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_122_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13178_ _13049_/X _14545_/A _13067_/X _19275_/A vssd1 vssd1 vccd1 vccd1 _13178_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17986_ _18612_/A _25724_/Q _18083_/C vssd1 vssd1 vccd1 vccd1 _17987_/C sky130_fd_sc_hd__nand3_1
Xhold1509 _25580_/Q vssd1 vssd1 vccd1 vccd1 _15808_/A sky130_fd_sc_hd__dlygate4sd3_1
X_19725_ _26256_/Q _19134_/X hold365/X vssd1 vssd1 vccd1 vccd1 _19725_/Y sky130_fd_sc_hd__a21oi_1
X_16937_ _16937_/A _16937_/B vssd1 vssd1 vccd1 vccd1 _16937_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_165_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19656_ _26251_/Q hold377/X vssd1 vssd1 vccd1 vccd1 _19656_/Y sky130_fd_sc_hd__nand2_1
X_16868_ _16869_/B _16869_/A vssd1 vssd1 vccd1 vccd1 _16868_/X sky130_fd_sc_hd__or2_1
X_18607_ _25884_/Q _22296_/A vssd1 vssd1 vccd1 vccd1 _18615_/A sky130_fd_sc_hd__or2_2
XFILLER_0_177_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15819_ _15830_/A _15820_/A vssd1 vssd1 vccd1 vccd1 _15819_/X sky130_fd_sc_hd__or2_1
X_19587_ _19584_/Y _19587_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19587_/X sky130_fd_sc_hd__and3b_1
X_16799_ _16858_/A _16799_/B vssd1 vssd1 vccd1 vccd1 _16799_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_133_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18538_ _18641_/A _19388_/A vssd1 vssd1 vccd1 vccd1 _18538_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18469_ _18955_/A _18469_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18470_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_185_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20500_ _20499_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20500_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21480_ _21480_/A _21480_/B _21480_/C vssd1 vssd1 vccd1 vccd1 _21484_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_133_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20431_ _20431_/A _25849_/Q vssd1 vssd1 vccd1 vccd1 _20435_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23150_ _23148_/X _23149_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _23150_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20362_ _20362_/A _20362_/B vssd1 vssd1 vccd1 vccd1 _20366_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22101_ _22101_/A _22101_/B vssd1 vssd1 vccd1 vccd1 _22791_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_144_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23081_ _23081_/A _23193_/B _23081_/C vssd1 vssd1 vccd1 vccd1 _23081_/X sky130_fd_sc_hd__and3_1
X_20293_ _21481_/A _21141_/C vssd1 vssd1 vccd1 vccd1 _20298_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22032_ _22004_/X _22031_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _22032_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2700 _26266_/Q vssd1 vssd1 vccd1 vccd1 hold2700/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2711 _15561_/Y vssd1 vssd1 vccd1 vccd1 _25460_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2722 _26327_/Q vssd1 vssd1 vccd1 vccd1 hold2722/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2733 _26273_/Q vssd1 vssd1 vccd1 vccd1 hold2733/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2744 _26292_/Q vssd1 vssd1 vccd1 vccd1 hold2744/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2755 _25901_/Q vssd1 vssd1 vccd1 vccd1 hold2755/X sky130_fd_sc_hd__dlygate4sd3_1
X_23983_ hold2178/X _26063_/Q _24001_/S vssd1 vssd1 vccd1 vccd1 _23983_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22934_ _16872_/B _22421_/X _22928_/X _22929_/Y _22933_/X vssd1 vssd1 vccd1 vccd1
+ _22935_/A sky130_fd_sc_hd__a221o_1
X_25722_ _25794_/CLK _25722_/D vssd1 vssd1 vccd1 vccd1 _25722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22865_ _26064_/Q vssd1 vssd1 vccd1 vccd1 _22866_/A sky130_fd_sc_hd__inv_2
X_25653_ _25743_/CLK _25653_/D vssd1 vssd1 vccd1 vccd1 _25653_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_39_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21816_ _21816_/A _21816_/B vssd1 vssd1 vccd1 vccd1 _22601_/A sky130_fd_sc_hd__nand2_2
X_24604_ _24604_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24605_/A sky130_fd_sc_hd__and2_1
X_25584_ _25587_/CLK _25584_/D vssd1 vssd1 vccd1 vccd1 _25584_/Q sky130_fd_sc_hd__dfxtp_2
X_22796_ _23188_/A _22796_/B vssd1 vssd1 vccd1 vccd1 _22796_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24535_ hold2626/X _26242_/Q _24587_/S vssd1 vssd1 vccd1 vccd1 _24535_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_94_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21747_ _22048_/A _23056_/A vssd1 vssd1 vccd1 vccd1 _21754_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_93_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24466_ _24466_/A vssd1 vssd1 vccd1 vccd1 _26219_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21678_ _21678_/A _21678_/B _21678_/C vssd1 vssd1 vccd1 vccd1 _21679_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_184_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26205_ _26205_/CLK _26205_/D vssd1 vssd1 vccd1 vccd1 _26205_/Q sky130_fd_sc_hd__dfxtp_1
X_23417_ _24940_/S hold362/A _23416_/X vssd1 vssd1 vccd1 vccd1 _23417_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20629_ _20631_/B _20631_/C vssd1 vssd1 vccd1 vccd1 _20630_/A sky130_fd_sc_hd__nand2_1
X_24397_ hold2514/X hold2363/X _24433_/S vssd1 vssd1 vccd1 vccd1 _24398_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_80_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26136_ _26136_/CLK _26136_/D vssd1 vssd1 vccd1 vccd1 _26136_/Q sky130_fd_sc_hd__dfxtp_1
X_14150_ _14236_/A hold825/X vssd1 vssd1 vccd1 vccd1 _14150_/Y sky130_fd_sc_hd__nand2_1
X_23348_ _23351_/A _23377_/B _23348_/C vssd1 vssd1 vccd1 vccd1 _23348_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13101_ _26152_/Q _13065_/X _13100_/X vssd1 vssd1 vccd1 vccd1 _13101_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26067_ _26069_/CLK _26067_/D vssd1 vssd1 vccd1 vccd1 _26067_/Q sky130_fd_sc_hd__dfxtp_1
X_14081_ hold489/X _14080_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold490/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23279_ _23279_/A _23377_/B _23284_/A vssd1 vssd1 vccd1 vccd1 _23279_/X sky130_fd_sc_hd__and3_1
XFILLER_0_120_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25018_ _26109_/CLK _25018_/D vssd1 vssd1 vccd1 vccd1 _25018_/Q sky130_fd_sc_hd__dfxtp_1
X_13032_ _17587_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13032_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17840_ _17840_/A _17840_/B vssd1 vssd1 vccd1 vccd1 _22307_/A sky130_fd_sc_hd__nand2_1
X_17771_ _17771_/A _17771_/B _17771_/C vssd1 vssd1 vccd1 vccd1 _17774_/B sky130_fd_sc_hd__nand3_2
X_14983_ _14962_/Y _14982_/A _14973_/B vssd1 vssd1 vccd1 vccd1 _14983_/Y sky130_fd_sc_hd__o21ai_1
X_19510_ _19508_/X _19509_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19510_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16722_ _16858_/A _16722_/B vssd1 vssd1 vccd1 vccd1 _16722_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13934_ _26287_/Q _13801_/X _13793_/X _13933_/Y vssd1 vssd1 vccd1 vccd1 _13935_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19441_ _26236_/Q hold599/X vssd1 vssd1 vccd1 vccd1 _19441_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_92_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16653_ hold942/X vssd1 vssd1 vccd1 vccd1 _16655_/A sky130_fd_sc_hd__inv_2
XFILLER_0_159_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13865_ _26276_/Q _13801_/X _13793_/X _13864_/Y vssd1 vssd1 vccd1 vccd1 _13866_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15604_ _15604_/A _16897_/A vssd1 vssd1 vccd1 vccd1 _15605_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12816_ _17200_/B _14264_/A vssd1 vssd1 vccd1 vccd1 _12816_/X sky130_fd_sc_hd__or2_1
X_19372_ _19369_/Y _19372_/B _19980_/B vssd1 vssd1 vccd1 vccd1 _19372_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16584_ hold962/X vssd1 vssd1 vccd1 vccd1 _16587_/B sky130_fd_sc_hd__inv_2
X_13796_ _26265_/Q _13612_/X _13793_/X _13795_/Y vssd1 vssd1 vccd1 vccd1 _13797_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18323_ _18445_/A _18327_/B vssd1 vssd1 vccd1 vccd1 _18325_/A sky130_fd_sc_hd__nand2_1
X_15535_ _15535_/A _15535_/B vssd1 vssd1 vccd1 vccd1 _15535_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_151_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _14120_/A vssd1 vssd1 vccd1 vccd1 _14262_/B sky130_fd_sc_hd__clkbuf_16
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ _19444_/A vssd1 vssd1 vccd1 vccd1 _21773_/B sky130_fd_sc_hd__inv_2
XFILLER_0_182_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12678_ _12678_/A vssd1 vssd1 vccd1 vccd1 _24987_/D sky130_fd_sc_hd__clkbuf_1
X_15466_ _15466_/A _15466_/B vssd1 vssd1 vccd1 vccd1 _15467_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_115_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17205_ _17202_/Y _17203_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _17205_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14417_ _14465_/A hold137/X vssd1 vssd1 vccd1 vccd1 hold138/A sky130_fd_sc_hd__nand2_1
XFILLER_0_181_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18185_ _25847_/Q _18185_/B _18184_/Y vssd1 vssd1 vccd1 vccd1 _18192_/A sky130_fd_sc_hd__or3b_2
XFILLER_0_170_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15397_ _15397_/A _15810_/B vssd1 vssd1 vccd1 vccd1 _15398_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17136_ _17134_/X _23187_/B _17135_/X vssd1 vssd1 vccd1 vccd1 _17137_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14348_ _14348_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14348_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold606 hold606/A vssd1 vssd1 vccd1 vccd1 hold606/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold617 hold617/A vssd1 vssd1 vccd1 vccd1 hold617/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold628 hold628/A vssd1 vssd1 vccd1 vccd1 hold628/X sky130_fd_sc_hd__dlygate4sd3_1
X_14279_ _14279_/A _14279_/B vssd1 vssd1 vccd1 vccd1 _14279_/Y sky130_fd_sc_hd__nand2_1
Xhold639 hold639/A vssd1 vssd1 vccd1 vccd1 hold639/X sky130_fd_sc_hd__dlygate4sd3_1
X_17067_ _20174_/B _25842_/Q _25778_/Q vssd1 vssd1 vccd1 vccd1 _17068_/B sky130_fd_sc_hd__mux2_2
X_16018_ _16212_/A _16018_/B vssd1 vssd1 vccd1 vccd1 _16018_/Y sky130_fd_sc_hd__nand2_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2007 _25935_/Q vssd1 vssd1 vccd1 vccd1 _23360_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2018 _25976_/Q vssd1 vssd1 vccd1 vccd1 hold2018/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2029 _25938_/Q vssd1 vssd1 vccd1 vccd1 _23376_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1306 _25572_/Q vssd1 vssd1 vccd1 vccd1 _16926_/B sky130_fd_sc_hd__clkbuf_2
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1317 _19368_/Y vssd1 vssd1 vccd1 vccd1 _25727_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1328 _13213_/X vssd1 vssd1 vccd1 vccd1 _25088_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17969_ _25650_/Q vssd1 vssd1 vccd1 vccd1 _21889_/A sky130_fd_sc_hd__inv_2
Xhold1339 _25061_/Q vssd1 vssd1 vccd1 vccd1 _17624_/B sky130_fd_sc_hd__dlygate4sd3_1
X_19708_ _19700_/X _19707_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19708_/Y sky130_fd_sc_hd__o21ai_1
X_20980_ _21467_/B _21513_/C vssd1 vssd1 vccd1 vccd1 _20981_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_177_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19639_ _19637_/Y _19638_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19639_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_178_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22650_ _22650_/A _22650_/B vssd1 vssd1 vccd1 vccd1 _22651_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_87_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21601_ _26333_/Q hold398/X vssd1 vssd1 vccd1 vccd1 _21601_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22581_ _22580_/A _22454_/X _22580_/B vssd1 vssd1 vccd1 vccd1 _22582_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24320_ hold2037/X _26172_/Q _24356_/S vssd1 vssd1 vccd1 vccd1 _24320_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21532_ _21532_/A _21532_/B _21532_/C vssd1 vssd1 vccd1 vccd1 _21533_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_157_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24251_ _24251_/A vssd1 vssd1 vccd1 vccd1 _26149_/D sky130_fd_sc_hd__clkbuf_1
X_21463_ _21514_/A _21466_/A vssd1 vssd1 vccd1 vccd1 _21464_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_141_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23202_ _23202_/A vssd1 vssd1 vccd1 vccd1 _25902_/D sky130_fd_sc_hd__inv_2
XFILLER_0_160_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20414_ _20414_/A _20414_/B _21141_/C vssd1 vssd1 vccd1 vccd1 _20418_/A sky130_fd_sc_hd__nand3_1
X_24182_ _24182_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24183_/A sky130_fd_sc_hd__and2_1
XFILLER_0_43_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21394_ _21394_/A _21394_/B vssd1 vssd1 vccd1 vccd1 _21395_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_120_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23133_ _23197_/A _23133_/B vssd1 vssd1 vccd1 vccd1 _23133_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_113_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20345_ _20345_/A _20345_/B vssd1 vssd1 vccd1 vccd1 _20346_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23064_ _23063_/A _22849_/X _23063_/B vssd1 vssd1 vccd1 vccd1 _23065_/C sky130_fd_sc_hd__o21ai_1
X_20276_ _22920_/B vssd1 vssd1 vccd1 vccd1 _22302_/B sky130_fd_sc_hd__inv_2
XFILLER_0_45_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22015_ _25810_/Q _22015_/B vssd1 vssd1 vccd1 vccd1 _22015_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2530 _25700_/Q vssd1 vssd1 vccd1 vccd1 _13407_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2541 _12697_/X vssd1 vssd1 vccd1 vccd1 _12698_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2552 _15251_/X vssd1 vssd1 vccd1 vccd1 hold2552/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2563 _26240_/Q vssd1 vssd1 vccd1 vccd1 hold2563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2574 _24483_/X vssd1 vssd1 vccd1 vccd1 _24484_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1840 _12550_/Y vssd1 vssd1 vccd1 vccd1 hold1840/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2585 _24467_/X vssd1 vssd1 vccd1 vccd1 _24469_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1851 _21829_/Y vssd1 vssd1 vccd1 vccd1 _25840_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2596 _26291_/Q vssd1 vssd1 vccd1 vccd1 hold2596/X sky130_fd_sc_hd__dlygate4sd3_1
X_23966_ _23966_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23967_/A sky130_fd_sc_hd__and2_1
Xhold1862 _25630_/Q vssd1 vssd1 vccd1 vccd1 _17546_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1873 _22034_/Y vssd1 vssd1 vccd1 vccd1 _25846_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1884 _25413_/Q vssd1 vssd1 vccd1 vccd1 _14916_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1895 _25983_/Q vssd1 vssd1 vccd1 vccd1 _14714_/B sky130_fd_sc_hd__dlygate4sd3_1
X_25705_ _26335_/CLK _25705_/D vssd1 vssd1 vccd1 vccd1 _25705_/Q sky130_fd_sc_hd__dfxtp_4
X_22917_ _16865_/B _22421_/X _22911_/X _22912_/Y _22916_/X vssd1 vssd1 vccd1 vccd1
+ _22918_/A sky130_fd_sc_hd__a221o_1
X_23897_ _23897_/A vssd1 vssd1 vccd1 vccd1 _26036_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22848_ _22848_/A _22848_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22851_/A sky130_fd_sc_hd__or3_1
XFILLER_0_39_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13650_ _13760_/A hold416/X vssd1 vssd1 vccd1 vccd1 hold417/A sky130_fd_sc_hd__nand2_1
X_25636_ _25636_/CLK _25636_/D vssd1 vssd1 vccd1 vccd1 _25636_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12601_/A _12644_/A vssd1 vssd1 vccd1 vccd1 _12602_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_112_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13581_ _17846_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13581_/Y sky130_fd_sc_hd__nor2_1
X_22779_ _23188_/A _22779_/B vssd1 vssd1 vccd1 vccd1 _22779_/X sky130_fd_sc_hd__or2_1
X_25567_ _26069_/CLK _25567_/D vssd1 vssd1 vccd1 vccd1 _25567_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15320_ _16787_/A _15320_/B vssd1 vssd1 vccd1 vccd1 _15321_/B sky130_fd_sc_hd__and2_1
X_12532_ _24745_/A vssd1 vssd1 vccd1 vccd1 _23629_/B sky130_fd_sc_hd__clkbuf_16
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24518_ _24518_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24519_/A sky130_fd_sc_hd__and2_1
XFILLER_0_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25498_ _25919_/CLK hold965/X vssd1 vssd1 vccd1 vccd1 hold964/A sky130_fd_sc_hd__dfxtp_1
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15251_ _15252_/B _15252_/A vssd1 vssd1 vccd1 vccd1 _15251_/X sky130_fd_sc_hd__or2_1
XFILLER_0_152_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24449_ hold2737/X hold2726/X _24510_/S vssd1 vssd1 vccd1 vccd1 _24450_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_62_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14202_ _18754_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14202_/Y sky130_fd_sc_hd__nor2_1
X_15182_ _15182_/A _15182_/B vssd1 vssd1 vccd1 vccd1 _15182_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_151_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14133_ _25816_/Q vssd1 vssd1 vccd1 vccd1 _18530_/B sky130_fd_sc_hd__inv_2
XFILLER_0_104_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26119_ _26119_/CLK _26119_/D vssd1 vssd1 vccd1 vccd1 _26119_/Q sky130_fd_sc_hd__dfxtp_1
X_19990_ _19990_/A _19990_/B vssd1 vssd1 vccd1 vccd1 _19990_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14064_ _14064_/A vssd1 vssd1 vccd1 vccd1 _14180_/A sky130_fd_sc_hd__clkbuf_8
X_18941_ _19026_/A _18941_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18941_/X sky130_fd_sc_hd__and3_1
XFILLER_0_24_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13015_ _26136_/Q _12907_/X _13014_/X vssd1 vssd1 vccd1 vccd1 _13015_/X sky130_fd_sc_hd__a21o_1
X_18872_ _18954_/A _25769_/Q vssd1 vssd1 vccd1 vccd1 _18874_/A sky130_fd_sc_hd__nand2_1
X_17823_ _17821_/Y _17822_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _25646_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
X_17754_ _17773_/B _17829_/A vssd1 vssd1 vccd1 vccd1 _17831_/B sky130_fd_sc_hd__nand2_1
X_14966_ _14946_/B _14964_/B _14956_/B vssd1 vssd1 vccd1 vccd1 _14967_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16705_ _21874_/B _13467_/A _15100_/A vssd1 vssd1 vccd1 vccd1 _16706_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13917_ _14345_/A vssd1 vssd1 vccd1 vccd1 _13917_/X sky130_fd_sc_hd__buf_8
XFILLER_0_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17685_ _17685_/A _17706_/A _17685_/C vssd1 vssd1 vccd1 vccd1 _23208_/A sky130_fd_sc_hd__nand3_1
X_14897_ _25860_/Q _12527_/A _15083_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14897_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19424_ _19452_/A _19424_/B vssd1 vssd1 vccd1 vccd1 _19424_/Y sky130_fd_sc_hd__nand2_1
X_16636_ _16698_/A hold948/X vssd1 vssd1 vccd1 vccd1 _16636_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13848_ _13941_/A _13848_/B vssd1 vssd1 vccd1 vccd1 _13848_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_175_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19355_ _26230_/Q _12537_/B hold786/X vssd1 vssd1 vccd1 vccd1 _19355_/Y sky130_fd_sc_hd__a21oi_1
X_16567_ _16565_/X _16566_/Y _16231_/A vssd1 vssd1 vccd1 vccd1 _16567_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_146_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13779_ _13774_/Y _13778_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold714/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18306_ _18951_/A hold981/X vssd1 vssd1 vccd1 vccd1 _18308_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15518_ _15505_/Y _15550_/A _15517_/Y vssd1 vssd1 vccd1 vccd1 _15518_/Y sky130_fd_sc_hd__o21ai_1
X_19286_ _26225_/Q hold419/X vssd1 vssd1 vccd1 vccd1 _19286_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16498_ _16498_/A _16691_/B vssd1 vssd1 vccd1 vccd1 _16501_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_183_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18237_ _18237_/A _18237_/B vssd1 vssd1 vccd1 vccd1 _21737_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_167_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15449_ _15449_/A vssd1 vssd1 vccd1 vccd1 _25454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18168_ _18529_/C vssd1 vssd1 vccd1 vccd1 _18952_/C sky130_fd_sc_hd__buf_8
XFILLER_0_81_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold403 hold403/A vssd1 vssd1 vccd1 vccd1 hold403/X sky130_fd_sc_hd__dlygate4sd3_1
X_17119_ _19715_/A _17119_/B vssd1 vssd1 vccd1 vccd1 _17541_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold414 hold414/A vssd1 vssd1 vccd1 vccd1 hold414/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 hold425/A vssd1 vssd1 vccd1 vccd1 hold425/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18099_ _18954_/A _25733_/Q vssd1 vssd1 vccd1 vccd1 _18102_/A sky130_fd_sc_hd__nand2_1
Xhold436 hold436/A vssd1 vssd1 vccd1 vccd1 hold436/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold447 hold447/A vssd1 vssd1 vccd1 vccd1 hold447/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold458 hold458/A vssd1 vssd1 vccd1 vccd1 hold458/X sky130_fd_sc_hd__dlygate4sd3_1
X_20130_ _20128_/Y _20129_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _20130_/Y sky130_fd_sc_hd__a21oi_1
Xhold469 hold469/A vssd1 vssd1 vccd1 vccd1 hold469/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20061_ _20061_/A _20061_/B vssd1 vssd1 vccd1 vccd1 _20063_/A sky130_fd_sc_hd__nand2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 _25043_/Q vssd1 vssd1 vccd1 vccd1 _17493_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 _13081_/X vssd1 vssd1 vccd1 vccd1 _25065_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1125 _25766_/Q vssd1 vssd1 vccd1 vccd1 _19917_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1136 _13157_/X vssd1 vssd1 vccd1 vccd1 _25079_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23820_ _23820_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23821_/A sky130_fd_sc_hd__and2_1
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1147 _25736_/Q vssd1 vssd1 vccd1 vccd1 _19498_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1158 _19284_/Y vssd1 vssd1 vccd1 vccd1 _25721_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 _25063_/Q vssd1 vssd1 vccd1 vccd1 _17639_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23751_ _14761_/B _14770_/B _23754_/S vssd1 vssd1 vccd1 vccd1 _23752_/A sky130_fd_sc_hd__mux2_1
X_20963_ _20961_/Y _20962_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _20963_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_92_clk clkbuf_leaf_95_clk/A vssd1 vssd1 vccd1 vccd1 _25919_/CLK sky130_fd_sc_hd__clkbuf_16
X_22702_ _22702_/A _22702_/B vssd1 vssd1 vccd1 vccd1 _22703_/B sky130_fd_sc_hd__nand2_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23682_ _23682_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23683_/A sky130_fd_sc_hd__and2_1
XFILLER_0_49_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20894_ _20894_/A _20894_/B _21419_/B vssd1 vssd1 vccd1 vccd1 _20898_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22633_ _22633_/A _23001_/B _22633_/C vssd1 vssd1 vccd1 vccd1 _22633_/X sky130_fd_sc_hd__and3_1
X_25421_ _25425_/CLK _25421_/D vssd1 vssd1 vccd1 vccd1 _25421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25352_ _26175_/CLK hold37/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfxtp_1
X_22564_ _25831_/Q _22564_/B vssd1 vssd1 vccd1 vccd1 _22564_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24303_ _24303_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24304_/A sky130_fd_sc_hd__and2_1
X_21515_ _21515_/A _21563_/A vssd1 vssd1 vccd1 vccd1 _21516_/C sky130_fd_sc_hd__nand2_1
X_25283_ _26235_/CLK hold364/X vssd1 vssd1 vccd1 vccd1 hold362/A sky130_fd_sc_hd__dfxtp_1
X_22495_ _23040_/B vssd1 vssd1 vccd1 vccd1 _23039_/A sky130_fd_sc_hd__inv_2
XFILLER_0_17_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24234_ hold2397/X hold2249/X _24279_/S vssd1 vssd1 vccd1 vccd1 _24235_/A sky130_fd_sc_hd__mux2_1
X_21446_ _21449_/A _21499_/A vssd1 vssd1 vccd1 vccd1 _21448_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24165_ _24165_/A vssd1 vssd1 vccd1 vccd1 _26121_/D sky130_fd_sc_hd__clkbuf_1
X_21377_ _21636_/A _21377_/B _21376_/X vssd1 vssd1 vccd1 vccd1 _21378_/B sky130_fd_sc_hd__or3b_2
XFILLER_0_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23116_ _23107_/Y _23115_/Y _19199_/A vssd1 vssd1 vccd1 vccd1 _23116_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20328_ _20330_/B vssd1 vssd1 vccd1 vccd1 _20329_/B sky130_fd_sc_hd__inv_2
X_24096_ _24096_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24097_/A sky130_fd_sc_hd__and2_1
Xhold970 hold970/A vssd1 vssd1 vccd1 vccd1 hold970/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 hold981/A vssd1 vssd1 vccd1 vccd1 hold981/X sky130_fd_sc_hd__dlygate4sd3_1
X_23047_ _23047_/A _23047_/B _23191_/C vssd1 vssd1 vccd1 vccd1 _23049_/A sky130_fd_sc_hd__or3_1
Xhold992 hold992/A vssd1 vssd1 vccd1 vccd1 hold992/X sky130_fd_sc_hd__dlygate4sd3_1
X_20259_ _20261_/A _20261_/B vssd1 vssd1 vccd1 vccd1 _20260_/A sky130_fd_sc_hd__nand2_1
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2360 _25920_/Q vssd1 vssd1 vccd1 vccd1 _23293_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2371 _12614_/X vssd1 vssd1 vccd1 vccd1 _12615_/A sky130_fd_sc_hd__dlygate4sd3_1
X_14820_ _25851_/Q _13466_/A _14819_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14821_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2382 _26104_/Q vssd1 vssd1 vccd1 vccd1 hold2382/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2393 _24353_/X vssd1 vssd1 vccd1 vccd1 _24354_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24998_ _26046_/CLK _24998_/D vssd1 vssd1 vccd1 vccd1 _24998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1670 _17337_/Y vssd1 vssd1 vccd1 vccd1 _25605_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ _14749_/Y _14750_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14751_/Y sky130_fd_sc_hd__a21oi_1
Xhold1681 _25831_/Q vssd1 vssd1 vccd1 vccd1 _21623_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23949_ _23949_/A vssd1 vssd1 vccd1 vccd1 _26051_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1692 _25756_/Q vssd1 vssd1 vccd1 vccd1 _19782_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_83_clk clkbuf_leaf_95_clk/A vssd1 vssd1 vccd1 vccd1 _26047_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _26250_/Q _13612_/X _13605_/X _13701_/Y vssd1 vssd1 vccd1 vccd1 _13703_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17470_ _17470_/A _17470_/B vssd1 vssd1 vccd1 vccd1 _17470_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_54_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682_ _14688_/A hold146/X vssd1 vssd1 vccd1 vccd1 hold147/A sky130_fd_sc_hd__nand2_1
X_16421_ _16421_/A _16697_/B _16428_/A vssd1 vssd1 vccd1 vccd1 _16421_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25619_ _25619_/CLK _25619_/D vssd1 vssd1 vccd1 vccd1 _25619_/Q sky130_fd_sc_hd__dfxtp_4
X_13633_ _26239_/Q _13612_/X _13605_/X _13632_/Y vssd1 vssd1 vccd1 vccd1 _13634_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19140_ _25654_/Q vssd1 vssd1 vccd1 vccd1 _22026_/A sky130_fd_sc_hd__inv_2
XFILLER_0_54_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16352_ _16350_/X _16351_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _16352_/X sky130_fd_sc_hd__a21o_1
X_13564_ _26228_/Q _13426_/X _13468_/X _13563_/Y vssd1 vssd1 vccd1 vccd1 _13565_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15303_ _16304_/A _16711_/A vssd1 vssd1 vccd1 vccd1 _15305_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_125_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12515_ _12515_/A _12515_/B _12515_/C vssd1 vssd1 vccd1 vccd1 _12515_/X sky130_fd_sc_hd__or3_2
X_19071_ _19186_/A _19071_/B vssd1 vssd1 vccd1 vccd1 _19071_/Y sky130_fd_sc_hd__nand2_1
X_16283_ _16285_/B _16285_/A vssd1 vssd1 vccd1 vccd1 _16284_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_164_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13495_ _26217_/Q _13426_/X _13468_/X _13494_/Y vssd1 vssd1 vccd1 vccd1 _13496_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18022_ _18022_/A _18022_/B vssd1 vssd1 vccd1 vccd1 _18023_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_87_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15234_ _15221_/X _15266_/B _15233_/X vssd1 vssd1 vccd1 vccd1 _15234_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15165_ _15165_/A _15165_/B vssd1 vssd1 vccd1 vccd1 _15166_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14116_ _14180_/A _14116_/B vssd1 vssd1 vccd1 vccd1 _14116_/Y sky130_fd_sc_hd__nand2_1
X_15096_ _15774_/B vssd1 vssd1 vccd1 vccd1 _15810_/B sky130_fd_sc_hd__clkbuf_16
X_19973_ _19971_/X _19972_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19973_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18924_ _21099_/A vssd1 vssd1 vccd1 vccd1 _18924_/X sky130_fd_sc_hd__clkbuf_8
X_14047_ _18244_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14047_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_158_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18855_ _20758_/B _22592_/A vssd1 vssd1 vccd1 vccd1 _20751_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_98_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17806_ _20663_/B _19275_/A vssd1 vssd1 vccd1 vccd1 _17807_/B sky130_fd_sc_hd__nand2_1
X_18786_ _20635_/B _19816_/A vssd1 vssd1 vccd1 vccd1 _18787_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15998_ _16026_/A vssd1 vssd1 vccd1 vccd1 _16006_/B sky130_fd_sc_hd__inv_2
X_17737_ _17737_/A _17737_/B vssd1 vssd1 vccd1 vccd1 _17771_/A sky130_fd_sc_hd__nand2_1
X_14949_ _14932_/B _14947_/B _14939_/B vssd1 vssd1 vccd1 vccd1 _14950_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_173_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17668_ _25656_/Q _20390_/B vssd1 vssd1 vccd1 vccd1 _17671_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_106_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19407_ _19407_/A _19407_/B vssd1 vssd1 vccd1 vccd1 _19407_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16619_ _16620_/A _16629_/B _16629_/A vssd1 vssd1 vccd1 vccd1 _16619_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_106_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17599_ _17597_/Y _17598_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _25637_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19338_ _19330_/X _19337_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19338_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19269_ _19267_/Y _19268_/Y _19086_/X vssd1 vssd1 vccd1 vccd1 _19269_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21300_ _21707_/C vssd1 vssd1 vccd1 vccd1 _21710_/B sky130_fd_sc_hd__inv_2
X_22280_ _22280_/A _22280_/B vssd1 vssd1 vccd1 vccd1 _22280_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_14_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold200 hold200/A vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__dlygate4sd3_1
X_21231_ _21230_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21231_/X
+ sky130_fd_sc_hd__a211o_1
Xhold211 hold211/A vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold222 hold222/A vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold233 hold233/A vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 hold244/A vssd1 vssd1 vccd1 vccd1 hold244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 hold255/A vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__dlygate4sd3_1
X_21162_ _21164_/C vssd1 vssd1 vccd1 vccd1 _21163_/B sky130_fd_sc_hd__inv_2
XFILLER_0_141_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold266 hold266/A vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold277 hold277/A vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 hold288/A vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20113_ _20113_/A _20113_/B vssd1 vssd1 vccd1 vccd1 _20114_/B sky130_fd_sc_hd__nand2_1
Xhold299 hold299/A vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
X_25970_ _26041_/CLK _25970_/D vssd1 vssd1 vccd1 vccd1 _25970_/Q sky130_fd_sc_hd__dfxtp_1
X_21093_ _26307_/Q hold796/X vssd1 vssd1 vccd1 vccd1 _21093_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_141_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24921_ _24946_/A _24921_/B vssd1 vssd1 vccd1 vccd1 _24921_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_176_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20044_ _20044_/A _20044_/B vssd1 vssd1 vccd1 vccd1 _20048_/A sky130_fd_sc_hd__nand2_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24852_ _24844_/X _24851_/X _24949_/S vssd1 vssd1 vccd1 vccd1 _24852_/X sky130_fd_sc_hd__mux2_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23803_ hold2067/X hold1967/X _23831_/S vssd1 vssd1 vccd1 vccd1 _23804_/A sky130_fd_sc_hd__mux2_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21995_ _21996_/A _21996_/B _23010_/A vssd1 vssd1 vccd1 vccd1 _21995_/X sky130_fd_sc_hd__a21o_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24783_ _24783_/A vssd1 vssd1 vccd1 vccd1 _26322_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_65_clk _25472_/CLK vssd1 vssd1 vccd1 vccd1 _26057_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23734_ _23734_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23735_/A sky130_fd_sc_hd__and2_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20946_ _21448_/C _21497_/C vssd1 vssd1 vccd1 vccd1 _20949_/A sky130_fd_sc_hd__nand2_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23665_ hold1993/X _25961_/Q _23677_/S vssd1 vssd1 vccd1 vccd1 _23665_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20877_ _21042_/A _20877_/B _20876_/X vssd1 vssd1 vccd1 vccd1 _20878_/B sky130_fd_sc_hd__or3b_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25404_ _25992_/CLK hold956/X vssd1 vssd1 vccd1 vccd1 hold955/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22616_ _18876_/A _25833_/Q _22614_/Y _22615_/Y vssd1 vssd1 vccd1 vccd1 _22617_/B
+ sky130_fd_sc_hd__a31o_1
X_23596_ _23923_/A _23596_/B _24970_/Q _24969_/Q vssd1 vssd1 vccd1 vccd1 _23599_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_187_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22547_ _23071_/B _22924_/A vssd1 vssd1 vccd1 vccd1 _22549_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25335_ _25797_/CLK hold322/X vssd1 vssd1 vccd1 vccd1 hold320/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13280_ _26182_/Q _13239_/X _13279_/X vssd1 vssd1 vccd1 vccd1 _13280_/X sky130_fd_sc_hd__a21o_1
X_22478_ _26046_/Q vssd1 vssd1 vccd1 vccd1 _22479_/A sky130_fd_sc_hd__inv_2
XFILLER_0_133_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25266_ _26219_/CLK hold13/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24217_ _24217_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24218_/A sky130_fd_sc_hd__and2_1
X_21429_ _21427_/Y _21428_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21429_/Y sky130_fd_sc_hd__a21oi_1
X_25197_ _26281_/CLK hold852/X vssd1 vssd1 vccd1 vccd1 hold851/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24148_ hold2284/X hold1955/X _24203_/S vssd1 vssd1 vccd1 vccd1 _24149_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16970_ _16977_/A _16970_/B vssd1 vssd1 vccd1 vccd1 _16970_/Y sky130_fd_sc_hd__nand2_1
X_24079_ _24079_/A vssd1 vssd1 vccd1 vccd1 _26093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15921_ _15921_/A _15921_/B vssd1 vssd1 vccd1 vccd1 _15941_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_21_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18640_ _18640_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18640_/Y sky130_fd_sc_hd__nand2_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15852_ hold692/X vssd1 vssd1 vccd1 vccd1 _15855_/B sky130_fd_sc_hd__inv_2
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2190 _24974_/Q vssd1 vssd1 vccd1 vccd1 _12643_/B sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_189_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ _14803_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14803_/Y sky130_fd_sc_hd__nand2_1
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ _18612_/A _18571_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18572_/C sky130_fd_sc_hd__nand3_1
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _15786_/A _15783_/B vssd1 vssd1 vccd1 vccd1 _15783_/X sky130_fd_sc_hd__or2_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_56_clk _25472_/CLK vssd1 vssd1 vccd1 vccd1 _25532_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12995_ _17536_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _12995_/X sky130_fd_sc_hd__or2_1
XFILLER_0_188_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ _17520_/X _17241_/X _17521_/X vssd1 vssd1 vccd1 vccd1 _17523_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14734_ _14740_/B _21865_/A vssd1 vssd1 vccd1 vccd1 _21864_/B sky130_fd_sc_hd__xnor2_2
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17453_ _17467_/A _17453_/B vssd1 vssd1 vccd1 vccd1 _17453_/Y sky130_fd_sc_hd__nand2_1
X_14665_ _14663_/Y hold39/X _14646_/X vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__a21oi_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16404_ _16404_/A _16404_/B vssd1 vssd1 vccd1 vccd1 _16406_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_145_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13616_ _13703_/A _13616_/B vssd1 vssd1 vccd1 vccd1 _13616_/Y sky130_fd_sc_hd__nand2_1
X_17384_ _17382_/X _17241_/X _17383_/X vssd1 vssd1 vccd1 vccd1 _17385_/A sky130_fd_sc_hd__a21o_1
X_14596_ _14596_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14596_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_156_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19123_ _26214_/Q _19483_/A hold497/X vssd1 vssd1 vccd1 vccd1 _19124_/C sky130_fd_sc_hd__a21o_1
X_16335_ _16335_/A vssd1 vssd1 vccd1 vccd1 _16380_/B sky130_fd_sc_hd__inv_2
X_13547_ hold420/X _13546_/Y _12558_/B vssd1 vssd1 vccd1 vccd1 hold421/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19054_ _19082_/A _19054_/B _22786_/A vssd1 vssd1 vccd1 vccd1 _19054_/X sky130_fd_sc_hd__and3_1
X_16266_ _16266_/A _16697_/B vssd1 vssd1 vccd1 vccd1 _16266_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13478_ _13583_/A _13478_/B vssd1 vssd1 vccd1 vccd1 _13478_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18005_ _18005_/A _20817_/A vssd1 vssd1 vccd1 vccd1 _18454_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_70_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15217_ _15218_/B _15218_/A vssd1 vssd1 vccd1 vccd1 _15217_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16197_ _16197_/A vssd1 vssd1 vccd1 vccd1 _16214_/A sky130_fd_sc_hd__inv_2
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15148_ _15149_/B _15149_/A vssd1 vssd1 vccd1 vccd1 _15148_/X sky130_fd_sc_hd__or2_1
XFILLER_0_121_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15079_ _15085_/B _15080_/A vssd1 vssd1 vccd1 vccd1 _15079_/X sky130_fd_sc_hd__or2_1
X_19956_ _19955_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19958_/A
+ sky130_fd_sc_hd__a211o_1
X_18907_ _25643_/Q _22665_/B vssd1 vssd1 vccd1 vccd1 _18908_/B sky130_fd_sc_hd__nor2_1
X_19887_ _19888_/B _19888_/A vssd1 vssd1 vccd1 vccd1 _19887_/X sky130_fd_sc_hd__or2_1
Xclkbuf_4_0__f_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _26093_/CLK sky130_fd_sc_hd__clkbuf_16
X_18838_ _18838_/A _18838_/B vssd1 vssd1 vccd1 vccd1 _18838_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_101_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18769_ _18792_/A _18773_/B vssd1 vssd1 vccd1 vccd1 _18771_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_47_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _26042_/CLK sky130_fd_sc_hd__clkbuf_16
X_20800_ _21416_/C _21693_/B vssd1 vssd1 vccd1 vccd1 _20803_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21780_ _23071_/A _22575_/A vssd1 vssd1 vccd1 vccd1 _21788_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20731_ _21228_/A vssd1 vssd1 vccd1 vccd1 _20731_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_175_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23450_ _23447_/Y _23449_/Y _24957_/S vssd1 vssd1 vccd1 vccd1 _23450_/X sky130_fd_sc_hd__mux2_1
X_20662_ _20662_/A _22278_/B vssd1 vssd1 vccd1 vccd1 _20663_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_147_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22401_ _22402_/A _22402_/C _23103_/A vssd1 vssd1 vccd1 vccd1 _22401_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_147_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23381_ _23379_/X hold477/X _12702_/A vssd1 vssd1 vccd1 vccd1 hold478/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20593_ _20592_/B _20593_/B _20593_/C vssd1 vssd1 vccd1 vccd1 _20594_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_61_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25120_ _26330_/CLK hold974/X vssd1 vssd1 vccd1 vccd1 hold973/A sky130_fd_sc_hd__dfxtp_1
X_22332_ _22332_/A _22332_/B vssd1 vssd1 vccd1 vccd1 _22333_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25051_ _25636_/CLK _25051_/D vssd1 vssd1 vccd1 vccd1 _25051_/Q sky130_fd_sc_hd__dfxtp_1
X_22263_ _22263_/A _22387_/B vssd1 vssd1 vccd1 vccd1 _22263_/Y sky130_fd_sc_hd__nand2_1
X_24002_ _24002_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _24003_/A sky130_fd_sc_hd__and2_1
XFILLER_0_131_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21214_ _25873_/Q _21214_/B _21214_/C vssd1 vssd1 vccd1 vccd1 _21217_/C sky130_fd_sc_hd__nand3b_1
X_22194_ _22195_/B _22195_/A vssd1 vssd1 vccd1 vccd1 _22196_/A sky130_fd_sc_hd__or2_2
XFILLER_0_111_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21145_ _21145_/A _21145_/B vssd1 vssd1 vccd1 vccd1 _21146_/A sky130_fd_sc_hd__nand2_1
X_25953_ _26021_/CLK _25953_/D vssd1 vssd1 vccd1 vccd1 _25953_/Q sky130_fd_sc_hd__dfxtp_1
X_21076_ _21078_/B _21078_/C vssd1 vssd1 vccd1 vccd1 _21077_/A sky130_fd_sc_hd__nand2_1
X_24904_ _15891_/B _15907_/B _24945_/S vssd1 vssd1 vccd1 vccd1 _24904_/X sky130_fd_sc_hd__mux2_1
X_20027_ _20949_/C vssd1 vssd1 vccd1 vccd1 _20952_/B sky130_fd_sc_hd__inv_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25884_ _26084_/CLK _25884_/D vssd1 vssd1 vccd1 vccd1 _25884_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24835_ hold2702/X hold2716/X _24835_/S vssd1 vssd1 vccd1 vccd1 _24836_/A sky130_fd_sc_hd__mux2_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_clk _25184_/CLK vssd1 vssd1 vccd1 vccd1 _26264_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12780_ _26091_/Q _12748_/X _12779_/X vssd1 vssd1 vccd1 vccd1 _12780_/X sky130_fd_sc_hd__a21o_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24766_ hold2589/X hold2532/X _24817_/S vssd1 vssd1 vccd1 vccd1 _24767_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_96_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21978_ _21978_/A _21978_/B vssd1 vssd1 vccd1 vccd1 _23168_/A sky130_fd_sc_hd__nand2_4
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23717_ hold2259/X hold2079/X _23754_/S vssd1 vssd1 vccd1 vccd1 _23718_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_139_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20929_ _20928_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20929_/X
+ sky130_fd_sc_hd__a211o_1
X_24697_ _24697_/A vssd1 vssd1 vccd1 vccd1 _26294_/D sky130_fd_sc_hd__clkbuf_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _14465_/A hold56/X vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__nand2_1
X_23648_ _23648_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23649_/A sky130_fd_sc_hd__and2_1
XFILLER_0_154_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13401_ _13401_/A vssd1 vssd1 vccd1 vccd1 _19788_/A sky130_fd_sc_hd__buf_6
XFILLER_0_181_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14381_ _14379_/Y hold108/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold109/A sky130_fd_sc_hd__a21oi_1
X_23579_ _23555_/X _24959_/A _23256_/B _23578_/X vssd1 vssd1 vccd1 vccd1 _23579_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16120_ hold644/X vssd1 vssd1 vccd1 vccd1 _16123_/B sky130_fd_sc_hd__inv_2
XFILLER_0_36_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25318_ _26252_/CLK hold193/X vssd1 vssd1 vccd1 vccd1 hold191/A sky130_fd_sc_hd__dfxtp_1
X_13332_ _26190_/Q _13239_/X _13331_/X vssd1 vssd1 vccd1 vccd1 _13332_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_106_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26298_ _26298_/CLK _26298_/D vssd1 vssd1 vccd1 vccd1 _26298_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_106_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16051_ _16084_/A vssd1 vssd1 vccd1 vccd1 _16062_/B sky130_fd_sc_hd__inv_2
XFILLER_0_161_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25249_ _25249_/CLK hold753/X vssd1 vssd1 vccd1 vccd1 hold751/A sky130_fd_sc_hd__dfxtp_1
X_13263_ _18638_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13263_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15002_ _15015_/B _15003_/A vssd1 vssd1 vccd1 vccd1 _15002_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13194_ _13109_/X _13191_/X _13192_/X _13193_/X vssd1 vssd1 vccd1 vccd1 _13194_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19810_ _19975_/A _19810_/B vssd1 vssd1 vccd1 vccd1 _19810_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_102_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16953_ _16953_/A _16953_/B vssd1 vssd1 vccd1 vccd1 _16953_/Y sky130_fd_sc_hd__nand2_1
X_19741_ _26257_/Q hold584/X vssd1 vssd1 vccd1 vccd1 _19741_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15904_ hold858/X vssd1 vssd1 vccd1 vccd1 _15907_/B sky130_fd_sc_hd__inv_2
X_19672_ _19669_/Y _19672_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19672_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16884_ _16882_/X _16711_/X _16883_/Y _25887_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16885_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_189_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18623_ _19701_/A vssd1 vssd1 vccd1 vccd1 _22327_/B sky130_fd_sc_hd__inv_2
X_15835_ _15828_/Y _15557_/Y _15834_/Y vssd1 vssd1 vccd1 vccd1 _15836_/B sky130_fd_sc_hd__a21oi_1
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_clk _25759_/CLK vssd1 vssd1 vccd1 vccd1 _25761_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_189_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18554_ _18758_/A _18899_/A vssd1 vssd1 vccd1 vccd1 _18555_/B sky130_fd_sc_hd__xnor2_1
X_15766_ _15764_/Y _15719_/X _15765_/Y vssd1 vssd1 vccd1 vccd1 _15766_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12978_ _26129_/Q _12907_/X _12977_/X vssd1 vssd1 vccd1 vccd1 _12978_/X sky130_fd_sc_hd__a21o_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _17505_/A _17555_/A vssd1 vssd1 vccd1 vccd1 _17506_/B sky130_fd_sc_hd__xnor2_1
X_14717_ _14717_/A vssd1 vssd1 vccd1 vccd1 _14913_/A sky130_fd_sc_hd__inv_2
XFILLER_0_87_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18485_ _18792_/A _18489_/B vssd1 vssd1 vccd1 vccd1 _18487_/A sky130_fd_sc_hd__nand2_1
X_15697_ _15659_/X _15693_/A _15696_/X vssd1 vssd1 vccd1 vccd1 _15698_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17436_ _17434_/X _17241_/X _17435_/X vssd1 vssd1 vccd1 vccd1 _17437_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_68_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14648_ _14648_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _14648_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 _18874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_28 _19031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17367_ _17365_/Y _17366_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _25608_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14579_ _14585_/A hold359/X vssd1 vssd1 vccd1 vccd1 hold360/A sky130_fd_sc_hd__nand2_1
XFILLER_0_103_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19106_ _19102_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19109_/A
+ sky130_fd_sc_hd__a211o_1
X_16318_ _16320_/B hold873/X vssd1 vssd1 vccd1 vccd1 _16319_/A sky130_fd_sc_hd__and2_1
XFILLER_0_55_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17298_ _17298_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17298_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19037_ _19035_/Y _19036_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25702_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16249_ _16250_/B _16250_/A vssd1 vssd1 vccd1 vccd1 _16264_/B sky130_fd_sc_hd__or2_1
XFILLER_0_140_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19939_ _19939_/A _19990_/A vssd1 vssd1 vccd1 vccd1 _19939_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_177_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22950_ _22950_/A _23001_/B _22950_/C vssd1 vssd1 vccd1 vccd1 _22950_/X sky130_fd_sc_hd__and3_1
XFILLER_0_173_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21901_ _21899_/X _14270_/A _21900_/Y _14750_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _21902_/A sky130_fd_sc_hd__a32o_1
X_22881_ _26065_/Q vssd1 vssd1 vccd1 vccd1 _22882_/A sky130_fd_sc_hd__inv_2
XFILLER_0_78_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24620_ _24620_/A vssd1 vssd1 vccd1 vccd1 _26269_/D sky130_fd_sc_hd__clkbuf_1
X_21832_ _21830_/X _14270_/A _21831_/Y _14731_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _21833_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21763_ _21763_/A _25858_/Q vssd1 vssd1 vccd1 vccd1 _21763_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24551_ _24551_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24552_/A sky130_fd_sc_hd__and2_1
XFILLER_0_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20714_ _20714_/A _25895_/Q vssd1 vssd1 vccd1 vccd1 _20720_/A sky130_fd_sc_hd__nand2_1
X_23502_ hold95/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23502_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_176_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24482_ _24482_/A vssd1 vssd1 vccd1 vccd1 _26224_/D sky130_fd_sc_hd__clkbuf_1
X_21694_ _21694_/A _21694_/B _21694_/C vssd1 vssd1 vccd1 vccd1 _21695_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26221_ _26221_/CLK _26221_/D vssd1 vssd1 vccd1 vccd1 _26221_/Q sky130_fd_sc_hd__dfxtp_2
X_23433_ hold47/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23433_/X sky130_fd_sc_hd__or2b_1
X_20645_ _21354_/B _21629_/B vssd1 vssd1 vccd1 vccd1 _20648_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_135_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23364_ _23366_/B _23366_/A vssd1 vssd1 vccd1 vccd1 _23365_/A sky130_fd_sc_hd__nor2_1
X_26152_ _26152_/CLK _26152_/D vssd1 vssd1 vccd1 vccd1 _26152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20576_ _20576_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20581_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25103_ _26317_/CLK _25103_/D vssd1 vssd1 vccd1 vccd1 _25103_/Q sky130_fd_sc_hd__dfxtp_1
X_22315_ _23039_/B vssd1 vssd1 vccd1 vccd1 _23186_/A sky130_fd_sc_hd__inv_2
X_23295_ _23307_/A _23306_/A vssd1 vssd1 vccd1 vccd1 _23298_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_143_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26083_ _26084_/CLK _26083_/D vssd1 vssd1 vccd1 vccd1 _26083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22246_ _22729_/A _22874_/B vssd1 vssd1 vccd1 vccd1 _22257_/C sky130_fd_sc_hd__nand2_1
X_25034_ _26119_/CLK _25034_/D vssd1 vssd1 vccd1 vccd1 _25034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22177_ _22177_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _22177_/X sky130_fd_sc_hd__and2_1
XFILLER_0_121_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21128_ _21128_/A _21878_/B vssd1 vssd1 vccd1 vccd1 _21129_/A sky130_fd_sc_hd__nand2_1
X_25936_ _25939_/CLK _25936_/D vssd1 vssd1 vccd1 vccd1 _25936_/Q sky130_fd_sc_hd__dfxtp_1
X_13950_ _14000_/A hold728/X vssd1 vssd1 vccd1 vccd1 hold729/A sky130_fd_sc_hd__nand2_1
X_21059_ _21059_/A _21059_/B _21059_/C vssd1 vssd1 vccd1 vccd1 _21063_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_89_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12901_ _12840_/X _12899_/X _12827_/X _12900_/X vssd1 vssd1 vccd1 vccd1 _12901_/X
+ sky130_fd_sc_hd__o211a_1
X_25867_ _25876_/CLK _25867_/D vssd1 vssd1 vccd1 vccd1 _25867_/Q sky130_fd_sc_hd__dfxtp_4
X_13881_ _20129_/B vssd1 vssd1 vccd1 vccd1 _17881_/B sky130_fd_sc_hd__inv_2
XFILLER_0_9_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15620_ _23012_/B _16369_/B vssd1 vssd1 vccd1 vccd1 _16548_/B sky130_fd_sc_hd__nand2_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24818_ _24818_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24819_/A sky130_fd_sc_hd__and2_1
XFILLER_0_115_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12832_ _26101_/Q _12748_/X _12831_/X vssd1 vssd1 vccd1 vccd1 _12832_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25798_ _25803_/CLK _25798_/D vssd1 vssd1 vccd1 vccd1 _25798_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_69_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15551_ _15551_/A _15551_/B vssd1 vssd1 vccd1 vccd1 _15552_/B sky130_fd_sc_hd__nor2_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12763_ _26216_/Q _25585_/Q vssd1 vssd1 vccd1 vccd1 _14298_/A sky130_fd_sc_hd__xor2_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24749_ _24749_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24750_/A sky130_fd_sc_hd__and2_1
XFILLER_0_96_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _14500_/Y hold135/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold136/A sky130_fd_sc_hd__a21oi_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _18535_/A _18270_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _18270_/X sky130_fd_sc_hd__and3_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15482_ _15470_/X _15502_/B _15233_/X vssd1 vssd1 vccd1 vccd1 _15482_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12694_ _12694_/A vssd1 vssd1 vccd1 vccd1 _12713_/A sky130_fd_sc_hd__inv_2
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _19345_/A _17221_/B vssd1 vssd1 vccd1 vccd1 _17520_/A sky130_fd_sc_hd__xor2_4
X_14433_ _14431_/Y hold171/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold172/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_166_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17152_ _17150_/Y _17151_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _25591_/D sky130_fd_sc_hd__a21oi_1
X_14364_ _14364_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14364_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16103_ _16103_/A _16103_/B vssd1 vssd1 vccd1 vccd1 _16106_/A sky130_fd_sc_hd__nor2_1
X_13315_ _14260_/A vssd1 vssd1 vccd1 vccd1 _13315_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17083_ _19176_/B _25843_/Q _25779_/Q vssd1 vssd1 vccd1 vccd1 _17084_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_161_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14295_ _14295_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14295_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16034_ _16032_/Y hold663/X _15805_/X vssd1 vssd1 vccd1 vccd1 hold664/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13246_ _13207_/X _13244_/X _13192_/X _13245_/X vssd1 vssd1 vccd1 vccd1 _13246_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13177_ _26294_/Q _19275_/A vssd1 vssd1 vccd1 vccd1 _14545_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_21_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17985_ _18611_/A _17989_/B vssd1 vssd1 vccd1 vccd1 _17987_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_165_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16936_ _16937_/B _16937_/A vssd1 vssd1 vccd1 vccd1 _16936_/X sky130_fd_sc_hd__or2_1
X_19724_ _19722_/Y _19723_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19724_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_189_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16867_ _16935_/A _16872_/B vssd1 vssd1 vccd1 vccd1 _16869_/B sky130_fd_sc_hd__nand2_1
X_19655_ _26251_/Q _19483_/X hold377/X vssd1 vssd1 vccd1 vccd1 _19655_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15818_ _15789_/Y _15830_/B _15800_/B vssd1 vssd1 vccd1 vccd1 _15820_/A sky130_fd_sc_hd__a21oi_1
X_18606_ _18606_/A _18606_/B vssd1 vssd1 vccd1 vccd1 _22296_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_133_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19586_ _19585_/Y _19272_/X _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19587_/B
+ sky130_fd_sc_hd__a211o_1
X_16798_ _16798_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16798_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18537_ _18537_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18537_/Y sky130_fd_sc_hd__nand2_1
X_15749_ _15750_/B _15750_/A vssd1 vssd1 vccd1 vccd1 _15749_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18468_ _18954_/A _25749_/Q vssd1 vssd1 vccd1 vccd1 _18470_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17419_ _25621_/Q vssd1 vssd1 vccd1 vccd1 _20011_/B sky130_fd_sc_hd__inv_2
XFILLER_0_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18399_ _22015_/B _25618_/Q vssd1 vssd1 vccd1 vccd1 _18401_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_172_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20430_ _20432_/B _20432_/C vssd1 vssd1 vccd1 vccd1 _20431_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20361_ _20361_/A _22348_/B vssd1 vssd1 vccd1 vccd1 _20362_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_9_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _26142_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_144_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22100_ _22100_/A _22805_/B vssd1 vssd1 vccd1 vccd1 _22101_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23080_ _23079_/A _22849_/X _23079_/B vssd1 vssd1 vccd1 vccd1 _23081_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20292_ _20292_/A _20292_/B vssd1 vssd1 vccd1 vccd1 _21141_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_144_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22031_ _22029_/X _22030_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _22031_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2701 _26257_/Q vssd1 vssd1 vccd1 vccd1 hold2701/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2712 _26329_/Q vssd1 vssd1 vccd1 vccd1 hold2712/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2723 _26222_/Q vssd1 vssd1 vccd1 vccd1 hold2723/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2734 _26282_/Q vssd1 vssd1 vccd1 vccd1 hold2734/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2745 _26307_/Q vssd1 vssd1 vccd1 vccd1 hold2745/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2756 _25656_/Q vssd1 vssd1 vccd1 vccd1 hold2756/X sky130_fd_sc_hd__dlygate4sd3_1
X_23982_ _23982_/A vssd1 vssd1 vccd1 vccd1 _26062_/D sky130_fd_sc_hd__clkbuf_1
X_25721_ _26236_/CLK _25721_/D vssd1 vssd1 vccd1 vccd1 _25721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22933_ _22933_/A _23001_/B _22933_/C vssd1 vssd1 vccd1 vccd1 _22933_/X sky130_fd_sc_hd__and3_1
XFILLER_0_39_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25652_ _25743_/CLK _25652_/D vssd1 vssd1 vccd1 vccd1 _25652_/Q sky130_fd_sc_hd__dfxtp_4
X_22864_ _15454_/B _22680_/X _22829_/X vssd1 vssd1 vccd1 vccd1 _22864_/Y sky130_fd_sc_hd__a21oi_1
X_24603_ hold2736/X hold2615/X _24664_/S vssd1 vssd1 vccd1 vccd1 _24604_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_149_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21815_ _21815_/A _22612_/B vssd1 vssd1 vccd1 vccd1 _21816_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_167_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25583_ _26121_/CLK _25583_/D vssd1 vssd1 vccd1 vccd1 _25583_/Q sky130_fd_sc_hd__dfxtp_2
X_22795_ _22795_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22795_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24534_ _24534_/A vssd1 vssd1 vccd1 vccd1 _26241_/D sky130_fd_sc_hd__clkbuf_1
X_21746_ _22550_/A vssd1 vssd1 vccd1 vccd1 _22048_/A sky130_fd_sc_hd__inv_2
XFILLER_0_94_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24465_ _24465_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24466_/A sky130_fd_sc_hd__and2_1
XFILLER_0_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21677_ _21677_/A _21677_/B vssd1 vssd1 vccd1 vccd1 _21678_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_47_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26204_ _26205_/CLK _26204_/D vssd1 vssd1 vccd1 vccd1 _26204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23416_ hold50/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23416_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_164_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20628_ _25854_/Q _20628_/B _20628_/C vssd1 vssd1 vccd1 vccd1 _20631_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24396_ _24396_/A vssd1 vssd1 vccd1 vccd1 _26196_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26135_ _26135_/CLK _26135_/D vssd1 vssd1 vccd1 vccd1 _26135_/Q sky130_fd_sc_hd__dfxtp_1
X_23347_ _23347_/A _23347_/B vssd1 vssd1 vccd1 vccd1 _23347_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20559_ _20562_/A _20562_/C vssd1 vssd1 vccd1 vccd1 _20560_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13100_ _13049_/X _14500_/A _13067_/X _25649_/Q vssd1 vssd1 vccd1 vccd1 _13100_/X
+ sky130_fd_sc_hd__a22o_1
X_26066_ _26066_/CLK _26066_/D vssd1 vssd1 vccd1 vccd1 _26066_/Q sky130_fd_sc_hd__dfxtp_1
X_14080_ _14180_/A _14080_/B vssd1 vssd1 vccd1 vccd1 _14080_/Y sky130_fd_sc_hd__nand2_1
X_23278_ _23278_/A _23278_/B _23278_/C vssd1 vssd1 vccd1 vccd1 _23284_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_21_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25017_ _26109_/CLK _25017_/D vssd1 vssd1 vccd1 vccd1 _25017_/Q sky130_fd_sc_hd__dfxtp_1
X_13031_ _26139_/Q _12907_/X _13030_/X vssd1 vssd1 vccd1 vccd1 _13031_/X sky130_fd_sc_hd__a21o_1
X_22229_ _22206_/X _22228_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _22229_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17770_ _17770_/A _17783_/C vssd1 vssd1 vccd1 vccd1 _17781_/A sky130_fd_sc_hd__nand2_2
X_14982_ _14982_/A _14982_/B vssd1 vssd1 vccd1 vccd1 _15032_/B sky130_fd_sc_hd__nor2_1
X_16721_ _16721_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16721_/Y sky130_fd_sc_hd__nand2_1
X_25919_ _25919_/CLK hold834/X vssd1 vssd1 vccd1 vccd1 hold832/A sky130_fd_sc_hd__dfxtp_1
X_13933_ _17801_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13933_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_156_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19440_ _26236_/Q _12537_/B hold599/X vssd1 vssd1 vccd1 vccd1 _19440_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16652_ hold942/X _16654_/A vssd1 vssd1 vccd1 vccd1 _16656_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_88_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13864_ _18955_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13864_/Y sky130_fd_sc_hd__nor2_1
X_15603_ _15603_/A vssd1 vssd1 vccd1 vccd1 _16897_/A sky130_fd_sc_hd__inv_2
X_19371_ _19370_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19372_/B
+ sky130_fd_sc_hd__a211o_1
X_12815_ _26098_/Q _12748_/X _12814_/X vssd1 vssd1 vccd1 vccd1 _12815_/X sky130_fd_sc_hd__a21o_1
X_16583_ _16581_/Y _16582_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 hold919/A sky130_fd_sc_hd__a21oi_1
X_13795_ _18733_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13795_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18322_ _25870_/Q _21877_/A vssd1 vssd1 vccd1 vccd1 _18330_/A sky130_fd_sc_hd__or2_2
X_15534_ _15535_/B _15535_/A vssd1 vssd1 vccd1 vccd1 _15534_/X sky130_fd_sc_hd__or2_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _14260_/A vssd1 vssd1 vccd1 vccd1 _12746_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_85_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ _18251_/Y _18252_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25657_/D sky130_fd_sc_hd__a21oi_1
X_15465_ _15462_/X hold2461/X _15464_/X vssd1 vssd1 vccd1 vccd1 _15465_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12677_ _12677_/A _24836_/B _12684_/B vssd1 vssd1 vccd1 vccd1 _12677_/X sky130_fd_sc_hd__and3_1
XFILLER_0_37_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17204_ _17568_/A vssd1 vssd1 vccd1 vccd1 _17204_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14416_ _14416_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14416_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18184_ _20350_/B _25655_/Q vssd1 vssd1 vccd1 vccd1 _18184_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_170_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15396_ _26021_/Q _25957_/Q _15773_/S vssd1 vssd1 vccd1 vccd1 _15397_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_154_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17135_ _17393_/A _25010_/Q _19994_/B vssd1 vssd1 vccd1 vccd1 _17135_/X sky130_fd_sc_hd__and3_1
XFILLER_0_4_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14347_ _14687_/B vssd1 vssd1 vccd1 vccd1 _14403_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold607 hold607/A vssd1 vssd1 vccd1 vccd1 hold607/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold618 hold618/A vssd1 vssd1 vccd1 vccd1 hold618/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold629 hold629/A vssd1 vssd1 vccd1 vccd1 hold629/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_64_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17066_ _25586_/Q vssd1 vssd1 vccd1 vccd1 _20174_/B sky130_fd_sc_hd__inv_2
X_14278_ _14279_/B _14279_/A vssd1 vssd1 vccd1 vccd1 _14278_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16017_ _16015_/X _16016_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _16017_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_111_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13229_ _13220_/X _14569_/A _13067_/X _19388_/A vssd1 vssd1 vccd1 vccd1 _13229_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2008 _23359_/X vssd1 vssd1 vccd1 vccd1 _23361_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2019 _23714_/X vssd1 vssd1 vccd1 vccd1 _23715_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1307 _16927_/Y vssd1 vssd1 vccd1 vccd1 _25572_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1318 _25395_/Q vssd1 vssd1 vccd1 vccd1 _14759_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17968_ _20174_/B _25650_/Q vssd1 vssd1 vccd1 vccd1 _17971_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_100_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1329 _25411_/Q vssd1 vssd1 vccd1 vccd1 _14900_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_19707_ _19705_/X _19706_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19707_/Y sky130_fd_sc_hd__a21oi_1
X_16919_ _16917_/Y _15656_/B _16918_/Y vssd1 vssd1 vccd1 vccd1 _16919_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17899_ _19303_/A vssd1 vssd1 vccd1 vccd1 _21729_/B sky130_fd_sc_hd__inv_2
XFILLER_0_178_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19638_ _19723_/A _19638_/B vssd1 vssd1 vccd1 vccd1 _19638_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_177_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19569_ _19567_/Y _19568_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 hold982/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21600_ _26333_/Q _19130_/X hold398/X vssd1 vssd1 vccd1 vccd1 _21603_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22580_ _22580_/A _22580_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22582_/A sky130_fd_sc_hd__or3_1
XFILLER_0_34_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21531_ _21531_/A _21579_/A vssd1 vssd1 vccd1 vccd1 _21532_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_91_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24250_ _24250_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24251_/A sky130_fd_sc_hd__and2_1
XFILLER_0_69_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21462_ _21465_/A _21515_/A vssd1 vssd1 vccd1 vccd1 _21464_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_160_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23201_ _23212_/A _23201_/B vssd1 vssd1 vccd1 vccd1 _23202_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20413_ _21530_/A _21222_/C vssd1 vssd1 vccd1 vccd1 _20414_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24181_ _26126_/Q hold2354/X _24203_/S vssd1 vssd1 vccd1 vccd1 _24181_/X sky130_fd_sc_hd__mux2_1
X_21393_ _21636_/A _21393_/B _21392_/X vssd1 vssd1 vccd1 vccd1 _21394_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_4_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23132_ _23123_/Y _23131_/Y _19199_/A vssd1 vssd1 vccd1 vccd1 _23132_/X sky130_fd_sc_hd__a21o_1
X_20344_ _21042_/A _20344_/B _20343_/X vssd1 vssd1 vccd1 vccd1 _20345_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23063_ _23063_/A _23063_/B _23191_/C vssd1 vssd1 vccd1 vccd1 _23065_/A sky130_fd_sc_hd__or3_1
X_20275_ _20275_/A _25884_/Q vssd1 vssd1 vccd1 vccd1 _20281_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_105_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22014_ _22014_/A _25874_/Q vssd1 vssd1 vccd1 vccd1 _22014_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2520 _17678_/Y vssd1 vssd1 vccd1 vccd1 _17679_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2531 _25701_/Q vssd1 vssd1 vccd1 vccd1 _13413_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2542 _25414_/Q vssd1 vssd1 vccd1 vccd1 _14913_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2553 _15253_/Y vssd1 vssd1 vccd1 vccd1 _25443_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2564 _24532_/X vssd1 vssd1 vccd1 vccd1 _24533_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1830 _17490_/Y vssd1 vssd1 vccd1 vccd1 _25622_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2575 _26258_/Q vssd1 vssd1 vccd1 vccd1 hold2575/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2586 _26267_/Q vssd1 vssd1 vccd1 vccd1 hold2586/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1841 _12557_/X vssd1 vssd1 vccd1 vccd1 _25581_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23965_ hold2390/X hold2357/X _24001_/S vssd1 vssd1 vccd1 vccd1 _23966_/A sky130_fd_sc_hd__mux2_1
Xhold1852 _25851_/Q vssd1 vssd1 vccd1 vccd1 _22171_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2597 _24689_/X vssd1 vssd1 vccd1 vccd1 _24690_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1863 _17547_/Y vssd1 vssd1 vccd1 vccd1 _25630_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1874 _25854_/Q vssd1 vssd1 vccd1 vccd1 _22260_/B sky130_fd_sc_hd__dlygate4sd3_1
X_25704_ _25708_/CLK _25704_/D vssd1 vssd1 vccd1 vccd1 _25704_/Q sky130_fd_sc_hd__dfxtp_4
X_22916_ _22916_/A _23001_/B _22916_/C vssd1 vssd1 vccd1 vccd1 _22916_/X sky130_fd_sc_hd__and3_1
Xhold1885 _14907_/Y vssd1 vssd1 vccd1 vccd1 _14909_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1896 _23736_/X vssd1 vssd1 vccd1 vccd1 _23737_/A sky130_fd_sc_hd__dlygate4sd3_1
X_23896_ _23896_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23897_/A sky130_fd_sc_hd__and2_1
XFILLER_0_155_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25635_ _25636_/CLK _25635_/D vssd1 vssd1 vccd1 vccd1 _25635_/Q sky130_fd_sc_hd__dfxtp_4
X_22847_ _26063_/Q vssd1 vssd1 vccd1 vccd1 _22848_/A sky130_fd_sc_hd__inv_2
XFILLER_0_184_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12600_ _12644_/A _12601_/A vssd1 vssd1 vccd1 vccd1 _12610_/A sky130_fd_sc_hd__nor2_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25566_ _26069_/CLK _25566_/D vssd1 vssd1 vccd1 vccd1 _25566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _25728_/Q vssd1 vssd1 vccd1 vccd1 _17846_/B sky130_fd_sc_hd__inv_2
XFILLER_0_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22778_ _22778_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22778_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12531_ _12724_/B _12529_/Y _12558_/B vssd1 vssd1 vccd1 vccd1 _25001_/D sky130_fd_sc_hd__a21oi_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24517_ hold2380/X hold1999/X _24587_/S vssd1 vssd1 vccd1 vccd1 _24518_/A sky130_fd_sc_hd__mux2_1
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21729_ _25793_/Q _21729_/B vssd1 vssd1 vccd1 vccd1 _21729_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_93_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25497_ _25919_/CLK hold646/X vssd1 vssd1 vccd1 vccd1 hold644/A sky130_fd_sc_hd__dfxtp_1
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15250_ _15221_/X _15266_/B _15232_/B vssd1 vssd1 vccd1 vccd1 _15252_/A sky130_fd_sc_hd__a21o_1
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24448_ _24448_/A vssd1 vssd1 vccd1 vccd1 _26213_/D sky130_fd_sc_hd__clkbuf_1
X_14201_ _25827_/Q vssd1 vssd1 vccd1 vccd1 _18754_/B sky130_fd_sc_hd__inv_2
XFILLER_0_124_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15181_ _15182_/B _15182_/A vssd1 vssd1 vccd1 vccd1 _15181_/X sky130_fd_sc_hd__or2_1
XFILLER_0_152_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24379_ hold2090/X _26191_/Q _24433_/S vssd1 vssd1 vccd1 vccd1 _24379_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_151_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26118_ _26119_/CLK _26118_/D vssd1 vssd1 vccd1 vccd1 _26118_/Q sky130_fd_sc_hd__dfxtp_1
X_14132_ _14236_/A hold731/X vssd1 vssd1 vccd1 vccd1 _14132_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26049_ _26051_/CLK _26049_/D vssd1 vssd1 vccd1 vccd1 _26049_/Q sky130_fd_sc_hd__dfxtp_1
X_14063_ _14118_/A hold620/X vssd1 vssd1 vccd1 vccd1 hold621/A sky130_fd_sc_hd__nand2_1
X_18940_ _18940_/A _18940_/B vssd1 vssd1 vccd1 vccd1 _18940_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13014_ _12891_/X _14449_/A _12909_/X _25633_/Q vssd1 vssd1 vccd1 vccd1 _13014_/X
+ sky130_fd_sc_hd__a22o_1
X_18871_ _18871_/A _25833_/Q _18871_/C vssd1 vssd1 vccd1 vccd1 _20797_/B sky130_fd_sc_hd__nand3_2
X_17822_ _18252_/A _21749_/A vssd1 vssd1 vccd1 vccd1 _17822_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
X_14965_ _14965_/A _14965_/B vssd1 vssd1 vccd1 vccd1 _14967_/A sky130_fd_sc_hd__nand2_1
X_17753_ _17753_/A _17757_/B vssd1 vssd1 vccd1 vccd1 _17874_/B sky130_fd_sc_hd__nor2b_1
X_16704_ _25861_/Q vssd1 vssd1 vccd1 vccd1 _21874_/B sky130_fd_sc_hd__inv_2
X_13916_ _13941_/A _13916_/B vssd1 vssd1 vccd1 vccd1 _13916_/Y sky130_fd_sc_hd__nand2_1
X_17684_ _17721_/B _17707_/B vssd1 vssd1 vccd1 vccd1 _17686_/A sky130_fd_sc_hd__nand2_1
X_14896_ _14896_/A vssd1 vssd1 vccd1 vccd1 _15083_/A sky130_fd_sc_hd__inv_2
XFILLER_0_18_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16635_ _16635_/A _16686_/B _16642_/A vssd1 vssd1 vccd1 vccd1 _16635_/Y sky130_fd_sc_hd__nand3_1
X_19423_ _19415_/X _19422_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19423_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13847_ _26273_/Q _13801_/X _13793_/X _13846_/Y vssd1 vssd1 vccd1 vccd1 _13848_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16566_ _16566_/A _16575_/A vssd1 vssd1 vccd1 vccd1 _16566_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_175_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19354_ _19352_/Y _19353_/Y _19086_/X vssd1 vssd1 vccd1 vccd1 _19354_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13778_ _13823_/A _13778_/B vssd1 vssd1 vccd1 vccd1 _13778_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_85_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15517_ _15505_/Y _15550_/A _15233_/X vssd1 vssd1 vccd1 vccd1 _15517_/Y sky130_fd_sc_hd__a21oi_1
X_18305_ _18305_/A _21844_/A _18305_/C vssd1 vssd1 vccd1 vccd1 _21109_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_85_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12729_ _14120_/A vssd1 vssd1 vccd1 vccd1 _13518_/B sky130_fd_sc_hd__buf_12
X_19285_ _26225_/Q _12537_/B hold419/X vssd1 vssd1 vccd1 vccd1 _19285_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16497_ hold745/X vssd1 vssd1 vccd1 vccd1 _16501_/B sky130_fd_sc_hd__inv_2
XFILLER_0_183_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18236_ _21022_/B _19430_/A vssd1 vssd1 vccd1 vccd1 _18237_/B sky130_fd_sc_hd__nand2_1
X_15448_ _15448_/A _23629_/B vssd1 vssd1 vccd1 vccd1 _15449_/A sky130_fd_sc_hd__and2_1
XFILLER_0_143_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18167_ _18445_/A _18172_/B vssd1 vssd1 vccd1 vccd1 _18170_/A sky130_fd_sc_hd__nand2_1
X_15379_ _15377_/X hold2399/X _15090_/X vssd1 vssd1 vccd1 vccd1 _25450_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17118_ _20362_/B _25886_/Q _25822_/Q vssd1 vssd1 vccd1 vccd1 _17119_/B sky130_fd_sc_hd__mux2_2
Xhold404 hold404/A vssd1 vssd1 vccd1 vccd1 hold404/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold415 hold415/A vssd1 vssd1 vccd1 vccd1 hold415/X sky130_fd_sc_hd__dlygate4sd3_1
X_18098_ _18098_/A vssd1 vssd1 vccd1 vccd1 _18954_/A sky130_fd_sc_hd__buf_12
Xhold426 hold426/A vssd1 vssd1 vccd1 vccd1 hold426/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold437 hold437/A vssd1 vssd1 vccd1 vccd1 hold437/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold448 hold448/A vssd1 vssd1 vccd1 vccd1 hold448/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17049_ _17047_/Y _17048_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _17049_/Y sky130_fd_sc_hd__a21oi_1
Xhold459 hold459/A vssd1 vssd1 vccd1 vccd1 hold459/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20060_ _20062_/C vssd1 vssd1 vccd1 vccd1 _20061_/B sky130_fd_sc_hd__inv_2
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 _12965_/X vssd1 vssd1 vccd1 vccd1 _25043_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1115 _25023_/Q vssd1 vssd1 vccd1 vccd1 _17309_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 _19919_/Y vssd1 vssd1 vccd1 vccd1 _25766_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1137 _25031_/Q vssd1 vssd1 vccd1 vccd1 _17393_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1148 _19499_/Y vssd1 vssd1 vccd1 vccd1 _25736_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 _25028_/Q vssd1 vssd1 vccd1 vccd1 _17363_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23750_ _23750_/A vssd1 vssd1 vccd1 vccd1 _25988_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20962_ _21235_/A _20962_/B vssd1 vssd1 vccd1 vccd1 _20962_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_178_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22701_ _23023_/A _23168_/B vssd1 vssd1 vccd1 vccd1 _22702_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23681_ hold1903/X _25966_/Q _23754_/S vssd1 vssd1 vccd1 vccd1 _23681_/X sky130_fd_sc_hd__mux2_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20893_ _21692_/A _21467_/B vssd1 vssd1 vccd1 vccd1 _20894_/B sky130_fd_sc_hd__nand2_1
X_25420_ _25420_/CLK _25420_/D vssd1 vssd1 vccd1 vccd1 _25420_/Q sky130_fd_sc_hd__dfxtp_1
X_22632_ _22631_/A _22454_/X _22631_/B vssd1 vssd1 vccd1 vccd1 _22633_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25351_ _26301_/CLK hold178/X vssd1 vssd1 vccd1 vccd1 hold176/A sky130_fd_sc_hd__dfxtp_1
X_22563_ _22563_/A _25895_/Q vssd1 vssd1 vccd1 vccd1 _22563_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_119_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24302_ hold2187/X hold2058/X _24356_/S vssd1 vssd1 vccd1 vccd1 _24303_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21514_ _21514_/A _21562_/A vssd1 vssd1 vccd1 vccd1 _21516_/A sky130_fd_sc_hd__nand2_1
X_25282_ _26235_/CLK hold256/X vssd1 vssd1 vccd1 vccd1 hold254/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22494_ _22494_/A _22494_/B vssd1 vssd1 vccd1 vccd1 _23040_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_118_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24233_ _24233_/A vssd1 vssd1 vccd1 vccd1 _26143_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21445_ _21443_/Y _21444_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21445_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_161_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24164_ _24164_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24165_/A sky130_fd_sc_hd__and2_1
X_21376_ _21375_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21376_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23115_ _23115_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _23115_/Y sky130_fd_sc_hd__nand2_1
X_20327_ _20330_/A _20330_/C vssd1 vssd1 vccd1 vccd1 _20329_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_141_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24095_ hold2267/X hold2218/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24096_/A sky130_fd_sc_hd__mux2_1
Xhold960 hold960/A vssd1 vssd1 vccd1 vccd1 hold960/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 hold971/A vssd1 vssd1 vccd1 vccd1 hold971/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold982 hold982/A vssd1 vssd1 vccd1 vccd1 hold982/X sky130_fd_sc_hd__dlygate4sd3_1
X_23046_ _26075_/Q vssd1 vssd1 vccd1 vccd1 _23047_/A sky130_fd_sc_hd__inv_2
Xhold993 hold993/A vssd1 vssd1 vccd1 vccd1 hold993/X sky130_fd_sc_hd__dlygate4sd3_1
X_20258_ _21466_/A _21114_/C vssd1 vssd1 vccd1 vccd1 _20261_/B sky130_fd_sc_hd__nand2_1
X_20189_ _20189_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20195_/A sky130_fd_sc_hd__nand2_2
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2350 _18622_/Y vssd1 vssd1 vccd1 vccd1 _25675_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2361 _23290_/A vssd1 vssd1 vccd1 vccd1 _23287_/C sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2372 _26284_/Q vssd1 vssd1 vccd1 vccd1 hold2372/X sky130_fd_sc_hd__buf_1
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24997_ _26046_/CLK _24997_/D vssd1 vssd1 vccd1 vccd1 _24997_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2383 _24114_/X vssd1 vssd1 vccd1 vccd1 _24115_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2394 _25663_/Q vssd1 vssd1 vccd1 vccd1 _13176_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1660 _21591_/Y vssd1 vssd1 vccd1 vccd1 _25829_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ _14900_/A _14750_/B vssd1 vssd1 vccd1 vccd1 _14750_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_118_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1671 _25600_/Q vssd1 vssd1 vccd1 vccd1 _17272_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23948_ _23948_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23949_/A sky130_fd_sc_hd__and2_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1682 _21624_/Y vssd1 vssd1 vccd1 vccd1 _25831_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1693 _19783_/Y vssd1 vssd1 vccd1 vccd1 _25756_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _18429_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13701_/Y sky130_fd_sc_hd__nor2_1
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _14681_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _14681_/Y sky130_fd_sc_hd__nand2_1
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23879_ _23879_/A vssd1 vssd1 vccd1 vccd1 _26030_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16420_ _16420_/A _16420_/B vssd1 vssd1 vccd1 vccd1 _16428_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_157_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25618_ _25619_/CLK _25618_/D vssd1 vssd1 vccd1 vccd1 _25618_/Q sky130_fd_sc_hd__dfxtp_2
X_13632_ _18202_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13632_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_39_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16351_ _16351_/A _16351_/B vssd1 vssd1 vccd1 vccd1 _16351_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25549_ _25875_/CLK _25549_/D vssd1 vssd1 vccd1 vccd1 _25549_/Q sky130_fd_sc_hd__dfxtp_1
X_13563_ _18034_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13563_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_41_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15302_ _15302_/A vssd1 vssd1 vccd1 vccd1 _16304_/A sky130_fd_sc_hd__inv_2
XFILLER_0_54_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12514_ _12514_/A _12514_/B _12514_/C _12514_/D vssd1 vssd1 vccd1 vccd1 _12515_/C
+ sky130_fd_sc_hd__or4_1
X_19070_ _19070_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _19070_/Y sky130_fd_sc_hd__nand2_1
X_16282_ _16676_/A _16282_/B vssd1 vssd1 vccd1 vccd1 _16285_/A sky130_fd_sc_hd__or2_1
X_13494_ _17974_/A _13518_/B vssd1 vssd1 vccd1 vccd1 _13494_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_70_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18021_ _18022_/B _18022_/A vssd1 vssd1 vccd1 vccd1 _20216_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15233_ _16231_/A vssd1 vssd1 vccd1 vccd1 _15233_/X sky130_fd_sc_hd__buf_12
XFILLER_0_87_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15164_ _15162_/A _15124_/B _15145_/A vssd1 vssd1 vccd1 vccd1 _15165_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14115_ _26316_/Q _13988_/X _13981_/X _14114_/Y vssd1 vssd1 vccd1 vccd1 _14116_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15095_ _22423_/B _15095_/B vssd1 vssd1 vccd1 vccd1 _22425_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19972_ _19972_/A _19972_/B vssd1 vssd1 vccd1 vccd1 _19972_/Y sky130_fd_sc_hd__nand2_1
X_14046_ _25802_/Q vssd1 vssd1 vccd1 vccd1 _18244_/B sky130_fd_sc_hd__inv_2
X_18923_ _18986_/A _19659_/A vssd1 vssd1 vccd1 vccd1 _18923_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_157_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18854_ _18854_/A _18854_/B _18854_/C vssd1 vssd1 vccd1 vccd1 _22592_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_158_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17805_ _22278_/B _25599_/Q vssd1 vssd1 vccd1 vccd1 _17807_/A sky130_fd_sc_hd__nand2_1
X_15997_ _16027_/A _15997_/B vssd1 vssd1 vccd1 vccd1 _16026_/A sky130_fd_sc_hd__nand2_1
X_18785_ _22513_/B _25637_/Q vssd1 vssd1 vccd1 vccd1 _18787_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_173_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14948_ _14948_/A _14948_/B vssd1 vssd1 vccd1 vccd1 _14950_/A sky130_fd_sc_hd__nand2_1
X_17736_ _17740_/B vssd1 vssd1 vccd1 vccd1 _17737_/B sky130_fd_sc_hd__inv_2
XFILLER_0_187_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14879_ _25858_/Q _12527_/A _15065_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14879_/X
+ sky130_fd_sc_hd__a22o_1
X_17667_ _17667_/A _19089_/A vssd1 vssd1 vccd1 vccd1 _19018_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_148_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19406_ _19407_/B _19407_/A vssd1 vssd1 vccd1 vccd1 _19406_/X sky130_fd_sc_hd__or2_1
X_16618_ _16618_/A _16618_/B vssd1 vssd1 vccd1 vccd1 _16629_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_159_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17598_ _17605_/A _17598_/B vssd1 vssd1 vccd1 vccd1 _17598_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_92_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16549_ _16551_/B _16551_/A vssd1 vssd1 vccd1 vccd1 _16550_/A sky130_fd_sc_hd__nor2_1
X_19337_ _19335_/X _19336_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19337_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19268_ _19452_/A _19268_/B vssd1 vssd1 vccd1 vccd1 _19268_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_183_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18219_ _18445_/A _18223_/B vssd1 vssd1 vccd1 vccd1 _18221_/A sky130_fd_sc_hd__nand2_1
X_19199_ _19199_/A vssd1 vssd1 vccd1 vccd1 _19452_/A sky130_fd_sc_hd__buf_8
XFILLER_0_131_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21230_ _26312_/Q hold569/X vssd1 vssd1 vccd1 vccd1 _21230_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_103_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold201 hold201/A vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 hold212/A vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 hold223/A vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21161_ _21164_/A _21164_/B vssd1 vssd1 vccd1 vccd1 _21163_/A sky130_fd_sc_hd__nand2_1
Xhold234 hold234/A vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 hold245/A vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 hold256/A vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 hold267/A vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold278 hold278/A vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
X_20112_ _19114_/A _21821_/A _25584_/Q vssd1 vssd1 vccd1 vccd1 _20113_/B sky130_fd_sc_hd__a21o_1
Xhold289 hold289/A vssd1 vssd1 vccd1 vccd1 hold289/X sky130_fd_sc_hd__dlygate4sd3_1
X_21092_ _26307_/Q _20731_/X hold796/X vssd1 vssd1 vccd1 vccd1 _21095_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_206_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _25594_/CLK sky130_fd_sc_hd__clkbuf_16
X_24920_ hold918/A hold962/A _24942_/S vssd1 vssd1 vccd1 vccd1 _24921_/B sky130_fd_sc_hd__mux2_1
X_20043_ _20043_/A _22692_/B vssd1 vssd1 vccd1 vccd1 _20044_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24851_ _24847_/X _24850_/X _25910_/Q vssd1 vssd1 vccd1 vccd1 _24851_/X sky130_fd_sc_hd__mux2_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23802_ _23802_/A vssd1 vssd1 vccd1 vccd1 _26005_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24782_ _24782_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24783_/A sky130_fd_sc_hd__and2_1
X_21994_ _21994_/A _21994_/B vssd1 vssd1 vccd1 vccd1 _23010_/A sky130_fd_sc_hd__xor2_4
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23733_ hold2244/X _14714_/B _23754_/S vssd1 vssd1 vccd1 vccd1 _23734_/A sky130_fd_sc_hd__mux2_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20945_ _20945_/A _20945_/B vssd1 vssd1 vccd1 vccd1 _21497_/C sky130_fd_sc_hd__nand2_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23664_ _23664_/A vssd1 vssd1 vccd1 vccd1 _25960_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20876_ _20875_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20876_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25403_ _25992_/CLK _25403_/D vssd1 vssd1 vccd1 vccd1 _25403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22615_ _25833_/Q _22615_/B vssd1 vssd1 vccd1 vccd1 _22615_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_119_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23595_ _23484_/Y hold1848/X _23593_/X _23594_/X vssd1 vssd1 vccd1 vccd1 _23595_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25334_ _26287_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22546_ _23072_/B vssd1 vssd1 vccd1 vccd1 _23071_/B sky130_fd_sc_hd__inv_2
XFILLER_0_119_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25265_ _26219_/CLK hold238/X vssd1 vssd1 vccd1 vccd1 hold236/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22477_ _15138_/B _22387_/B _14273_/X vssd1 vssd1 vccd1 vccd1 _22477_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24216_ hold2268/X hold2234/X _24279_/S vssd1 vssd1 vccd1 vccd1 _24217_/A sky130_fd_sc_hd__mux2_1
X_21428_ _21573_/A _21428_/B vssd1 vssd1 vccd1 vccd1 _21428_/Y sky130_fd_sc_hd__nand2_1
X_25196_ _26251_/CLK hold709/X vssd1 vssd1 vccd1 vccd1 hold707/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24147_ _24147_/A vssd1 vssd1 vccd1 vccd1 _26115_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21359_ _21358_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21359_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24078_ _24078_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24079_/A sky130_fd_sc_hd__and2_1
Xhold790 hold790/A vssd1 vssd1 vccd1 vccd1 hold790/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15920_ _15940_/A vssd1 vssd1 vccd1 vccd1 _15925_/B sky130_fd_sc_hd__inv_2
X_23029_ _15635_/B _22893_/A _22829_/X vssd1 vssd1 vccd1 vccd1 _23029_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15851_ _15849_/X hold507/X _15805_/X vssd1 vssd1 vccd1 vccd1 hold508/A sky130_fd_sc_hd__a21oi_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2180 _26051_/Q vssd1 vssd1 vccd1 vccd1 hold2180/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _25849_/Q _13466_/A _14801_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14803_/A
+ sky130_fd_sc_hd__a22o_1
Xhold2191 _12605_/Y vssd1 vssd1 vccd1 vccd1 _12606_/C sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15782_ _15787_/A _15762_/B _15760_/A vssd1 vssd1 vccd1 vccd1 _15783_/B sky130_fd_sc_hd__a21o_1
X_18570_ _18611_/A _25754_/Q vssd1 vssd1 vccd1 vccd1 _18572_/A sky130_fd_sc_hd__nand2_1
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12994_ _26132_/Q _12907_/X _12993_/X vssd1 vssd1 vccd1 vccd1 _12994_/X sky130_fd_sc_hd__a21o_1
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1490 _19769_/Y vssd1 vssd1 vccd1 vccd1 _25755_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14733_ _15839_/A _14733_/B vssd1 vssd1 vccd1 vccd1 _21865_/A sky130_fd_sc_hd__nand2_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17521_ _17624_/A _25047_/Q _17572_/C vssd1 vssd1 vccd1 vccd1 _17521_/X sky130_fd_sc_hd__and3_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _17452_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17452_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_86_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14664_ _14688_/A hold38/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__nand2_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16403_ _16403_/A vssd1 vssd1 vccd1 vccd1 _16416_/A sky130_fd_sc_hd__inv_2
XFILLER_0_131_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13615_ _26236_/Q _13612_/X _13605_/X _13614_/Y vssd1 vssd1 vccd1 vccd1 _13616_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17383_ _17393_/A _17383_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17383_/X sky130_fd_sc_hd__and3_1
XFILLER_0_39_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14595_ _14593_/Y hold387/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold388/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16334_ _16334_/A _16334_/B vssd1 vssd1 vccd1 vccd1 _16335_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_171_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19122_ _19121_/Y _21228_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19124_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_109_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13546_ _13583_/A _13546_/B vssd1 vssd1 vccd1 vccd1 _13546_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_109_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19053_ _19053_/A _19053_/B vssd1 vssd1 vccd1 vccd1 _19053_/X sky130_fd_sc_hd__xor2_1
X_16265_ _16269_/A _16265_/B vssd1 vssd1 vccd1 vccd1 _16266_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13477_ _26214_/Q _13426_/X _13468_/X _13476_/Y vssd1 vssd1 vccd1 vccd1 _13478_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_180_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15216_ _15188_/X _15268_/B _15199_/B vssd1 vssd1 vccd1 vccd1 _15218_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_124_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18004_ _20824_/B _21803_/A vssd1 vssd1 vccd1 vccd1 _20817_/A sky130_fd_sc_hd__nand2_2
X_16196_ _16208_/B _16196_/B vssd1 vssd1 vccd1 vccd1 _16197_/A sky130_fd_sc_hd__and2_1
XFILLER_0_65_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15147_ _15112_/X _15162_/B _15124_/B vssd1 vssd1 vccd1 vccd1 _15149_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_26_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15078_ _15073_/A _15066_/A _15066_/B vssd1 vssd1 vccd1 vccd1 _15080_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_26_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19955_ _26273_/Q hold780/X vssd1 vssd1 vccd1 vccd1 _19955_/Y sky130_fd_sc_hd__nand2_1
X_14029_ _26302_/Q _13988_/X _13981_/X _14028_/Y vssd1 vssd1 vccd1 vccd1 _14030_/B
+ sky130_fd_sc_hd__a22o_1
X_18906_ _25707_/Q vssd1 vssd1 vccd1 vccd1 _22665_/B sky130_fd_sc_hd__inv_2
X_19886_ _19959_/A _19901_/B vssd1 vssd1 vccd1 vccd1 _19888_/A sky130_fd_sc_hd__xnor2_1
X_18837_ _18988_/A _19038_/B vssd1 vssd1 vccd1 vccd1 _18838_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18768_ _25892_/Q _22487_/A vssd1 vssd1 vccd1 vccd1 _18776_/A sky130_fd_sc_hd__or2_2
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17719_ _17719_/A _17719_/B _23208_/B vssd1 vssd1 vccd1 vccd1 _17725_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_171_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18699_ _19026_/A _18699_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18699_/X sky130_fd_sc_hd__and3_1
XFILLER_0_78_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20730_ _20730_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20736_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20661_ _20659_/Y _20660_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _20661_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22400_ _22823_/B _22975_/B vssd1 vssd1 vccd1 vccd1 _22402_/C sky130_fd_sc_hd__nand2_1
X_23380_ _23380_/A hold476/X vssd1 vssd1 vccd1 vccd1 hold477/A sky130_fd_sc_hd__nand2_1
XFILLER_0_144_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20592_ _20592_/A _20592_/B vssd1 vssd1 vccd1 vccd1 _20594_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22331_ _22332_/B _22332_/A vssd1 vssd1 vccd1 vccd1 _22333_/A sky130_fd_sc_hd__or2_1
XFILLER_0_14_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25050_ _26135_/CLK _25050_/D vssd1 vssd1 vccd1 vccd1 _25050_/Q sky130_fd_sc_hd__dfxtp_1
X_22262_ _22653_/A _22262_/B vssd1 vssd1 vccd1 vccd1 _22262_/X sky130_fd_sc_hd__or2_1
XFILLER_0_143_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24001_ hold2437/X hold2449/X _24001_/S vssd1 vssd1 vccd1 vccd1 _24002_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21213_ _21213_/A _25873_/Q vssd1 vssd1 vccd1 vccd1 _21217_/B sky130_fd_sc_hd__nand2_1
X_22193_ _19230_/A _22192_/A _22192_/Y vssd1 vssd1 vccd1 vccd1 _22195_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21144_ _21144_/A _21144_/B _21144_/C vssd1 vssd1 vccd1 vccd1 _21145_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25952_ _26021_/CLK _25952_/D vssd1 vssd1 vccd1 vccd1 _25952_/Q sky130_fd_sc_hd__dfxtp_1
X_21075_ _21075_/A _21075_/B vssd1 vssd1 vccd1 vccd1 _21078_/B sky130_fd_sc_hd__nand2_1
X_24903_ _15918_/B _15932_/B _24945_/S vssd1 vssd1 vccd1 vccd1 _24903_/X sky130_fd_sc_hd__mux2_1
X_20026_ _20026_/A _20026_/B vssd1 vssd1 vccd1 vccd1 _20949_/C sky130_fd_sc_hd__xnor2_4
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25883_ _25883_/CLK _25883_/D vssd1 vssd1 vccd1 vccd1 _25883_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24834_ _24834_/A vssd1 vssd1 vccd1 vccd1 _26339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24765_ _24765_/A vssd1 vssd1 vccd1 vccd1 _26316_/D sky130_fd_sc_hd__clkbuf_1
X_21977_ _21977_/A _21977_/B vssd1 vssd1 vccd1 vccd1 _21978_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_68_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23716_ _23716_/A vssd1 vssd1 vccd1 vccd1 _25977_/D sky130_fd_sc_hd__clkbuf_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20928_ _26301_/Q hold635/X vssd1 vssd1 vccd1 vccd1 _20928_/Y sky130_fd_sc_hd__nand2_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24696_ _24696_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24697_/A sky130_fd_sc_hd__and2_1
XFILLER_0_68_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23647_ hold2086/X hold2068/X _23677_/S vssd1 vssd1 vccd1 vccd1 _23648_/A sky130_fd_sc_hd__mux2_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20859_ _25860_/Q vssd1 vssd1 vccd1 vccd1 _21840_/B sky130_fd_sc_hd__inv_2
X_13400_ _13315_/X _13398_/X _13300_/X _13399_/X vssd1 vssd1 vccd1 vccd1 _13400_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14380_ _14404_/A hold107/X vssd1 vssd1 vccd1 vccd1 hold108/A sky130_fd_sc_hd__nand2_1
X_23578_ _23566_/X _23577_/X _24949_/S vssd1 vssd1 vccd1 vccd1 _23578_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_187_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25317_ _26142_/CLK hold481/X vssd1 vssd1 vccd1 vccd1 hold479/A sky130_fd_sc_hd__dfxtp_1
X_13331_ _13220_/X _14620_/A _13242_/X _19616_/A vssd1 vssd1 vccd1 vccd1 _13331_/X
+ sky130_fd_sc_hd__a22o_1
X_22529_ _22529_/A _22529_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22531_/A sky130_fd_sc_hd__or3_1
XFILLER_0_36_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26297_ _26297_/CLK _26297_/D vssd1 vssd1 vccd1 vccd1 _26297_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_135_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16050_ _16071_/B _16050_/B vssd1 vssd1 vccd1 vccd1 _16084_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_122_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25248_ _25249_/CLK hold475/X vssd1 vssd1 vccd1 vccd1 hold473/A sky130_fd_sc_hd__dfxtp_1
X_13262_ _26179_/Q _13239_/X _13261_/X vssd1 vssd1 vccd1 vccd1 _13262_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_107_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15001_ _15033_/A _15032_/B _15032_/C _15000_/X vssd1 vssd1 vccd1 vccd1 _15003_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13193_ _18415_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13193_/X sky130_fd_sc_hd__or2_1
X_25179_ _25773_/CLK hold714/X vssd1 vssd1 vccd1 vccd1 hold713/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19740_ _26257_/Q _19134_/X hold584/X vssd1 vssd1 vccd1 vccd1 _19740_/Y sky130_fd_sc_hd__a21oi_1
X_16952_ _16953_/B _16953_/A vssd1 vssd1 vccd1 vccd1 _16952_/X sky130_fd_sc_hd__or2_1
X_15903_ _15901_/Y hold654/X _15805_/X vssd1 vssd1 vccd1 vccd1 hold655/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19671_ _19670_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19672_/B
+ sky130_fd_sc_hd__a211o_1
X_16883_ _16883_/A _16883_/B vssd1 vssd1 vccd1 vccd1 _16883_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18622_ _18620_/Y _18621_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _18622_/Y sky130_fd_sc_hd__a21oi_1
X_15834_ _15834_/A _15834_/B vssd1 vssd1 vccd1 vccd1 _15834_/Y sky130_fd_sc_hd__nand2_1
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ _18553_/A _20162_/A vssd1 vssd1 vccd1 vccd1 _18899_/A sky130_fd_sc_hd__xor2_4
X_15765_ _15764_/B _15731_/B _15746_/B vssd1 vssd1 vccd1 vccd1 _15765_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12977_ _12891_/X _14428_/A _12909_/X _25626_/Q vssd1 vssd1 vccd1 vccd1 _12977_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _17502_/Y _17503_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _25624_/D sky130_fd_sc_hd__a21oi_1
X_14716_ _21796_/B _15543_/B vssd1 vssd1 vccd1 vccd1 _14717_/A sky130_fd_sc_hd__nand2_1
X_15696_ _15675_/A _15657_/B _15674_/A vssd1 vssd1 vccd1 vccd1 _15696_/X sky130_fd_sc_hd__a21o_1
X_18484_ _25878_/Q _22119_/A vssd1 vssd1 vccd1 vccd1 _18492_/A sky130_fd_sc_hd__or2_2
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14647_ _14644_/Y hold153/X _14646_/X vssd1 vssd1 vccd1 vccd1 hold154/A sky130_fd_sc_hd__a21oi_1
X_17435_ _17624_/A _17435_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17435_/X sky130_fd_sc_hd__and3_1
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_18 _15384_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17366_ _17467_/A _17366_/B vssd1 vssd1 vccd1 vccd1 _17366_/Y sky130_fd_sc_hd__nand2_1
X_14578_ _14578_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14578_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_29 _19031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19105_ _20957_/A vssd1 vssd1 vccd1 vccd1 _19105_/X sky130_fd_sc_hd__buf_12
XFILLER_0_172_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16317_ _22731_/B _16369_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _16320_/B sky130_fd_sc_hd__and3_1
X_13529_ _14125_/A vssd1 vssd1 vccd1 vccd1 _13642_/A sky130_fd_sc_hd__clkbuf_8
X_17297_ _17295_/X _17241_/X _17296_/X vssd1 vssd1 vccd1 vccd1 _17298_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_125_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16248_ _16676_/A _16248_/B vssd1 vssd1 vccd1 vccd1 _16250_/A sky130_fd_sc_hd__or2_1
X_19036_ _19186_/A _19830_/A vssd1 vssd1 vccd1 vccd1 _19036_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16179_ _16179_/A hold860/X _16401_/C vssd1 vssd1 vccd1 vccd1 _16180_/B sky130_fd_sc_hd__and3_1
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19938_ _19990_/A _19939_/A vssd1 vssd1 vccd1 vccd1 _19938_/X sky130_fd_sc_hd__or2_1
XFILLER_0_177_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19869_ _26266_/Q _19134_/X hold617/X vssd1 vssd1 vccd1 vccd1 _19870_/C sky130_fd_sc_hd__a21o_1
X_21900_ _21900_/A _22145_/B vssd1 vssd1 vccd1 vccd1 _21900_/Y sky130_fd_sc_hd__nand2_1
X_22880_ _15474_/B _22680_/X _22829_/X vssd1 vssd1 vccd1 vccd1 _22880_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21831_ _21831_/A _22145_/B vssd1 vssd1 vccd1 vccd1 _21831_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24550_ hold2642/X _26247_/Q _24587_/S vssd1 vssd1 vccd1 vccd1 _24550_/X sky130_fd_sc_hd__mux2_1
X_21762_ _21762_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _21762_/X sky130_fd_sc_hd__and2_1
XFILLER_0_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23501_ _23498_/Y _23500_/Y _24858_/S vssd1 vssd1 vccd1 vccd1 _23501_/X sky130_fd_sc_hd__mux2_1
X_20713_ _20716_/A _20716_/C vssd1 vssd1 vccd1 vccd1 _20714_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_109_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24481_ _24481_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24482_/A sky130_fd_sc_hd__and2_1
XFILLER_0_92_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21693_ _21693_/A _21693_/B vssd1 vssd1 vccd1 vccd1 _21694_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_19_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26220_ _26221_/CLK _26220_/D vssd1 vssd1 vccd1 vccd1 _26220_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_11_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23432_ _23407_/X _23431_/X _25912_/Q vssd1 vssd1 vccd1 vccd1 _23432_/X sky130_fd_sc_hd__mux2_4
XFILLER_0_50_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20644_ _20644_/A _20644_/B vssd1 vssd1 vccd1 vccd1 _21629_/B sky130_fd_sc_hd__nand2_8
XFILLER_0_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26151_ _26151_/CLK _26151_/D vssd1 vssd1 vccd1 vccd1 _26151_/Q sky130_fd_sc_hd__dfxtp_1
X_23363_ _23363_/A vssd1 vssd1 vccd1 vccd1 _23366_/B sky130_fd_sc_hd__inv_2
XFILLER_0_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20575_ _20575_/A _20575_/B vssd1 vssd1 vccd1 vccd1 _20576_/A sky130_fd_sc_hd__nand2_1
X_25102_ _26317_/CLK _25102_/D vssd1 vssd1 vccd1 vccd1 _25102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22314_ _22314_/A _22314_/B vssd1 vssd1 vccd1 vccd1 _23039_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_108_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26082_ _26084_/CLK _26082_/D vssd1 vssd1 vccd1 vccd1 _26082_/Q sky130_fd_sc_hd__dfxtp_1
X_23294_ _23294_/A vssd1 vssd1 vccd1 vccd1 _23306_/A sky130_fd_sc_hd__inv_2
XFILLER_0_147_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25033_ _26117_/CLK _25033_/D vssd1 vssd1 vccd1 vccd1 _25033_/Q sky130_fd_sc_hd__dfxtp_1
X_22245_ _22245_/A _22875_/A vssd1 vssd1 vccd1 vccd1 _22257_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22176_ _22173_/X _15839_/B _22175_/Y _14831_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _22177_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_44_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21127_ _21125_/Y _21126_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21127_/Y sky130_fd_sc_hd__a21oi_1
X_25935_ _25938_/CLK _25935_/D vssd1 vssd1 vccd1 vccd1 _25935_/Q sky130_fd_sc_hd__dfxtp_1
X_21058_ _21516_/B _21564_/B vssd1 vssd1 vccd1 vccd1 _21059_/B sky130_fd_sc_hd__nand2_1
X_12900_ _17393_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12900_/X sky130_fd_sc_hd__or2_1
X_20009_ _21677_/A vssd1 vssd1 vccd1 vccd1 _21676_/A sky130_fd_sc_hd__inv_2
X_25866_ _25876_/CLK _25866_/D vssd1 vssd1 vccd1 vccd1 _25866_/Q sky130_fd_sc_hd__dfxtp_4
X_13880_ _13880_/A hold707/X vssd1 vssd1 vccd1 vccd1 hold708/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24817_ hold2695/X hold2561/X _24817_/S vssd1 vssd1 vccd1 vccd1 _24818_/A sky130_fd_sc_hd__mux2_1
X_12831_ _12726_/B _14337_/A _12752_/X _25598_/Q vssd1 vssd1 vccd1 vccd1 _12831_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25797_ _25797_/CLK _25797_/D vssd1 vssd1 vccd1 vccd1 _25797_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15550_ _15550_/A _15550_/B vssd1 vssd1 vccd1 vccd1 _15551_/A sky130_fd_sc_hd__nand2_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12762_ _12746_/X _12760_/X _14910_/B _12761_/X vssd1 vssd1 vccd1 vccd1 _12762_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24748_ hold2604/X _26311_/Q _24817_/S vssd1 vssd1 vccd1 vccd1 _24748_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_96_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14501_ _14525_/A hold134/X vssd1 vssd1 vccd1 vccd1 hold135/A sky130_fd_sc_hd__nand2_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _15481_/A _15481_/B vssd1 vssd1 vccd1 vccd1 _15502_/B sky130_fd_sc_hd__nor2_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12693_ _12693_/A vssd1 vssd1 vccd1 vccd1 _24990_/D sky130_fd_sc_hd__clkbuf_1
X_24679_ _24679_/A vssd1 vssd1 vccd1 vccd1 _26288_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _20856_/B _25860_/Q _20880_/B vssd1 vssd1 vccd1 vccd1 _17221_/B sky130_fd_sc_hd__mux2_2
X_14432_ _14465_/A hold170/X vssd1 vssd1 vccd1 vccd1 hold171/A sky130_fd_sc_hd__nand2_1
XFILLER_0_65_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17151_ _17272_/A _17151_/B vssd1 vssd1 vccd1 vccd1 _17151_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14363_ _14361_/Y hold51/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16102_ _16100_/X hold594/X _16076_/X vssd1 vssd1 vccd1 vccd1 hold595/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13314_ _13207_/X _13312_/X _13300_/X _13313_/X vssd1 vssd1 vccd1 vccd1 _13314_/X
+ sky130_fd_sc_hd__o211a_1
X_17082_ _25587_/Q vssd1 vssd1 vccd1 vccd1 _19176_/B sky130_fd_sc_hd__inv_2
XFILLER_0_126_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14294_ _14292_/Y hold156/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold157/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16033_ _16212_/A hold662/X vssd1 vssd1 vccd1 vccd1 hold663/A sky130_fd_sc_hd__nand2_1
X_13245_ _18577_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13245_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13176_ _13176_/A vssd1 vssd1 vccd1 vccd1 _19275_/A sky130_fd_sc_hd__buf_4
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17984_ _25852_/Q _22189_/A vssd1 vssd1 vccd1 vccd1 _17992_/A sky130_fd_sc_hd__or2_2
X_19723_ _19723_/A _19723_/B vssd1 vssd1 vccd1 vccd1 _19723_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_165_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16935_ _16935_/A _16940_/B vssd1 vssd1 vccd1 vccd1 _16937_/B sky130_fd_sc_hd__nand2_1
X_19654_ _19651_/Y _19652_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19654_/Y sky130_fd_sc_hd__a21oi_1
X_16866_ _16864_/Y _16865_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16866_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_189_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18605_ _20273_/B _19687_/A vssd1 vssd1 vccd1 vccd1 _18606_/B sky130_fd_sc_hd__nand2_1
X_15817_ _15817_/A _15817_/B vssd1 vssd1 vccd1 vccd1 _15830_/A sky130_fd_sc_hd__nor2_1
X_19585_ _26246_/Q hold545/X vssd1 vssd1 vccd1 vccd1 _19585_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_189_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16797_ _16795_/X _16711_/X _16796_/Y _25874_/Q _14170_/X vssd1 vssd1 vccd1 vccd1
+ _16798_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_181_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18536_ _18534_/X _18269_/X _18535_/X vssd1 vssd1 vccd1 vccd1 _18537_/A sky130_fd_sc_hd__a21o_1
X_15748_ _15720_/X _15764_/A _15731_/B vssd1 vssd1 vccd1 vccd1 _15750_/A sky130_fd_sc_hd__a21o_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18467_ _18467_/A _25813_/Q _18467_/C vssd1 vssd1 vccd1 vccd1 _20018_/C sky130_fd_sc_hd__nand3_2
X_15679_ _15677_/X hold2433/X _15464_/X vssd1 vssd1 vccd1 vccd1 _15679_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17418_ _17416_/Y _17417_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _17418_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18398_ _19546_/A vssd1 vssd1 vccd1 vccd1 _22015_/B sky130_fd_sc_hd__inv_2
XFILLER_0_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17349_ _21129_/B _25870_/Q _25806_/Q vssd1 vssd1 vccd1 vccd1 _17350_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_126_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20360_ _21195_/C vssd1 vssd1 vccd1 vccd1 _21198_/B sky130_fd_sc_hd__inv_2
XFILLER_0_31_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19019_ _19026_/A hold973/X _22786_/A vssd1 vssd1 vccd1 vccd1 _19019_/X sky130_fd_sc_hd__and3_1
XFILLER_0_114_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20291_ _20290_/B _20291_/B _20291_/C vssd1 vssd1 vccd1 vccd1 _20292_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22030_ _22030_/A _22030_/B _23026_/A vssd1 vssd1 vccd1 vccd1 _22030_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2702 _26339_/Q vssd1 vssd1 vccd1 vccd1 hold2702/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2713 _24805_/X vssd1 vssd1 vccd1 vccd1 _24806_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2724 _25909_/Q vssd1 vssd1 vccd1 vccd1 _23222_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2735 _26272_/Q vssd1 vssd1 vccd1 vccd1 hold2735/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2746 _26312_/Q vssd1 vssd1 vccd1 vccd1 hold2746/X sky130_fd_sc_hd__dlygate4sd3_1
X_23981_ _23981_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23982_/A sky130_fd_sc_hd__and2_1
Xhold2757 _25585_/Q vssd1 vssd1 vccd1 vccd1 hold2757/X sky130_fd_sc_hd__dlygate4sd3_1
X_25720_ _25783_/CLK _25720_/D vssd1 vssd1 vccd1 vccd1 _25720_/Q sky130_fd_sc_hd__dfxtp_1
X_22932_ _22931_/A _22849_/X _22931_/B vssd1 vssd1 vccd1 vccd1 _22933_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25651_ _26283_/CLK _25651_/D vssd1 vssd1 vccd1 vccd1 _25651_/Q sky130_fd_sc_hd__dfxtp_1
X_22863_ _23188_/A _22863_/B vssd1 vssd1 vccd1 vccd1 _22863_/X sky130_fd_sc_hd__or2_1
XFILLER_0_155_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24602_ _24602_/A vssd1 vssd1 vccd1 vccd1 _26263_/D sky130_fd_sc_hd__clkbuf_1
X_21814_ _22612_/B _21815_/A vssd1 vssd1 vccd1 vccd1 _21816_/A sky130_fd_sc_hd__or2_1
X_25582_ _25619_/CLK _25582_/D vssd1 vssd1 vccd1 vccd1 _25582_/Q sky130_fd_sc_hd__dfxtp_2
X_22794_ _22943_/A _22794_/B vssd1 vssd1 vccd1 vccd1 _22795_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24533_ _24533_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24534_/A sky130_fd_sc_hd__and2_1
X_21745_ _23055_/A _22550_/A vssd1 vssd1 vccd1 vccd1 _21754_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24464_ hold2690/X hold2584/X _24510_/S vssd1 vssd1 vccd1 vccd1 _24465_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21676_ _21676_/A _21676_/B vssd1 vssd1 vccd1 vccd1 _21678_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_175_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26203_ _26205_/CLK _26203_/D vssd1 vssd1 vccd1 vccd1 _26203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23415_ _24863_/S vssd1 vssd1 vccd1 vccd1 _24860_/S sky130_fd_sc_hd__buf_12
XFILLER_0_46_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20627_ _20627_/A _25854_/Q vssd1 vssd1 vccd1 vccd1 _20631_/B sky130_fd_sc_hd__nand2_1
X_24395_ _24395_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24396_/A sky130_fd_sc_hd__and2_1
XFILLER_0_61_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26134_ _26135_/CLK _26134_/D vssd1 vssd1 vccd1 vccd1 _26134_/Q sky130_fd_sc_hd__dfxtp_1
X_23346_ _23347_/B _23347_/A vssd1 vssd1 vccd1 vccd1 _23351_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_132_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20558_ _20558_/A _20558_/B vssd1 vssd1 vccd1 vccd1 _20562_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26065_ _26065_/CLK _26065_/D vssd1 vssd1 vccd1 vccd1 _26065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23277_ _23278_/A _23278_/B _23278_/C vssd1 vssd1 vccd1 vccd1 _23277_/X sky130_fd_sc_hd__a21o_1
X_20489_ _21276_/C _21563_/A vssd1 vssd1 vccd1 vccd1 _20492_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25016_ _26109_/CLK _25016_/D vssd1 vssd1 vccd1 vccd1 _25016_/Q sky130_fd_sc_hd__dfxtp_1
X_13030_ _12891_/X _14458_/A _12909_/X _25636_/Q vssd1 vssd1 vccd1 vccd1 _13030_/X
+ sky130_fd_sc_hd__a22o_1
X_22228_ _22226_/X _22227_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _22228_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_131_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22159_ _22159_/A _25851_/Q vssd1 vssd1 vccd1 vccd1 _22159_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14981_ _14981_/A _14981_/B vssd1 vssd1 vccd1 vccd1 _14998_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16720_ _16718_/X _16711_/X _16719_/Y _25863_/Q _14170_/X vssd1 vssd1 vccd1 vccd1
+ _16721_/A sky130_fd_sc_hd__a32o_1
X_25918_ _26341_/CLK _25918_/D vssd1 vssd1 vccd1 vccd1 _25918_/Q sky130_fd_sc_hd__dfxtp_1
X_13932_ _25784_/Q vssd1 vssd1 vccd1 vccd1 _17801_/B sky130_fd_sc_hd__inv_2
X_16651_ _16676_/A _16651_/B vssd1 vssd1 vccd1 vccd1 _16654_/A sky130_fd_sc_hd__nor2_1
X_13863_ _25773_/Q vssd1 vssd1 vccd1 vccd1 _18955_/B sky130_fd_sc_hd__inv_2
X_25849_ _26207_/CLK _25849_/D vssd1 vssd1 vccd1 vccd1 _25849_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15602_ _15602_/A vssd1 vssd1 vccd1 vccd1 _15604_/A sky130_fd_sc_hd__inv_2
X_12814_ _12726_/B _14328_/A _12752_/X _25595_/Q vssd1 vssd1 vccd1 vccd1 _12814_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19370_ _26231_/Q hold464/X vssd1 vssd1 vccd1 vccd1 _19370_/Y sky130_fd_sc_hd__nand2_1
X_16582_ _16698_/A hold918/X vssd1 vssd1 vccd1 vccd1 _16582_/Y sky130_fd_sc_hd__nand2_1
X_13794_ _25762_/Q vssd1 vssd1 vccd1 vccd1 _18733_/B sky130_fd_sc_hd__inv_2
XFILLER_0_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18321_ _18321_/A _18321_/B vssd1 vssd1 vccd1 vccd1 _21877_/A sky130_fd_sc_hd__nand2_1
X_15533_ _15505_/Y _15550_/A _15516_/B vssd1 vssd1 vccd1 vccd1 _15535_/A sky130_fd_sc_hd__a21o_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _12743_/X hold78/X _12558_/B vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15464_ _15464_/A vssd1 vssd1 vccd1 vccd1 _15464_/X sky130_fd_sc_hd__buf_6
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18252_ _18252_/A _18252_/B vssd1 vssd1 vccd1 vccd1 _18252_/Y sky130_fd_sc_hd__nand2_1
X_12676_ _12676_/A _12676_/B vssd1 vssd1 vccd1 vccd1 _12680_/A sky130_fd_sc_hd__nand2_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17203_ _17272_/A _17203_/B vssd1 vssd1 vccd1 vccd1 _17203_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_38_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14415_ _14413_/Y hold309/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold310/A sky130_fd_sc_hd__a21oi_1
X_15395_ _16827_/B vssd1 vssd1 vccd1 vccd1 _22815_/B sky130_fd_sc_hd__inv_2
X_18183_ _25655_/Q _20350_/B vssd1 vssd1 vccd1 vccd1 _18185_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_52_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14346_ _14343_/Y hold339/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold340/A sky130_fd_sc_hd__a21oi_1
X_17134_ _17413_/A _17134_/B vssd1 vssd1 vccd1 vccd1 _17134_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_25_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold608 hold608/A vssd1 vssd1 vccd1 vccd1 hold608/X sky130_fd_sc_hd__dlygate4sd3_1
X_17065_ _17063_/Y _17064_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _25585_/D sky130_fd_sc_hd__a21oi_1
X_14277_ _14277_/A _14277_/B _14277_/C vssd1 vssd1 vccd1 vccd1 _14279_/A sky130_fd_sc_hd__nor3_1
Xhold619 hold619/A vssd1 vssd1 vccd1 vccd1 hold619/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16016_ _16016_/A _16027_/B vssd1 vssd1 vccd1 vccd1 _16016_/Y sky130_fd_sc_hd__nand2_1
X_13228_ _26302_/Q _19388_/A vssd1 vssd1 vccd1 vccd1 _14569_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_21_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _26291_/Q _19230_/A vssd1 vssd1 vccd1 vccd1 _14536_/A sky130_fd_sc_hd__xor2_2
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2009 _23361_/X vssd1 vssd1 vccd1 vccd1 _23362_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1308 _25735_/Q vssd1 vssd1 vccd1 vccd1 _19481_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17967_ _17965_/Y _17966_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _25649_/D sky130_fd_sc_hd__a21oi_1
Xhold1319 _14760_/Y vssd1 vssd1 vccd1 vccd1 _25395_/D sky130_fd_sc_hd__dlygate4sd3_1
X_19706_ _19706_/A _19706_/B vssd1 vssd1 vccd1 vccd1 _19706_/Y sky130_fd_sc_hd__nand2_1
X_16918_ _16571_/B _16917_/Y _15621_/A vssd1 vssd1 vccd1 vccd1 _16918_/Y sky130_fd_sc_hd__a21oi_1
X_17898_ _17898_/A _20467_/A vssd1 vssd1 vccd1 vccd1 _19052_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_174_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19637_ _19629_/X _19636_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19637_/Y sky130_fd_sc_hd__o21ai_1
X_16849_ _16847_/X _16711_/X _16848_/Y _25882_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16850_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_137_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19568_ _19723_/A hold981/X vssd1 vssd1 vccd1 vccd1 _19568_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_48_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18519_ _18517_/Y _18518_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25670_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19499_ _19497_/Y _19498_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19499_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21530_ _21530_/A _21578_/A vssd1 vssd1 vccd1 vccd1 _21532_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21461_ _21459_/Y _21460_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21461_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23200_ _23200_/A vssd1 vssd1 vccd1 vccd1 _23212_/A sky130_fd_sc_hd__clkbuf_2
X_20412_ _21531_/A vssd1 vssd1 vccd1 vccd1 _21530_/A sky130_fd_sc_hd__inv_4
XFILLER_0_181_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24180_ _24180_/A vssd1 vssd1 vccd1 vccd1 _26126_/D sky130_fd_sc_hd__clkbuf_1
X_21392_ _21391_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21392_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23131_ _23131_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _23131_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20343_ _20342_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20343_/X
+ sky130_fd_sc_hd__a211o_1
X_23062_ _26076_/Q vssd1 vssd1 vccd1 vccd1 _23063_/A sky130_fd_sc_hd__inv_2
X_20274_ _20277_/A _20277_/C vssd1 vssd1 vccd1 vccd1 _20275_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22013_ _23184_/A vssd1 vssd1 vccd1 vccd1 _23183_/A sky130_fd_sc_hd__inv_2
XFILLER_0_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2510 _26059_/Q vssd1 vssd1 vccd1 vccd1 hold2510/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2521 _17691_/B vssd1 vssd1 vccd1 vccd1 _23205_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2532 _26317_/Q vssd1 vssd1 vccd1 vccd1 hold2532/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2543 _25680_/Q vssd1 vssd1 vccd1 vccd1 _13283_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2554 _25703_/Q vssd1 vssd1 vccd1 vccd1 _13427_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2565 _26221_/Q vssd1 vssd1 vccd1 vccd1 hold2565/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1820 _17525_/Y vssd1 vssd1 vccd1 vccd1 _25627_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1831 _26131_/Q vssd1 vssd1 vccd1 vccd1 hold1831/X sky130_fd_sc_hd__dlygate4sd3_1
X_23964_ _23964_/A vssd1 vssd1 vccd1 vccd1 _26056_/D sky130_fd_sc_hd__clkbuf_1
Xhold2576 _24587_/X vssd1 vssd1 vccd1 vccd1 _24588_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2587 _24615_/X vssd1 vssd1 vccd1 vccd1 _24616_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1842 _25709_/Q vssd1 vssd1 vccd1 vccd1 _19085_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1853 _22172_/Y vssd1 vssd1 vccd1 vccd1 _25851_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2598 _26158_/Q vssd1 vssd1 vccd1 vccd1 hold2598/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1864 _25633_/Q vssd1 vssd1 vccd1 vccd1 _17567_/B sky130_fd_sc_hd__dlygate4sd3_1
X_22915_ _22914_/A _22849_/X _22914_/B vssd1 vssd1 vccd1 vccd1 _22916_/C sky130_fd_sc_hd__o21ai_1
Xhold1875 _22261_/Y vssd1 vssd1 vccd1 vccd1 _25854_/D sky130_fd_sc_hd__dlygate4sd3_1
X_25703_ _26335_/CLK _25703_/D vssd1 vssd1 vccd1 vccd1 _25703_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1886 _14917_/A vssd1 vssd1 vccd1 vccd1 _14910_/C sky130_fd_sc_hd__dlygate4sd3_1
X_23895_ _26035_/Q hold2061/X _23907_/S vssd1 vssd1 vccd1 vccd1 _23895_/X sky130_fd_sc_hd__mux2_1
Xhold1897 _25706_/Q vssd1 vssd1 vccd1 vccd1 _19064_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22846_ _15435_/B _22680_/X _22829_/X vssd1 vssd1 vccd1 vccd1 _22846_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25634_ _26151_/CLK _25634_/D vssd1 vssd1 vccd1 vccd1 _25634_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25565_ _26069_/CLK _25565_/D vssd1 vssd1 vccd1 vccd1 _25565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22777_ _22926_/A _22777_/B vssd1 vssd1 vccd1 vccd1 _22778_/A sky130_fd_sc_hd__xor2_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12530_ _23245_/A vssd1 vssd1 vccd1 vccd1 _12558_/B sky130_fd_sc_hd__buf_12
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24516_ _24516_/A vssd1 vssd1 vccd1 vccd1 _26235_/D sky130_fd_sc_hd__clkbuf_1
X_21728_ _21728_/A _25857_/Q vssd1 vssd1 vccd1 vccd1 _21728_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_52_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25496_ _25919_/CLK hold430/X vssd1 vssd1 vccd1 vccd1 hold428/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24447_ _24447_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24448_/A sky130_fd_sc_hd__and2_1
XFILLER_0_19_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21659_ _21659_/A _21659_/B _21659_/C vssd1 vssd1 vccd1 vccd1 _21663_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_34_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14200_ _14236_/A hold783/X vssd1 vssd1 vccd1 vccd1 hold784/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15180_ _15166_/B _15184_/B _15161_/B vssd1 vssd1 vccd1 vccd1 _15180_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_105_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24378_ _24378_/A vssd1 vssd1 vccd1 vccd1 _26190_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26117_ _26117_/CLK _26117_/D vssd1 vssd1 vccd1 vccd1 _26117_/Q sky130_fd_sc_hd__dfxtp_1
X_14131_ hold758/X _14130_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold759/A sky130_fd_sc_hd__a21oi_1
X_23329_ _23336_/A vssd1 vssd1 vccd1 vccd1 _23334_/A sky130_fd_sc_hd__inv_2
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26048_ _26051_/CLK _26048_/D vssd1 vssd1 vccd1 vccd1 _26048_/Q sky130_fd_sc_hd__dfxtp_1
X_14062_ _14057_/Y _14061_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold797/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13013_ _26264_/Q _25633_/Q vssd1 vssd1 vccd1 vccd1 _14449_/A sky130_fd_sc_hd__xor2_2
X_18870_ _18952_/A _25769_/Q _18891_/C vssd1 vssd1 vccd1 vccd1 _18871_/C sky130_fd_sc_hd__nand3_1
X_17821_ _17821_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _17821_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_146_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17752_ _17830_/A _17752_/B vssd1 vssd1 vccd1 vccd1 _17757_/B sky130_fd_sc_hd__nand2_1
X_14964_ _14964_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14965_/B sky130_fd_sc_hd__nor2_1
X_16703_ _16976_/B vssd1 vssd1 vccd1 vccd1 _16857_/B sky130_fd_sc_hd__clkbuf_8
X_13915_ _26284_/Q _13801_/X _13793_/X _13914_/Y vssd1 vssd1 vccd1 vccd1 _13916_/B
+ sky130_fd_sc_hd__a22o_1
X_17683_ _17688_/A _17683_/B vssd1 vssd1 vccd1 vccd1 _17750_/B sky130_fd_sc_hd__nand2_2
X_14895_ _22386_/B _15543_/B vssd1 vssd1 vccd1 vccd1 _14896_/A sky130_fd_sc_hd__nand2_1
X_19422_ _19420_/X _19421_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19422_/Y sky130_fd_sc_hd__a21oi_1
X_16634_ _16634_/A _16647_/A vssd1 vssd1 vccd1 vccd1 _16642_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13846_ _18894_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13846_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_186_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19353_ _19452_/A _19353_/B vssd1 vssd1 vccd1 vccd1 _19353_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16565_ _16575_/A _16566_/A vssd1 vssd1 vccd1 vccd1 _16565_/X sky130_fd_sc_hd__or2_1
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13777_ _26262_/Q _13612_/X _13605_/X _13776_/Y vssd1 vssd1 vccd1 vccd1 _13778_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18304_ _18446_/A hold981/X _18952_/C vssd1 vssd1 vccd1 vccd1 _18305_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_73_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15516_ _15516_/A _15516_/B vssd1 vssd1 vccd1 vccd1 _15550_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_73_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12728_ _16774_/B vssd1 vssd1 vccd1 vccd1 _14120_/A sky130_fd_sc_hd__inv_8
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19284_ _19282_/Y _19283_/Y _19086_/X vssd1 vssd1 vccd1 vccd1 _19284_/Y sky130_fd_sc_hd__a21oi_1
X_16496_ _16599_/A vssd1 vssd1 vccd1 vccd1 _16503_/B sky130_fd_sc_hd__inv_2
XFILLER_0_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18235_ _21738_/B _25610_/Q vssd1 vssd1 vccd1 vccd1 _18237_/A sky130_fd_sc_hd__nand2_1
X_15447_ _15466_/B _15447_/B vssd1 vssd1 vccd1 vccd1 _15448_/A sky130_fd_sc_hd__xor2_1
X_12659_ _12659_/A vssd1 vssd1 vccd1 vccd1 _12664_/A sky130_fd_sc_hd__inv_2
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18166_ _25863_/Q _21937_/A vssd1 vssd1 vccd1 vccd1 _18175_/A sky130_fd_sc_hd__or2_2
X_15378_ _15378_/A _15405_/B vssd1 vssd1 vccd1 vccd1 _15378_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_25_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17117_ _25630_/Q vssd1 vssd1 vccd1 vccd1 _20362_/B sky130_fd_sc_hd__inv_2
XFILLER_0_25_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14329_ _14344_/A hold206/X vssd1 vssd1 vccd1 vccd1 hold207/A sky130_fd_sc_hd__nand2_1
Xhold405 hold405/A vssd1 vssd1 vccd1 vccd1 hold405/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18097_ _18097_/A _25797_/Q _18097_/C vssd1 vssd1 vccd1 vccd1 _20888_/B sky130_fd_sc_hd__nand3_2
Xhold416 hold416/A vssd1 vssd1 vccd1 vccd1 hold416/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 hold427/A vssd1 vssd1 vccd1 vccd1 hold427/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold438 hold438/A vssd1 vssd1 vccd1 vccd1 hold438/X sky130_fd_sc_hd__dlygate4sd3_1
X_17048_ _17272_/A _17048_/B vssd1 vssd1 vccd1 vccd1 _17048_/Y sky130_fd_sc_hd__nand2_1
Xhold449 hold449/A vssd1 vssd1 vccd1 vccd1 hold449/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1105 _25542_/Q vssd1 vssd1 vccd1 vccd1 _16722_/B sky130_fd_sc_hd__buf_1
X_18999_ _18997_/X _18879_/X _18998_/X vssd1 vssd1 vccd1 vccd1 _19000_/A sky130_fd_sc_hd__a21o_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1116 _12860_/X vssd1 vssd1 vccd1 vccd1 _25023_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1127 _25489_/Q vssd1 vssd1 vccd1 vccd1 _16018_/B sky130_fd_sc_hd__buf_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1138 _12901_/X vssd1 vssd1 vccd1 vccd1 _25031_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 _25080_/Q vssd1 vssd1 vccd1 vccd1 _18313_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20961_ _20961_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _20961_/Y sky130_fd_sc_hd__nand2_1
X_22700_ _23167_/B _23024_/B vssd1 vssd1 vccd1 vccd1 _22702_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23680_ _23920_/S vssd1 vssd1 vccd1 vccd1 _23754_/S sky130_fd_sc_hd__buf_12
XFILLER_0_45_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20892_ _21464_/C _21693_/A vssd1 vssd1 vccd1 vccd1 _20894_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22631_ _22631_/A _22631_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22633_/A sky130_fd_sc_hd__or3_1
XFILLER_0_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25350_ _26301_/CLK hold121/X vssd1 vssd1 vccd1 vccd1 hold119/A sky130_fd_sc_hd__dfxtp_1
X_22562_ _22560_/X _22561_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22562_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24301_ _24301_/A vssd1 vssd1 vccd1 vccd1 _26165_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21513_ _21513_/A _21513_/B _21513_/C vssd1 vssd1 vccd1 vccd1 _21517_/A sky130_fd_sc_hd__nand3_1
X_25281_ _26235_/CLK hold292/X vssd1 vssd1 vccd1 vccd1 hold290/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22493_ _22493_/A _22493_/B vssd1 vssd1 vccd1 vccd1 _22494_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_133_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24232_ _24232_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24233_/A sky130_fd_sc_hd__and2_1
XFILLER_0_106_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21444_ _21573_/A _21444_/B vssd1 vssd1 vccd1 vccd1 _21444_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_185_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24163_ hold2233/X hold2046/X _24203_/S vssd1 vssd1 vccd1 vccd1 _24164_/A sky130_fd_sc_hd__mux2_1
X_21375_ _26319_/Q hold731/X vssd1 vssd1 vccd1 vccd1 _21375_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23114_ _16949_/B _22421_/A _23108_/X _23109_/Y _23113_/X vssd1 vssd1 vccd1 vccd1
+ _23115_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20326_ _20326_/A _22332_/B _20326_/C vssd1 vssd1 vccd1 vccd1 _20330_/C sky130_fd_sc_hd__nand3_1
X_24094_ _24094_/A vssd1 vssd1 vccd1 vccd1 _26098_/D sky130_fd_sc_hd__clkbuf_1
Xhold950 hold950/A vssd1 vssd1 vccd1 vccd1 hold950/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold961 hold961/A vssd1 vssd1 vccd1 vccd1 hold961/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold972 hold972/A vssd1 vssd1 vccd1 vccd1 hold972/X sky130_fd_sc_hd__dlygate4sd3_1
X_23045_ _15650_/B _22893_/A _22829_/X vssd1 vssd1 vccd1 vccd1 _23045_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold983 hold983/A vssd1 vssd1 vccd1 vccd1 hold983/X sky130_fd_sc_hd__dlygate4sd3_1
X_20257_ _21465_/A _21117_/B vssd1 vssd1 vccd1 vccd1 _20261_/A sky130_fd_sc_hd__nand2_1
Xhold994 hold994/A vssd1 vssd1 vccd1 vccd1 hold994/X sky130_fd_sc_hd__dlygate4sd3_1
X_20188_ _20188_/A _20188_/B vssd1 vssd1 vccd1 vccd1 _20189_/A sky130_fd_sc_hd__nand2_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2340 _26123_/Q vssd1 vssd1 vccd1 vccd1 hold2340/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2351 _26102_/Q vssd1 vssd1 vccd1 vccd1 hold2351/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2362 _26170_/Q vssd1 vssd1 vccd1 vccd1 hold2362/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2373 _24668_/X vssd1 vssd1 vccd1 vccd1 _24669_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24996_ _26004_/CLK _24996_/D vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dfxtp_1
Xhold2384 _26172_/Q vssd1 vssd1 vccd1 vccd1 hold2384/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1650 _17139_/Y vssd1 vssd1 vccd1 vccd1 _25590_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2395 _25435_/Q vssd1 vssd1 vccd1 vccd1 _15092_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1661 _25875_/Q vssd1 vssd1 vccd1 vccd1 _22772_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23947_ hold2401/X hold2180/X _24001_/S vssd1 vssd1 vccd1 vccd1 _23948_/A sky130_fd_sc_hd__mux2_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1672 _17273_/Y vssd1 vssd1 vccd1 vccd1 _25600_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1683 _25878_/Q vssd1 vssd1 vccd1 vccd1 _22821_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1694 _25715_/Q vssd1 vssd1 vccd1 vccd1 _19200_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _25747_/Q vssd1 vssd1 vccd1 vccd1 _18429_/B sky130_fd_sc_hd__inv_2
XFILLER_0_86_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ _14678_/Y hold351/X _14646_/X vssd1 vssd1 vccd1 vccd1 hold352/A sky130_fd_sc_hd__a21oi_1
X_23878_ _23878_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23879_/A sky130_fd_sc_hd__and2_1
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13631_ _25736_/Q vssd1 vssd1 vccd1 vccd1 _18202_/B sky130_fd_sc_hd__inv_2
XFILLER_0_169_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22829_ _22829_/A vssd1 vssd1 vccd1 vccd1 _22829_/X sky130_fd_sc_hd__clkbuf_8
X_25617_ _25619_/CLK _25617_/D vssd1 vssd1 vccd1 vccd1 _25617_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_79_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16350_ _16351_/B _16351_/A vssd1 vssd1 vccd1 vccd1 _16350_/X sky130_fd_sc_hd__or2_1
X_13562_ _25725_/Q vssd1 vssd1 vccd1 vccd1 _18034_/B sky130_fd_sc_hd__inv_2
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25548_ _25875_/CLK _25548_/D vssd1 vssd1 vccd1 vccd1 _25548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12513_ _24987_/Q _24986_/Q _24985_/Q _24984_/Q vssd1 vssd1 vccd1 vccd1 _12514_/D
+ sky130_fd_sc_hd__or4_1
X_15301_ _22706_/B _15812_/B vssd1 vssd1 vccd1 vccd1 _15302_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_125_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16281_ hold701/X vssd1 vssd1 vccd1 vccd1 _16285_/B sky130_fd_sc_hd__inv_2
X_25479_ _25483_/CLK hold463/X vssd1 vssd1 vccd1 vccd1 hold461/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13493_ hold818/A vssd1 vssd1 vccd1 vccd1 _17974_/A sky130_fd_sc_hd__inv_2
XFILLER_0_54_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_160_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _26167_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18020_ _25715_/Q _18020_/B vssd1 vssd1 vccd1 vccd1 _18022_/A sky130_fd_sc_hd__xor2_2
X_15232_ _15232_/A _15232_/B vssd1 vssd1 vccd1 vccd1 _15266_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15163_ _15185_/A _15112_/X vssd1 vssd1 vccd1 vccd1 _15165_/A sky130_fd_sc_hd__or2b_1
XFILLER_0_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14114_ _18470_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14114_/Y sky130_fd_sc_hd__nor2_1
X_15094_ _26004_/Q _15809_/S _15774_/B vssd1 vssd1 vccd1 vccd1 _15095_/B sky130_fd_sc_hd__o21ai_4
X_19971_ _19972_/B _19972_/A vssd1 vssd1 vccd1 vccd1 _19971_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14045_ _14118_/A hold482/X vssd1 vssd1 vccd1 vccd1 hold483/A sky130_fd_sc_hd__nand2_1
X_18922_ _18922_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18922_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18853_ _18955_/A _18853_/B _18894_/C vssd1 vssd1 vccd1 vccd1 _18854_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_101_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17804_ _19275_/A vssd1 vssd1 vccd1 vccd1 _22278_/B sky130_fd_sc_hd__inv_2
X_18784_ _19816_/A vssd1 vssd1 vccd1 vccd1 _22513_/B sky130_fd_sc_hd__inv_2
X_15996_ _15996_/A _15996_/B vssd1 vssd1 vccd1 vccd1 _15997_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17735_ _17771_/C _17735_/B vssd1 vssd1 vccd1 vccd1 _17740_/B sky130_fd_sc_hd__nand2_1
X_14947_ _14947_/A _14947_/B vssd1 vssd1 vccd1 vccd1 _14948_/B sky130_fd_sc_hd__nor2_1
X_17666_ _20026_/A _17666_/B vssd1 vssd1 vccd1 vccd1 _19089_/A sky130_fd_sc_hd__nand2_2
X_14878_ _14878_/A vssd1 vssd1 vccd1 vccd1 _15065_/A sky130_fd_sc_hd__inv_2
XFILLER_0_159_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19405_ _19421_/B _19493_/B vssd1 vssd1 vccd1 vccd1 _19407_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16617_ _16617_/A hold887/X _16691_/B vssd1 vssd1 vccd1 vccd1 _16618_/B sky130_fd_sc_hd__and3_1
XFILLER_0_147_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13829_ _26270_/Q _13801_/X _13793_/X _13828_/Y vssd1 vssd1 vccd1 vccd1 _13830_/B
+ sky130_fd_sc_hd__a22o_1
X_17597_ _17597_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _17597_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19336_ _19336_/A _19336_/B vssd1 vssd1 vccd1 vccd1 _19336_/Y sky130_fd_sc_hd__nand2_1
X_16548_ _16676_/A _16548_/B vssd1 vssd1 vccd1 vccd1 _16551_/A sky130_fd_sc_hd__or2_1
X_19267_ _19267_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _19267_/Y sky130_fd_sc_hd__nand2_1
X_16479_ _16479_/A _16479_/B vssd1 vssd1 vccd1 vccd1 _16485_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_151_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _26175_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18218_ _25865_/Q _22005_/A vssd1 vssd1 vccd1 vccd1 _18226_/A sky130_fd_sc_hd__or2_2
XFILLER_0_26_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19198_ _19198_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _19198_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18149_ _25654_/Q _20310_/B vssd1 vssd1 vccd1 vccd1 _18151_/B sky130_fd_sc_hd__nor2_1
Xhold202 hold202/A vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 hold213/A vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold224 hold224/A vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21160_ _25871_/Q _21160_/B _21160_/C vssd1 vssd1 vccd1 vccd1 _21164_/B sky130_fd_sc_hd__nand3b_1
Xhold235 hold235/A vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold246 hold246/A vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 hold257/A vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold268 hold268/A vssd1 vssd1 vccd1 vccd1 hold268/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20111_ _20111_/A vssd1 vssd1 vccd1 vccd1 _20115_/A sky130_fd_sc_hd__inv_2
XFILLER_0_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold279 hold279/A vssd1 vssd1 vccd1 vccd1 hold279/X sky130_fd_sc_hd__dlygate4sd3_1
X_21091_ _21091_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _21096_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_102_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20042_ _20040_/Y _20041_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _20042_/Y sky130_fd_sc_hd__a21oi_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24850_ _24848_/X _24849_/X _24946_/A vssd1 vssd1 vccd1 vccd1 _24850_/X sky130_fd_sc_hd__mux2_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23801_ _23801_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23802_/A sky130_fd_sc_hd__and2_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24781_ hold2655/X _26322_/Q _24817_/S vssd1 vssd1 vccd1 vccd1 _24781_/X sky130_fd_sc_hd__mux2_1
X_21993_ _18124_/B _17125_/B _18126_/A vssd1 vssd1 vccd1 vccd1 _21994_/B sky130_fd_sc_hd__o21ai_2
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23732_ _23732_/A vssd1 vssd1 vccd1 vccd1 _25982_/D sky130_fd_sc_hd__clkbuf_1
X_20944_ _20944_/A _20944_/B _20944_/C vssd1 vssd1 vccd1 vccd1 _20945_/B sky130_fd_sc_hd__nand3_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23663_ _23663_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23664_/A sky130_fd_sc_hd__and2_1
XFILLER_0_113_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20875_ _26299_/Q hold578/X vssd1 vssd1 vccd1 vccd1 _20875_/Y sky130_fd_sc_hd__nand2_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25402_ _25425_/CLK _25402_/D vssd1 vssd1 vccd1 vccd1 _25402_/Q sky130_fd_sc_hd__dfxtp_1
X_22614_ _22614_/A _25897_/Q vssd1 vssd1 vccd1 vccd1 _22614_/Y sky130_fd_sc_hd__nand2_1
X_23594_ _23593_/X output9/A vssd1 vssd1 vccd1 vccd1 _23594_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_64_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25333_ _25796_/CLK hold181/X vssd1 vssd1 vccd1 vccd1 hold179/A sky130_fd_sc_hd__dfxtp_1
X_22545_ _22545_/A _22545_/B vssd1 vssd1 vccd1 vccd1 _23072_/B sky130_fd_sc_hd__nand2_4
Xclkbuf_leaf_142_clk clkbuf_4_11__f_clk/X vssd1 vssd1 vccd1 vccd1 _25678_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_187_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25264_ _26089_/CLK hold184/X vssd1 vssd1 vccd1 vccd1 hold182/A sky130_fd_sc_hd__dfxtp_1
X_22476_ _22653_/A _22476_/B vssd1 vssd1 vccd1 vccd1 _22476_/X sky130_fd_sc_hd__or2_1
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24215_ _24215_/A vssd1 vssd1 vccd1 vccd1 _26137_/D sky130_fd_sc_hd__clkbuf_1
X_21427_ _21427_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21427_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_115_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25195_ _26251_/CLK hold604/X vssd1 vssd1 vccd1 vccd1 hold602/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24146_ _24146_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24147_/A sky130_fd_sc_hd__and2_1
X_21358_ _26318_/Q hold757/X vssd1 vssd1 vccd1 vccd1 _21358_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20309_ _20309_/A _22026_/A vssd1 vssd1 vccd1 vccd1 _20310_/A sky130_fd_sc_hd__nand2_1
X_24077_ hold2255/X hold1/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24078_/A sky130_fd_sc_hd__mux2_1
X_21289_ _21287_/Y _21288_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21289_/Y sky130_fd_sc_hd__a21oi_1
Xhold780 hold780/A vssd1 vssd1 vccd1 vccd1 hold780/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold791 hold791/A vssd1 vssd1 vccd1 vccd1 hold791/X sky130_fd_sc_hd__dlygate4sd3_1
X_23028_ _23188_/A _23028_/B vssd1 vssd1 vccd1 vccd1 _23028_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15850_ _15956_/A hold506/X vssd1 vssd1 vccd1 vccd1 hold507/A sky130_fd_sc_hd__nand2_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2170 _23348_/X vssd1 vssd1 vccd1 vccd1 _23349_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2181 _23950_/X vssd1 vssd1 vccd1 vccd1 _23951_/A sky130_fd_sc_hd__dlygate4sd3_1
X_14801_ _25849_/Q _12527_/A _14989_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14801_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2192 _12606_/X vssd1 vssd1 vccd1 vccd1 _12607_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _15781_/A _15781_/B vssd1 vssd1 vccd1 vccd1 _15786_/A sky130_fd_sc_hd__nand2_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24979_ _24983_/CLK _24979_/D vssd1 vssd1 vccd1 vccd1 _24979_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _12891_/X _14437_/A _12909_/X _25629_/Q vssd1 vssd1 vccd1 vccd1 _12993_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17520_ _17520_/A _17520_/B vssd1 vssd1 vccd1 vccd1 _17520_/X sky130_fd_sc_hd__xor2_2
Xhold1480 _13012_/X vssd1 vssd1 vccd1 vccd1 _25052_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ _14730_/Y _14731_/Y _14646_/X vssd1 vssd1 vccd1 vccd1 _14732_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1491 _25815_/Q vssd1 vssd1 vccd1 vccd1 _21363_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _21791_/A vssd1 vssd1 vccd1 vccd1 _17582_/B sky130_fd_sc_hd__buf_6
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14663_ _14663_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _14663_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_170_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16402_ _16402_/A _16402_/B vssd1 vssd1 vccd1 vccd1 _16403_/A sky130_fd_sc_hd__nor2_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13614_ _18101_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13614_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_131_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17382_ _17645_/A _17382_/B vssd1 vssd1 vccd1 vccd1 _17382_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_95_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14594_ _14645_/A hold386/X vssd1 vssd1 vccd1 vccd1 hold387/A sky130_fd_sc_hd__nand2_1
XFILLER_0_184_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19121_ _26214_/Q hold497/X vssd1 vssd1 vccd1 vccd1 _19121_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_109_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16333_ _16333_/A _16336_/B vssd1 vssd1 vccd1 vccd1 _16334_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13545_ _26225_/Q _13426_/X _13468_/X _13544_/Y vssd1 vssd1 vccd1 vccd1 _13546_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_133_clk clkbuf_leaf_82_clk/A vssd1 vssd1 vccd1 vccd1 _25257_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_125_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19052_ _19052_/A _19052_/B vssd1 vssd1 vccd1 vccd1 _19053_/B sky130_fd_sc_hd__xnor2_1
X_16264_ _16264_/A _16264_/B vssd1 vssd1 vccd1 vccd1 _16265_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_180_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13476_ _17832_/A _13518_/B vssd1 vssd1 vccd1 vccd1 _13476_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_109_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18003_ _18003_/A _18003_/B _18003_/C vssd1 vssd1 vccd1 vccd1 _21803_/A sky130_fd_sc_hd__nand3_2
X_15215_ _15268_/C vssd1 vssd1 vccd1 vccd1 _15218_/B sky130_fd_sc_hd__inv_2
X_16195_ _16195_/A _16195_/B vssd1 vssd1 vccd1 vccd1 _16196_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_129_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15146_ _15162_/A vssd1 vssd1 vccd1 vccd1 _15149_/B sky130_fd_sc_hd__inv_2
XFILLER_0_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15077_ _15077_/A _15077_/B vssd1 vssd1 vccd1 vccd1 _15085_/B sky130_fd_sc_hd__nand2_1
X_19954_ _19952_/Y _19953_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _19954_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14028_ _18173_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14028_/Y sky130_fd_sc_hd__nor2_1
X_18905_ _25707_/Q _20000_/B vssd1 vssd1 vccd1 vccd1 _18908_/A sky130_fd_sc_hd__nor2_1
X_19885_ _20828_/A _18888_/A _20833_/C vssd1 vssd1 vccd1 vccd1 _19959_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_184_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18836_ _18836_/A _20711_/A vssd1 vssd1 vccd1 vccd1 _19038_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_101_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18767_ _18767_/A _18767_/B vssd1 vssd1 vccd1 vccd1 _22487_/A sky130_fd_sc_hd__nand2_1
X_15979_ _15979_/A _16697_/B _15987_/A vssd1 vssd1 vccd1 vccd1 _15979_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_89_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17718_ _17764_/A _17722_/A vssd1 vssd1 vccd1 vccd1 _17725_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18698_ _18698_/A _18698_/B vssd1 vssd1 vccd1 vccd1 _18698_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_187_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17649_ _18252_/A _17649_/B vssd1 vssd1 vccd1 vccd1 _17649_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_33_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20660_ _20660_/A _20660_/B vssd1 vssd1 vccd1 vccd1 _20660_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19319_ _20779_/A _19317_/Y _20784_/C vssd1 vssd1 vccd1 vccd1 _19407_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_124_clk clkbuf_4_14__f_clk/X vssd1 vssd1 vccd1 vccd1 _26324_/CLK sky130_fd_sc_hd__clkbuf_16
X_20591_ _20593_/B _20593_/C vssd1 vssd1 vccd1 vccd1 _20592_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22330_ _19701_/A _22329_/A _22329_/Y vssd1 vssd1 vccd1 vccd1 _22332_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22261_ _22259_/Y _22260_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _22261_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24000_ _24000_/A vssd1 vssd1 vccd1 vccd1 _26068_/D sky130_fd_sc_hd__clkbuf_1
X_21212_ _21214_/B _21214_/C vssd1 vssd1 vccd1 vccd1 _21213_/A sky130_fd_sc_hd__nand2_1
X_22192_ _22192_/A _22192_/B vssd1 vssd1 vccd1 vccd1 _22192_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_130_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21143_ _21564_/B _21610_/C vssd1 vssd1 vccd1 vccd1 _21144_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25951_ _26021_/CLK _25951_/D vssd1 vssd1 vccd1 vccd1 _25951_/Q sky130_fd_sc_hd__dfxtp_1
X_21074_ _21074_/A _21810_/B vssd1 vssd1 vccd1 vccd1 _21075_/A sky130_fd_sc_hd__nand2_1
X_24902_ _24900_/X _24901_/X _24957_/S vssd1 vssd1 vccd1 vccd1 _24902_/X sky130_fd_sc_hd__mux2_1
X_20025_ _20025_/A _20025_/B vssd1 vssd1 vccd1 vccd1 _20026_/B sky130_fd_sc_hd__xor2_2
X_25882_ _25901_/CLK _25882_/D vssd1 vssd1 vccd1 vccd1 _25882_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24833_ _24833_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24834_/A sky130_fd_sc_hd__and2_1
XFILLER_0_77_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21976_ _21977_/B _21977_/A vssd1 vssd1 vccd1 vccd1 _21978_/A sky130_fd_sc_hd__or2_1
XFILLER_0_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24764_ _24764_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24765_/A sky130_fd_sc_hd__and2_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23715_ _23715_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23716_/A sky130_fd_sc_hd__and2_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20927_ _26301_/Q _20731_/X hold635/X vssd1 vssd1 vccd1 vccd1 _20930_/B sky130_fd_sc_hd__a21oi_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24695_ hold2638/X hold2613/X _24740_/S vssd1 vssd1 vccd1 vccd1 _24696_/A sky130_fd_sc_hd__mux2_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23646_ _23646_/A vssd1 vssd1 vccd1 vccd1 _25954_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20858_ _20858_/A _25860_/Q vssd1 vssd1 vccd1 vccd1 _20863_/B sky130_fd_sc_hd__nand2_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_115_clk clkbuf_4_14__f_clk/X vssd1 vssd1 vccd1 vccd1 _26205_/CLK sky130_fd_sc_hd__clkbuf_16
X_23577_ _23571_/X _23576_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _23577_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20789_ _21419_/B vssd1 vssd1 vccd1 vccd1 _21416_/C sky130_fd_sc_hd__inv_2
XFILLER_0_153_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13330_ _26318_/Q _19616_/A vssd1 vssd1 vccd1 vccd1 _14620_/A sky130_fd_sc_hd__xor2_1
X_22528_ _26048_/Q vssd1 vssd1 vccd1 vccd1 _22529_/A sky130_fd_sc_hd__inv_2
XFILLER_0_18_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25316_ _26263_/CLK hold31/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26296_ _26296_/CLK _26296_/D vssd1 vssd1 vccd1 vccd1 _26296_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_84_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13261_ _13220_/X _14584_/A _13242_/X _19458_/A vssd1 vssd1 vccd1 vccd1 _13261_/X
+ sky130_fd_sc_hd__a22o_1
X_22459_ _22448_/Y _22458_/Y _23197_/A vssd1 vssd1 vccd1 vccd1 _22459_/X sky130_fd_sc_hd__a21o_1
X_25247_ _25709_/CLK hold785/X vssd1 vssd1 vccd1 vccd1 hold783/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15000_ _14983_/Y _15032_/C _14999_/Y vssd1 vssd1 vccd1 vccd1 _15000_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_121_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13192_ _23377_/B vssd1 vssd1 vccd1 vccd1 _13192_/X sky130_fd_sc_hd__buf_4
X_25178_ _25761_/CLK hold406/X vssd1 vssd1 vccd1 vccd1 hold404/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24129_ _24835_/S vssd1 vssd1 vccd1 vccd1 _24203_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16951_ _22145_/B _16956_/B vssd1 vssd1 vccd1 vccd1 _16953_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15902_ _15956_/A hold653/X vssd1 vssd1 vccd1 vccd1 hold654/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19670_ _26252_/Q hold542/X vssd1 vssd1 vccd1 vccd1 _19670_/Y sky130_fd_sc_hd__nand2_1
X_16882_ _16883_/B _16883_/A vssd1 vssd1 vccd1 vccd1 _16882_/X sky130_fd_sc_hd__or2_1
X_18621_ _18641_/A _19444_/A vssd1 vssd1 vccd1 vccd1 _18621_/Y sky130_fd_sc_hd__nand2_1
X_15833_ _15766_/Y _15824_/A _15832_/Y vssd1 vssd1 vccd1 vccd1 _15834_/B sky130_fd_sc_hd__a21oi_1
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18552_ _20171_/B _22210_/A vssd1 vssd1 vccd1 vccd1 _20162_/A sky130_fd_sc_hd__nand2_2
X_15764_ _15764_/A _15764_/B vssd1 vssd1 vccd1 vccd1 _15764_/Y sky130_fd_sc_hd__nand2_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _26257_/Q _25626_/Q vssd1 vssd1 vccd1 vccd1 _14428_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ _17605_/A _17503_/B vssd1 vssd1 vccd1 vccd1 _17503_/Y sky130_fd_sc_hd__nand2_1
X_14715_ _14721_/B _21797_/A vssd1 vssd1 vccd1 vccd1 _21796_/B sky130_fd_sc_hd__xnor2_2
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18483_ _18483_/A _18483_/B vssd1 vssd1 vccd1 vccd1 _22119_/A sky130_fd_sc_hd__nand2_1
X_15695_ _15695_/A _15695_/B vssd1 vssd1 vccd1 vccd1 _15698_/A sky130_fd_sc_hd__nand2_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17434_ _17434_/A _17434_/B vssd1 vssd1 vccd1 vccd1 _17434_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_184_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14646_ _15464_/A vssd1 vssd1 vccd1 vccd1 _14646_/X sky130_fd_sc_hd__buf_6
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_106_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _25422_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_19 _17456_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17365_ _17365_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17365_/Y sky130_fd_sc_hd__nand2_1
X_14577_ _14575_/Y hold36/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19104_ _20986_/A vssd1 vssd1 vccd1 vccd1 _19104_/X sky130_fd_sc_hd__buf_12
X_16316_ _16314_/Y _16315_/Y _16076_/X vssd1 vssd1 vccd1 vccd1 hold959/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_166_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ hold534/X _13527_/Y _12558_/B vssd1 vssd1 vccd1 vccd1 hold535/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17296_ _17393_/A _17296_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17296_/X sky130_fd_sc_hd__and3_1
XFILLER_0_42_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19035_ _19035_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _19035_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16247_ hold889/X vssd1 vssd1 vccd1 vccd1 _16250_/B sky130_fd_sc_hd__inv_2
X_13459_ _13220_/A _14687_/A _13242_/A _25709_/Q vssd1 vssd1 vccd1 vccd1 _13459_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16178_ _16676_/A _15141_/A _16177_/Y vssd1 vssd1 vccd1 vccd1 _16180_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_141_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15129_ _15112_/X _15162_/B _15128_/Y vssd1 vssd1 vccd1 vccd1 _15129_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19937_ _19937_/A _19948_/A vssd1 vssd1 vccd1 vccd1 _19939_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_177_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19868_ _19867_/Y _19130_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19870_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_177_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18819_ _19026_/A _18819_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18819_/X sky130_fd_sc_hd__and3_1
X_19799_ _26261_/Q hold404/X vssd1 vssd1 vccd1 vccd1 _19799_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_179_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21830_ _22653_/A _21830_/B vssd1 vssd1 vccd1 vccd1 _21830_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21761_ _21759_/X _14270_/A _21760_/Y _14712_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _21762_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_148_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20712_ _20712_/A _20712_/B vssd1 vssd1 vccd1 vccd1 _20716_/A sky130_fd_sc_hd__nand2_1
X_23500_ _24944_/S hold320/A _23499_/X vssd1 vssd1 vccd1 vccd1 _23500_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24480_ hold2617/X hold2573/X _24510_/S vssd1 vssd1 vccd1 vccd1 _24481_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_53_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21692_ _21692_/A _21692_/B vssd1 vssd1 vccd1 vccd1 _21694_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23431_ _23419_/X _23430_/X _24949_/S vssd1 vssd1 vccd1 vccd1 _23431_/X sky130_fd_sc_hd__mux2_1
X_20643_ _20643_/A _20643_/B _20643_/C vssd1 vssd1 vccd1 vccd1 _20644_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_19_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26150_ _26151_/CLK _26150_/D vssd1 vssd1 vccd1 vccd1 _26150_/Q sky130_fd_sc_hd__dfxtp_1
X_23362_ _23362_/A vssd1 vssd1 vccd1 vccd1 _25935_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20574_ _20574_/A _21252_/B _20574_/C vssd1 vssd1 vccd1 vccd1 _20575_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_18_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22313_ _22313_/A _25856_/Q vssd1 vssd1 vccd1 vccd1 _22314_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_15_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25101_ _26184_/CLK _25101_/D vssd1 vssd1 vccd1 vccd1 _25101_/Q sky130_fd_sc_hd__dfxtp_1
X_26081_ _26084_/CLK _26081_/D vssd1 vssd1 vccd1 vccd1 _26081_/Q sky130_fd_sc_hd__dfxtp_1
X_23293_ hold855/X _23293_/B vssd1 vssd1 vccd1 vccd1 _23294_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25032_ _26117_/CLK _25032_/D vssd1 vssd1 vccd1 vccd1 _25032_/Q sky130_fd_sc_hd__dfxtp_1
X_22244_ _22874_/B vssd1 vssd1 vccd1 vccd1 _22875_/A sky130_fd_sc_hd__inv_2
XFILLER_0_30_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22175_ _22175_/A _22387_/B vssd1 vssd1 vccd1 vccd1 _22175_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21126_ _21235_/A _21844_/A vssd1 vssd1 vccd1 vccd1 _21126_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_100_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25934_ _25938_/CLK _25934_/D vssd1 vssd1 vccd1 vccd1 _25934_/Q sky130_fd_sc_hd__dfxtp_1
X_21057_ _21561_/C _21513_/C vssd1 vssd1 vccd1 vccd1 _21059_/A sky130_fd_sc_hd__nand2_1
X_20008_ _20008_/A _20008_/B vssd1 vssd1 vccd1 vccd1 _21677_/A sky130_fd_sc_hd__nand2_4
X_25865_ _25865_/CLK _25865_/D vssd1 vssd1 vccd1 vccd1 _25865_/Q sky130_fd_sc_hd__dfxtp_2
X_24816_ _24816_/A vssd1 vssd1 vccd1 vccd1 _26333_/D sky130_fd_sc_hd__clkbuf_1
X_12830_ _26229_/Q _25598_/Q vssd1 vssd1 vccd1 vccd1 _14337_/A sky130_fd_sc_hd__xor2_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25796_ _25796_/CLK _25796_/D vssd1 vssd1 vccd1 vccd1 _25796_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _17045_/B _14264_/A vssd1 vssd1 vccd1 vccd1 _12761_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24747_ _24747_/A vssd1 vssd1 vccd1 vccd1 _26310_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21959_ _18073_/B _17112_/B _18075_/A vssd1 vssd1 vccd1 vccd1 _21960_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_57_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _14500_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14500_/Y sky130_fd_sc_hd__nand2_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12692_/A _24836_/B _12696_/A vssd1 vssd1 vccd1 vccd1 _12692_/X sky130_fd_sc_hd__and3_1
X_15480_ _15480_/A _16848_/A vssd1 vssd1 vccd1 vccd1 _15481_/B sky130_fd_sc_hd__nor2_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24678_ _24678_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24679_/A sky130_fd_sc_hd__and2_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _14431_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14431_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_181_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23629_ _23629_/A _23629_/B vssd1 vssd1 vccd1 vccd1 _23630_/A sky130_fd_sc_hd__and2_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17150_ _17150_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17150_/Y sky130_fd_sc_hd__nand2_1
X_14362_ _14404_/A hold50/X vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16101_ _16212_/A hold593/X vssd1 vssd1 vccd1 vccd1 hold594/A sky130_fd_sc_hd__nand2_1
X_13313_ _18799_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13313_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17081_ _17079_/Y _17080_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _17081_/Y sky130_fd_sc_hd__a21oi_1
X_14293_ _14344_/A hold155/X vssd1 vssd1 vccd1 vccd1 hold156/A sky130_fd_sc_hd__nand2_1
XFILLER_0_80_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26279_ _26279_/CLK _26279_/D vssd1 vssd1 vccd1 vccd1 _26279_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_150_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16032_ _16032_/A _16697_/B _16040_/A vssd1 vssd1 vccd1 vccd1 _16032_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_122_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13244_ _26176_/Q _13239_/X _13243_/X vssd1 vssd1 vccd1 vccd1 _13244_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_62_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ _13109_/X _13173_/X _13096_/X _13174_/X vssd1 vssd1 vccd1 vccd1 hold980/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17983_ _17983_/A _17983_/B vssd1 vssd1 vccd1 vccd1 _22189_/A sky130_fd_sc_hd__nand2_1
X_19722_ _19714_/X _19721_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19722_/Y sky130_fd_sc_hd__o21ai_1
X_16934_ _16932_/Y _16933_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16934_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19653_ _21099_/A vssd1 vssd1 vccd1 vccd1 _19653_/X sky130_fd_sc_hd__buf_8
X_16865_ _16977_/A _16865_/B vssd1 vssd1 vccd1 vccd1 _16865_/Y sky130_fd_sc_hd__nand2_1
X_18604_ _22297_/B _25628_/Q vssd1 vssd1 vccd1 vccd1 _18606_/A sky130_fd_sc_hd__nand2_1
X_15816_ _15816_/A _15816_/B vssd1 vssd1 vccd1 vccd1 _15817_/B sky130_fd_sc_hd__and2_1
X_19584_ _26246_/Q _19483_/X hold545/X vssd1 vssd1 vccd1 vccd1 _19584_/Y sky130_fd_sc_hd__a21oi_1
X_16796_ _16796_/A _16796_/B vssd1 vssd1 vccd1 vccd1 _16796_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18535_ _18535_/A _18535_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18535_/X sky130_fd_sc_hd__and3_1
X_15747_ _15764_/B vssd1 vssd1 vccd1 vccd1 _15750_/B sky130_fd_sc_hd__inv_2
XFILLER_0_133_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12959_ _17486_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12959_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18466_ _18793_/A _25749_/Q _18891_/C vssd1 vssd1 vccd1 vccd1 _18467_/C sky130_fd_sc_hd__nand3_1
X_15678_ _15678_/A _15692_/B vssd1 vssd1 vccd1 vccd1 _15678_/Y sky130_fd_sc_hd__nand2_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17417_ _17467_/A _17417_/B vssd1 vssd1 vccd1 vccd1 _17417_/Y sky130_fd_sc_hd__nand2_1
X_14629_ _14629_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14629_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_157_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18397_ _18395_/Y _18396_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25664_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17348_ _25614_/Q vssd1 vssd1 vccd1 vccd1 _21129_/B sky130_fd_sc_hd__inv_2
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17279_ _25706_/Q _17279_/B vssd1 vssd1 vccd1 vccd1 _17629_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_28_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19018_ _19018_/A _19018_/B vssd1 vssd1 vccd1 vccd1 _19018_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20290_ _20290_/A _20290_/B vssd1 vssd1 vccd1 vccd1 _20292_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2703 _24832_/X vssd1 vssd1 vccd1 vccd1 _24833_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2714 _26328_/Q vssd1 vssd1 vccd1 vccd1 hold2714/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2725 _26278_/Q vssd1 vssd1 vccd1 vccd1 hold2725/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2736 _26263_/Q vssd1 vssd1 vccd1 vccd1 hold2736/X sky130_fd_sc_hd__dlygate4sd3_1
X_23980_ hold2422/X hold2178/X _24001_/S vssd1 vssd1 vccd1 vccd1 _23981_/A sky130_fd_sc_hd__mux2_1
Xhold2747 _24998_/Q vssd1 vssd1 vccd1 vccd1 _12491_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2758 _25890_/Q vssd1 vssd1 vccd1 vccd1 hold2758/X sky130_fd_sc_hd__dlygate4sd3_1
X_22931_ _22931_/A _22931_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22933_/A sky130_fd_sc_hd__or3_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25650_ _25650_/CLK _25650_/D vssd1 vssd1 vccd1 vccd1 _25650_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_79_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22862_ _22862_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22862_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24601_ _24601_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24602_/A sky130_fd_sc_hd__and2_1
X_21813_ _19458_/A _21812_/A _21812_/Y vssd1 vssd1 vccd1 vccd1 _21815_/A sky130_fd_sc_hd__o21ai_2
X_22793_ _22793_/A _22793_/B vssd1 vssd1 vccd1 vccd1 _22794_/B sky130_fd_sc_hd__nand2_1
X_25581_ _26269_/CLK _25581_/D vssd1 vssd1 vccd1 vccd1 _25581_/Q sky130_fd_sc_hd__dfxtp_4
X_21744_ _21744_/A _21744_/B vssd1 vssd1 vccd1 vccd1 _22550_/A sky130_fd_sc_hd__nand2_2
X_24532_ hold2563/X _26241_/Q _24587_/S vssd1 vssd1 vccd1 vccd1 _24532_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_182_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24463_ _24463_/A vssd1 vssd1 vccd1 vccd1 _26218_/D sky130_fd_sc_hd__clkbuf_1
X_21675_ _21675_/A _21675_/B _21675_/C vssd1 vssd1 vccd1 vccd1 _21679_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_171_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26202_ _26202_/CLK _26202_/D vssd1 vssd1 vccd1 vccd1 _26202_/Q sky130_fd_sc_hd__dfxtp_1
X_23414_ _24940_/S hold290/A _23413_/X vssd1 vssd1 vccd1 vccd1 _23414_/Y sky130_fd_sc_hd__o21ai_1
X_20626_ _20628_/B _20628_/C vssd1 vssd1 vccd1 vccd1 _20627_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24394_ hold2464/X _26196_/Q _24433_/S vssd1 vssd1 vccd1 vccd1 _24394_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23345_ _23345_/A vssd1 vssd1 vccd1 vccd1 _23347_/B sky130_fd_sc_hd__inv_2
XFILLER_0_116_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26133_ _26136_/CLK _26133_/D vssd1 vssd1 vccd1 vccd1 _26133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20557_ _20557_/A _22463_/B vssd1 vssd1 vccd1 vccd1 _20558_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23276_ _23276_/A hold829/X _23276_/C vssd1 vssd1 vccd1 vccd1 _23278_/A sky130_fd_sc_hd__and3_1
X_26064_ _26064_/CLK _26064_/D vssd1 vssd1 vccd1 vccd1 _26064_/Q sky130_fd_sc_hd__dfxtp_1
X_20488_ _20488_/A _20488_/B vssd1 vssd1 vccd1 vccd1 _21563_/A sky130_fd_sc_hd__nand2_4
X_22227_ _22227_/A _23138_/A _22227_/C vssd1 vssd1 vccd1 vccd1 _22227_/Y sky130_fd_sc_hd__nand3_1
X_25015_ _25596_/CLK _25015_/D vssd1 vssd1 vccd1 vccd1 _25015_/Q sky130_fd_sc_hd__dfxtp_1
X_22158_ _22651_/A _22823_/B vssd1 vssd1 vccd1 vccd1 _22168_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_100_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21109_ _21109_/A _21109_/B _21109_/C vssd1 vssd1 vccd1 vccd1 _21110_/B sky130_fd_sc_hd__nand3_1
X_14980_ _14980_/A _14980_/B vssd1 vssd1 vccd1 vccd1 _14981_/B sky130_fd_sc_hd__nand2_1
X_22089_ _22086_/Y _22088_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _22089_/Y sky130_fd_sc_hd__a21oi_1
X_25917_ _26341_/CLK hold831/X vssd1 vssd1 vccd1 vccd1 hold829/A sky130_fd_sc_hd__dfxtp_1
X_13931_ _14000_/A hold686/X vssd1 vssd1 vccd1 vccd1 hold687/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16650_ _16650_/A _16650_/B vssd1 vssd1 vccd1 vccd1 _16658_/A sky130_fd_sc_hd__nand2_1
X_25848_ _26208_/CLK _25848_/D vssd1 vssd1 vccd1 vccd1 _25848_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13862_ _13880_/A hold725/X vssd1 vssd1 vccd1 vccd1 hold726/A sky130_fd_sc_hd__nand2_1
X_15601_ _15602_/A _15603_/A vssd1 vssd1 vccd1 vccd1 _15605_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12813_ _26226_/Q _25595_/Q vssd1 vssd1 vccd1 vccd1 _14328_/A sky130_fd_sc_hd__xor2_2
X_16581_ _16581_/A _16686_/B _16581_/C vssd1 vssd1 vccd1 vccd1 _16581_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_187_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25779_ _25779_/CLK _25779_/D vssd1 vssd1 vccd1 vccd1 _25779_/Q sky130_fd_sc_hd__dfxtp_1
X_13793_ _14170_/A vssd1 vssd1 vccd1 vccd1 _13793_/X sky130_fd_sc_hd__buf_12
XFILLER_0_186_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18320_ _21129_/B _19488_/A vssd1 vssd1 vccd1 vccd1 _18321_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15532_ _15550_/B vssd1 vssd1 vccd1 vccd1 _15535_/B sky130_fd_sc_hd__inv_2
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _14260_/A hold77/X vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _18251_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18251_/Y sky130_fd_sc_hd__nand2_1
X_15463_ _15463_/A _15463_/B vssd1 vssd1 vccd1 vccd1 _15463_/Y sky130_fd_sc_hd__nand2_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _12676_/B _12676_/A vssd1 vssd1 vccd1 vccd1 _12677_/A sky130_fd_sc_hd__or2_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17202_ _17202_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17202_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_38_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14414_ _14465_/A hold308/X vssd1 vssd1 vccd1 vccd1 hold309/A sky130_fd_sc_hd__nand2_1
XFILLER_0_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18182_ _18180_/Y _18181_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25654_/D sky130_fd_sc_hd__a21oi_1
X_15394_ _15394_/A vssd1 vssd1 vccd1 vccd1 _15403_/B sky130_fd_sc_hd__inv_2
XFILLER_0_182_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17133_ _17470_/A _17548_/A vssd1 vssd1 vccd1 vccd1 _17134_/B sky130_fd_sc_hd__xnor2_1
X_14345_ _14345_/A vssd1 vssd1 vccd1 vccd1 _14345_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold609 hold609/A vssd1 vssd1 vccd1 vccd1 hold609/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17064_ _17272_/A _17064_/B vssd1 vssd1 vccd1 vccd1 _17064_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_64_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14276_ _14277_/C _14274_/X _12482_/A _14275_/Y _14910_/B vssd1 vssd1 vccd1 vccd1
+ _14276_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16015_ _16027_/B _16016_/A vssd1 vssd1 vccd1 vccd1 _16015_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13227_ _13227_/A vssd1 vssd1 vccd1 vccd1 _19388_/A sky130_fd_sc_hd__buf_4
XFILLER_0_110_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13158_ _13158_/A vssd1 vssd1 vccd1 vccd1 _19230_/A sky130_fd_sc_hd__buf_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17966_ _18252_/A _17966_/B vssd1 vssd1 vccd1 vccd1 _17966_/Y sky130_fd_sc_hd__nand2_1
X_13089_ _13049_/X _14494_/A _13067_/X _25647_/Q vssd1 vssd1 vccd1 vccd1 _13089_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1309 _19482_/Y vssd1 vssd1 vccd1 vccd1 _25735_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16917_ _16980_/A _25571_/Q vssd1 vssd1 vccd1 vccd1 _16917_/Y sky130_fd_sc_hd__nand2_1
X_19705_ _19706_/B _19706_/A vssd1 vssd1 vccd1 vccd1 _19705_/X sky130_fd_sc_hd__or2_1
X_17897_ _20474_/B _22133_/A vssd1 vssd1 vccd1 vccd1 _20467_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16848_ _16848_/A _16848_/B vssd1 vssd1 vccd1 vccd1 _16848_/Y sky130_fd_sc_hd__nand2_1
X_19636_ _19634_/X _19635_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19636_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_189_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19567_ _19559_/X _19566_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19567_/Y sky130_fd_sc_hd__o21ai_1
X_16779_ _22683_/B _16977_/A _16775_/Y _16778_/Y _12702_/A vssd1 vssd1 vccd1 vccd1
+ _16779_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_0_34_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18518_ _18641_/A _19373_/A vssd1 vssd1 vccd1 vccd1 _18518_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_34_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19498_ _19723_/A _19498_/B vssd1 vssd1 vccd1 vccd1 _19498_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18449_ _18955_/A _18449_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18450_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21460_ _21573_/A _21460_/B vssd1 vssd1 vccd1 vccd1 _21460_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_69_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20411_ _21225_/B _21531_/A vssd1 vssd1 vccd1 vccd1 _20414_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21391_ _26320_/Q hold748/X vssd1 vssd1 vccd1 vccd1 _21391_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_172_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_6__f_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _25759_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23130_ _16956_/B _22421_/A _23124_/X _23125_/Y _23129_/X vssd1 vssd1 vccd1 vccd1
+ _23131_/A sky130_fd_sc_hd__a221o_1
X_20342_ _26285_/Q hold389/X vssd1 vssd1 vccd1 vccd1 _20342_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23061_ _15668_/B _22893_/A _22829_/X vssd1 vssd1 vccd1 vccd1 _23061_/Y sky130_fd_sc_hd__a21oi_1
X_20273_ _20273_/A _20273_/B vssd1 vssd1 vccd1 vccd1 _20277_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_113_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22012_ _22012_/A _22012_/B vssd1 vssd1 vccd1 vccd1 _23184_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2500 _12670_/Y vssd1 vssd1 vccd1 vccd1 _12672_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2511 _23974_/X vssd1 vssd1 vccd1 vccd1 _23975_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2522 _25685_/Q vssd1 vssd1 vccd1 vccd1 _13316_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2533 _24769_/X vssd1 vssd1 vccd1 vccd1 _24770_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2544 _25903_/Q vssd1 vssd1 vccd1 vccd1 _17706_/A sky130_fd_sc_hd__buf_1
Xhold2555 _26226_/Q vssd1 vssd1 vccd1 vccd1 hold2555/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1810 _25625_/Q vssd1 vssd1 vccd1 vccd1 _17510_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1821 _25412_/Q vssd1 vssd1 vccd1 vccd1 _14903_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2566 _24474_/X vssd1 vssd1 vccd1 vccd1 _24475_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2577 _25471_/Q vssd1 vssd1 vccd1 vccd1 _15743_/A sky130_fd_sc_hd__dlygate4sd3_1
X_23963_ _23963_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23964_/A sky130_fd_sc_hd__and2_1
Xhold1832 _26096_/Q vssd1 vssd1 vccd1 vccd1 hold1832/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2588 _25908_/Q vssd1 vssd1 vccd1 vccd1 _23215_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1843 _25841_/Q vssd1 vssd1 vccd1 vccd1 _21862_/B sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_95_clk clkbuf_leaf_95_clk/A vssd1 vssd1 vccd1 vccd1 _26001_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1854 _25844_/Q vssd1 vssd1 vccd1 vccd1 _21965_/B sky130_fd_sc_hd__dlygate4sd3_1
X_25702_ _25708_/CLK _25702_/D vssd1 vssd1 vccd1 vccd1 _25702_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2599 _26231_/Q vssd1 vssd1 vccd1 vccd1 hold2599/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22914_ _22914_/A _22914_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22916_/A sky130_fd_sc_hd__or3_1
Xhold1865 _17569_/Y vssd1 vssd1 vccd1 vccd1 _25633_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1876 _25628_/Q vssd1 vssd1 vccd1 vccd1 _17532_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1887 _14910_/Y vssd1 vssd1 vccd1 vccd1 _14911_/A sky130_fd_sc_hd__dlygate4sd3_1
X_23894_ _23894_/A vssd1 vssd1 vccd1 vccd1 _26035_/D sky130_fd_sc_hd__clkbuf_1
Xhold1898 _25708_/Q vssd1 vssd1 vccd1 vccd1 _19078_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25633_ _25716_/CLK _25633_/D vssd1 vssd1 vccd1 vccd1 _25633_/Q sky130_fd_sc_hd__dfxtp_4
X_22845_ _23188_/A _22845_/B vssd1 vssd1 vccd1 vccd1 _22845_/X sky130_fd_sc_hd__or2_1
XFILLER_0_6_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25564_ _26066_/CLK _25564_/D vssd1 vssd1 vccd1 vccd1 _25564_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22776_ _22776_/A _22776_/B vssd1 vssd1 vccd1 vccd1 _22777_/B sky130_fd_sc_hd__nand2_1
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24515_ _24515_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24516_/A sky130_fd_sc_hd__and2_1
XFILLER_0_176_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21727_ _21727_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _21727_/X sky130_fd_sc_hd__and2_1
XFILLER_0_137_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25495_ _25495_/CLK hold595/X vssd1 vssd1 vccd1 vccd1 hold593/A sky130_fd_sc_hd__dfxtp_1
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24446_ input6/X hold2737/X _24510_/S vssd1 vssd1 vccd1 vccd1 _24447_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21658_ _21660_/B _21709_/B vssd1 vssd1 vccd1 vccd1 _21659_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_124_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20609_ _21611_/A _21335_/C vssd1 vssd1 vccd1 vccd1 _20610_/B sky130_fd_sc_hd__nand2_1
X_21589_ _22586_/A vssd1 vssd1 vccd1 vccd1 _22058_/A sky130_fd_sc_hd__clkbuf_8
X_24377_ _24377_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24378_/A sky130_fd_sc_hd__and2_1
XFILLER_0_22_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26116_ _26116_/CLK _26116_/D vssd1 vssd1 vccd1 vccd1 _26116_/Q sky130_fd_sc_hd__dfxtp_1
X_14130_ _14180_/A _14130_/B vssd1 vssd1 vccd1 vccd1 _14130_/Y sky130_fd_sc_hd__nand2_1
X_23328_ _23330_/B _23330_/A vssd1 vssd1 vccd1 vccd1 _23336_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_34_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26047_ _26047_/CLK _26047_/D vssd1 vssd1 vccd1 vccd1 _26047_/Q sky130_fd_sc_hd__dfxtp_1
X_14061_ _14061_/A _14061_/B vssd1 vssd1 vccd1 vccd1 _14061_/Y sky130_fd_sc_hd__nand2_1
X_23259_ _23484_/B _23267_/B vssd1 vssd1 vccd1 vccd1 _23264_/A sky130_fd_sc_hd__or2_1
XFILLER_0_104_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13012_ _12930_/X _13010_/X _13005_/X _13011_/X vssd1 vssd1 vccd1 vccd1 _13012_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17820_ _17818_/X _17528_/X _17819_/X vssd1 vssd1 vccd1 vccd1 _17821_/A sky130_fd_sc_hd__a21o_1
X_17751_ _17752_/B _17830_/A vssd1 vssd1 vccd1 vccd1 _17753_/A sky130_fd_sc_hd__nor2_1
X_14963_ _14963_/A _14963_/B vssd1 vssd1 vccd1 vccd1 _14982_/B sky130_fd_sc_hd__nand2_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_86_clk clkbuf_leaf_95_clk/A vssd1 vssd1 vccd1 vccd1 _26053_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16702_ _16702_/A vssd1 vssd1 vccd1 vccd1 _16976_/B sky130_fd_sc_hd__buf_6
XFILLER_0_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13914_ _18124_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13914_/Y sky130_fd_sc_hd__nor2_1
X_17682_ _17719_/B _25905_/Q vssd1 vssd1 vccd1 vccd1 _17717_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_187_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14894_ _14900_/B _22387_/A vssd1 vssd1 vccd1 vccd1 _22386_/B sky130_fd_sc_hd__xnor2_2
X_19421_ _19421_/A _19421_/B vssd1 vssd1 vccd1 vccd1 _19421_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16633_ _16647_/A _16634_/A vssd1 vssd1 vccd1 vccd1 _16635_/A sky130_fd_sc_hd__or2_1
X_13845_ _25770_/Q vssd1 vssd1 vccd1 vccd1 _18894_/B sky130_fd_sc_hd__inv_2
XFILLER_0_162_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19352_ _19344_/X _19351_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19352_/Y sky130_fd_sc_hd__o21ai_1
X_16564_ _16564_/A _16564_/B vssd1 vssd1 vccd1 vccd1 _16566_/A sky130_fd_sc_hd__nand2_1
X_13776_ _18673_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13776_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18303_ _18445_/A _18307_/B vssd1 vssd1 vccd1 vccd1 _18305_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15515_ _15515_/A _16862_/A vssd1 vssd1 vccd1 vccd1 _15516_/B sky130_fd_sc_hd__nor2_1
X_12727_ _13465_/A _14267_/A vssd1 vssd1 vccd1 vccd1 _16774_/B sky130_fd_sc_hd__nand2_2
X_19283_ _19452_/A _19283_/B vssd1 vssd1 vccd1 vccd1 _19283_/Y sky130_fd_sc_hd__nand2_1
X_16495_ _16495_/A _16495_/B vssd1 vssd1 vccd1 vccd1 _16599_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_45_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18234_ _19430_/A vssd1 vssd1 vccd1 vccd1 _21738_/B sky130_fd_sc_hd__inv_2
XFILLER_0_183_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15446_ _15446_/A _15446_/B vssd1 vssd1 vccd1 vccd1 _15447_/B sky130_fd_sc_hd__nand2_1
X_12658_ _12658_/A vssd1 vssd1 vccd1 vccd1 _24983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18165_ _18165_/A _18165_/B vssd1 vssd1 vccd1 vccd1 _21937_/A sky130_fd_sc_hd__nand2_1
X_15377_ _15405_/B _15378_/A vssd1 vssd1 vccd1 vccd1 _15377_/X sky130_fd_sc_hd__or2_1
XFILLER_0_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12589_ _12589_/A vssd1 vssd1 vccd1 vccd1 _24970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_10_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _26263_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17116_ _19230_/A _17116_/B vssd1 vssd1 vccd1 vccd1 _17463_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14328_ _14328_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14328_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_64_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18096_ _18446_/A _25733_/Q _21716_/A vssd1 vssd1 vccd1 vccd1 _18097_/C sky130_fd_sc_hd__nand3_1
Xhold406 hold406/A vssd1 vssd1 vccd1 vccd1 hold406/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold417 hold417/A vssd1 vssd1 vccd1 vccd1 hold417/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 hold428/A vssd1 vssd1 vccd1 vccd1 hold428/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17047_ _17047_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17047_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold439 hold439/A vssd1 vssd1 vccd1 vccd1 hold439/X sky130_fd_sc_hd__dlygate4sd3_1
X_14259_ hold432/X _14258_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold433/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_14__f_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_14__f_clk/X
+ sky130_fd_sc_hd__clkbuf_16
X_18998_ _19026_/A _18998_/B _22786_/A vssd1 vssd1 vccd1 vccd1 _18998_/X sky130_fd_sc_hd__and3_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 _16723_/Y vssd1 vssd1 vccd1 vccd1 _25542_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 _25565_/Q vssd1 vssd1 vccd1 vccd1 _16879_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1128 _16019_/Y vssd1 vssd1 vccd1 vccd1 _25489_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17949_ _21764_/B _25602_/Q vssd1 vssd1 vccd1 vccd1 _17951_/A sky130_fd_sc_hd__nand2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_clk clkbuf_leaf_82_clk/A vssd1 vssd1 vccd1 vccd1 _25876_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1139 _25029_/Q vssd1 vssd1 vccd1 vccd1 _17373_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20960_ _20960_/A _20960_/B vssd1 vssd1 vccd1 vccd1 _20961_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_174_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19619_ _19635_/B _19706_/B vssd1 vssd1 vccd1 vccd1 _19621_/A sky130_fd_sc_hd__xnor2_1
X_20891_ _21467_/B vssd1 vssd1 vccd1 vccd1 _21464_/C sky130_fd_sc_hd__inv_2
XFILLER_0_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22630_ _26052_/Q vssd1 vssd1 vccd1 vccd1 _22631_/A sky130_fd_sc_hd__inv_2
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22561_ _22561_/A _22561_/B vssd1 vssd1 vccd1 vccd1 _22561_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_119_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24300_ _24300_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24301_/A sky130_fd_sc_hd__and2_1
X_21512_ _21514_/A _21563_/A vssd1 vssd1 vccd1 vccd1 _21513_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_57_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22492_ _22493_/B _22493_/A vssd1 vssd1 vccd1 vccd1 _22494_/A sky130_fd_sc_hd__or2_1
XFILLER_0_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25280_ _26235_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24231_ hold2312/X _26143_/Q _24279_/S vssd1 vssd1 vccd1 vccd1 _24231_/X sky130_fd_sc_hd__mux2_1
X_21443_ _21443_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21443_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24162_ _24162_/A vssd1 vssd1 vccd1 vccd1 _26120_/D sky130_fd_sc_hd__clkbuf_1
X_21374_ _26319_/Q _21228_/X hold731/X vssd1 vssd1 vccd1 vccd1 _21377_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23113_ _23113_/A _23193_/B _23113_/C vssd1 vssd1 vccd1 vccd1 _23113_/X sky130_fd_sc_hd__and3_1
X_20325_ _22937_/B vssd1 vssd1 vccd1 vccd1 _22332_/B sky130_fd_sc_hd__inv_2
X_24093_ _24093_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24094_/A sky130_fd_sc_hd__and2_1
Xhold940 hold940/A vssd1 vssd1 vccd1 vccd1 hold940/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold951 hold951/A vssd1 vssd1 vccd1 vccd1 hold951/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 hold962/A vssd1 vssd1 vccd1 vccd1 hold962/X sky130_fd_sc_hd__dlygate4sd3_1
X_23044_ _23188_/A _23044_/B vssd1 vssd1 vccd1 vccd1 _23044_/X sky130_fd_sc_hd__or2_1
Xhold973 hold973/A vssd1 vssd1 vccd1 vccd1 hold973/X sky130_fd_sc_hd__dlygate4sd3_1
X_20256_ _21114_/C vssd1 vssd1 vccd1 vccd1 _21117_/B sky130_fd_sc_hd__inv_2
Xhold984 hold984/A vssd1 vssd1 vccd1 vccd1 hold984/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 hold995/A vssd1 vssd1 vccd1 vccd1 hold995/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20187_ _20187_/A _20187_/B _20981_/B vssd1 vssd1 vccd1 vccd1 _20188_/B sky130_fd_sc_hd__nand3_1
Xhold2330 _24600_/X vssd1 vssd1 vccd1 vccd1 _24601_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2341 _24172_/X vssd1 vssd1 vccd1 vccd1 _24173_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2352 _26147_/Q vssd1 vssd1 vccd1 vccd1 hold2352/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24995_ _25422_/CLK hold412/X vssd1 vssd1 vccd1 vccd1 hold410/A sky130_fd_sc_hd__dfxtp_1
Xhold2363 _26197_/Q vssd1 vssd1 vccd1 vccd1 hold2363/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2374 _25428_/Q vssd1 vssd1 vccd1 vccd1 _15027_/B sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_68_clk _25472_/CLK vssd1 vssd1 vccd1 vccd1 _25878_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1640 _17454_/Y vssd1 vssd1 vccd1 vccd1 _25617_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2385 _24323_/X vssd1 vssd1 vccd1 vccd1 _24324_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2396 _15105_/Y vssd1 vssd1 vccd1 vccd1 _25435_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1651 _25830_/Q vssd1 vssd1 vccd1 vccd1 _21606_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23946_ _23946_/A vssd1 vssd1 vccd1 vccd1 _26050_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1662 _22773_/Y vssd1 vssd1 vccd1 vccd1 _25875_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1673 hold2753/X vssd1 vssd1 vccd1 vccd1 _17867_/B sky130_fd_sc_hd__buf_2
XFILLER_0_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1684 _22822_/Y vssd1 vssd1 vccd1 vccd1 _25878_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1695 _19201_/Y vssd1 vssd1 vccd1 vccd1 _25715_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23877_ hold2240/X hold2075/X _23907_/S vssd1 vssd1 vccd1 vccd1 _23878_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_98_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25616_ _26119_/CLK _25616_/D vssd1 vssd1 vccd1 vccd1 _25616_/Q sky130_fd_sc_hd__dfxtp_2
X_13630_ _13642_/A hold841/X vssd1 vssd1 vccd1 vccd1 _13630_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_184_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22828_ _23188_/A _22828_/B vssd1 vssd1 vccd1 vccd1 _22828_/X sky130_fd_sc_hd__or2_1
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25547_ _25875_/CLK _25547_/D vssd1 vssd1 vccd1 vccd1 _25547_/Q sky130_fd_sc_hd__dfxtp_1
X_13561_ _13642_/A hold560/X vssd1 vssd1 vccd1 vccd1 hold561/A sky130_fd_sc_hd__nand2_1
XFILLER_0_183_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22759_ _22759_/A _23072_/B vssd1 vssd1 vccd1 vccd1 _22760_/B sky130_fd_sc_hd__nand2_1
X_15300_ _22709_/B _15300_/B vssd1 vssd1 vccd1 vccd1 _22706_/B sky130_fd_sc_hd__xor2_1
X_12512_ _24983_/Q _24982_/Q _24981_/Q _24980_/Q vssd1 vssd1 vccd1 vccd1 _12514_/C
+ sky130_fd_sc_hd__or4_1
X_16280_ _16490_/A vssd1 vssd1 vccd1 vccd1 _16287_/B sky130_fd_sc_hd__inv_2
X_25478_ _25495_/CLK hold776/X vssd1 vssd1 vccd1 vccd1 hold774/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13492_ _13522_/A hold766/X vssd1 vssd1 vccd1 vccd1 _13492_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15231_ _15231_/A _16754_/A vssd1 vssd1 vccd1 vccd1 _15232_/B sky130_fd_sc_hd__nor2_1
X_24429_ _24429_/A vssd1 vssd1 vccd1 vccd1 _26207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15162_ _15162_/A _15162_/B vssd1 vssd1 vccd1 vccd1 _15185_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14113_ _25813_/Q vssd1 vssd1 vccd1 vccd1 _18470_/B sky130_fd_sc_hd__inv_2
X_15093_ _15773_/S vssd1 vssd1 vccd1 vccd1 _15809_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_120_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19970_ _19970_/A _19981_/A vssd1 vssd1 vccd1 vccd1 _19972_/A sky130_fd_sc_hd__xnor2_1
X_14044_ hold372/X _14043_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold373/A sky130_fd_sc_hd__a21oi_1
X_18921_ _18919_/X _18879_/X _18920_/X vssd1 vssd1 vccd1 vccd1 _18922_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18852_ _18954_/A _25768_/Q vssd1 vssd1 vccd1 vccd1 _18854_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_98_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17803_ _17803_/A _20389_/A vssd1 vssd1 vccd1 vccd1 _19038_/A sky130_fd_sc_hd__xor2_4
X_18783_ _18781_/Y _18782_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25683_/D sky130_fd_sc_hd__a21oi_1
X_15995_ _15996_/B _15996_/A vssd1 vssd1 vccd1 vccd1 _16027_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_59_clk _25472_/CLK vssd1 vssd1 vccd1 vccd1 _25535_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17734_ _17734_/A _17734_/B _17794_/A vssd1 vssd1 vccd1 vccd1 _17735_/B sky130_fd_sc_hd__nand3_1
X_14946_ _14946_/A _14946_/B vssd1 vssd1 vccd1 vccd1 _14964_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17665_ _17665_/A _17665_/B vssd1 vssd1 vccd1 vccd1 _17666_/B sky130_fd_sc_hd__nand2_1
X_14877_ _22343_/B _15543_/B vssd1 vssd1 vccd1 vccd1 _14878_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_148_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16616_ _16676_/A _15709_/A _24952_/A vssd1 vssd1 vccd1 vccd1 _16618_/A sky130_fd_sc_hd__o21a_1
X_19404_ _20964_/A _19402_/Y _20969_/C vssd1 vssd1 vccd1 vccd1 _19493_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_134_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13828_ _18833_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13828_/Y sky130_fd_sc_hd__nor2_1
X_17596_ _17594_/X _17528_/X _17595_/X vssd1 vssd1 vccd1 vccd1 _17597_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_147_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16547_ hold904/X vssd1 vssd1 vccd1 vccd1 _16551_/B sky130_fd_sc_hd__inv_2
X_19335_ _19336_/B _19336_/A vssd1 vssd1 vccd1 vccd1 _19335_/X sky130_fd_sc_hd__or2_1
X_13759_ hold501/X _13758_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold502/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19266_ _19261_/X _18879_/X _19265_/X vssd1 vssd1 vccd1 vccd1 _19267_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_72_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16478_ _16478_/A vssd1 vssd1 vccd1 vccd1 _16479_/B sky130_fd_sc_hd__inv_2
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18217_ _18217_/A _18217_/B vssd1 vssd1 vccd1 vccd1 _22005_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_171_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15429_ _15443_/B _15430_/A vssd1 vssd1 vccd1 vccd1 _15429_/X sky130_fd_sc_hd__or2_1
XFILLER_0_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19197_ _21791_/A vssd1 vssd1 vccd1 vccd1 _20503_/B sky130_fd_sc_hd__buf_8
XFILLER_0_60_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18148_ _18146_/Y _18147_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25653_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold203 hold203/A vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold214 hold214/A vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
X_18079_ _20625_/B _19257_/A vssd1 vssd1 vccd1 vccd1 _18080_/B sky130_fd_sc_hd__nand2_1
Xhold225 hold225/A vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 hold236/A vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 hold247/A vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 hold258/A vssd1 vssd1 vccd1 vccd1 hold258/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20110_ _21401_/A _21709_/A vssd1 vssd1 vccd1 vccd1 _20117_/B sky130_fd_sc_hd__nand2_1
Xhold269 hold269/A vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__dlygate4sd3_1
X_21090_ _21090_/A _21090_/B vssd1 vssd1 vccd1 vccd1 _21091_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20041_ _20660_/A _20041_/B vssd1 vssd1 vccd1 vccd1 _20041_/Y sky130_fd_sc_hd__nand2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23800_ hold2256/X hold2067/X _23831_/S vssd1 vssd1 vccd1 vccd1 _23801_/A sky130_fd_sc_hd__mux2_1
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24780_ _24780_/A vssd1 vssd1 vccd1 vccd1 _26321_/D sky130_fd_sc_hd__clkbuf_1
X_21992_ _21992_/A _21992_/B vssd1 vssd1 vccd1 vccd1 _21994_/A sky130_fd_sc_hd__xor2_4
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23731_ _23731_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23732_/A sky130_fd_sc_hd__and2_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20943_ _20943_/A _20943_/B vssd1 vssd1 vccd1 vccd1 _20945_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23662_ hold1936/X _25960_/Q _23677_/S vssd1 vssd1 vccd1 vccd1 _23662_/X sky130_fd_sc_hd__mux2_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20874_ _26299_/Q _20731_/X hold578/X vssd1 vssd1 vccd1 vccd1 _20877_/B sky130_fd_sc_hd__a21oi_1
X_25401_ _25998_/CLK _25401_/D vssd1 vssd1 vccd1 vccd1 _25401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22613_ _22611_/X _22612_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22613_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23593_ _23593_/A _23593_/B vssd1 vssd1 vccd1 vccd1 _23593_/X sky130_fd_sc_hd__and2_1
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25332_ _26249_/CLK hold127/X vssd1 vssd1 vccd1 vccd1 hold125/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22544_ _22544_/A _22544_/B vssd1 vssd1 vccd1 vccd1 _22545_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25263_ _26219_/CLK hold103/X vssd1 vssd1 vccd1 vccd1 hold101/A sky130_fd_sc_hd__dfxtp_1
X_22475_ _22475_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _22475_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24214_ _24214_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24215_/A sky130_fd_sc_hd__and2_1
XFILLER_0_134_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21426_ _21426_/A _21426_/B vssd1 vssd1 vccd1 vccd1 _21427_/A sky130_fd_sc_hd__nand2_1
X_25194_ _26251_/CLK hold724/X vssd1 vssd1 vccd1 vccd1 hold722/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24145_ hold2323/X hold2284/X _24203_/S vssd1 vssd1 vccd1 vccd1 _24146_/A sky130_fd_sc_hd__mux2_1
X_21357_ _26318_/Q _21228_/X hold757/X vssd1 vssd1 vccd1 vccd1 _21360_/B sky130_fd_sc_hd__a21oi_1
X_20308_ _20306_/Y _20307_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _20308_/Y sky130_fd_sc_hd__a21oi_1
X_24076_ _24076_/A vssd1 vssd1 vccd1 vccd1 _26092_/D sky130_fd_sc_hd__clkbuf_1
X_21288_ _21573_/A _21288_/B vssd1 vssd1 vccd1 vccd1 _21288_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_102_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold770 hold770/A vssd1 vssd1 vccd1 vccd1 hold770/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold781 hold781/A vssd1 vssd1 vccd1 vccd1 hold781/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 hold792/A vssd1 vssd1 vccd1 vccd1 hold792/X sky130_fd_sc_hd__dlygate4sd3_1
X_23027_ _23027_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _23027_/Y sky130_fd_sc_hd__nand2_1
X_20239_ _22903_/B vssd1 vssd1 vccd1 vccd1 _22272_/B sky130_fd_sc_hd__inv_2
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2160 _24184_/X vssd1 vssd1 vccd1 vccd1 _24185_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ _14800_/A vssd1 vssd1 vccd1 vccd1 _14989_/A sky130_fd_sc_hd__inv_2
Xhold2171 _26163_/Q vssd1 vssd1 vccd1 vccd1 hold2171/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2182 _26156_/Q vssd1 vssd1 vccd1 vccd1 hold2182/X sky130_fd_sc_hd__dlygate4sd3_1
X_15780_ _16967_/A _15780_/B vssd1 vssd1 vccd1 vccd1 _15781_/B sky130_fd_sc_hd__nand2_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24978_ _24983_/CLK _24978_/D vssd1 vssd1 vccd1 vccd1 _24978_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2193 _26025_/Q vssd1 vssd1 vccd1 vccd1 hold2193/X sky130_fd_sc_hd__dlygate4sd3_1
X_12992_ _26260_/Q _25629_/Q vssd1 vssd1 vccd1 vccd1 _14437_/A sky130_fd_sc_hd__xor2_2
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1470 _21720_/Y vssd1 vssd1 vccd1 vccd1 _25837_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1481 _25550_/Q vssd1 vssd1 vccd1 vccd1 _16776_/B sky130_fd_sc_hd__buf_1
X_14731_ _14900_/A _14731_/B vssd1 vssd1 vccd1 vccd1 _14731_/Y sky130_fd_sc_hd__nand2_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23929_ input4/X hold2456/X _24001_/S vssd1 vssd1 vccd1 vccd1 _23930_/A sky130_fd_sc_hd__mux2_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1492 _21364_/Y vssd1 vssd1 vccd1 vccd1 _25815_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _17448_/X _17241_/X _17449_/X vssd1 vssd1 vccd1 vccd1 _17452_/A sky130_fd_sc_hd__a21o_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _14660_/Y hold393/X _14646_/X vssd1 vssd1 vccd1 vccd1 hold394/A sky130_fd_sc_hd__a21oi_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16401_ _16401_/A hold966/X _16401_/C vssd1 vssd1 vccd1 vccd1 _16402_/B sky130_fd_sc_hd__and3_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13613_ _25733_/Q vssd1 vssd1 vccd1 vccd1 _18101_/B sky130_fd_sc_hd__inv_2
XFILLER_0_67_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17381_ _17563_/A _17615_/B vssd1 vssd1 vccd1 vccd1 _17382_/B sky130_fd_sc_hd__xnor2_1
X_14593_ _14593_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14593_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_184_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19120_ _19950_/B _19120_/B vssd1 vssd1 vccd1 vccd1 _19120_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_95_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16332_ _16332_/A _16332_/B vssd1 vssd1 vccd1 vccd1 _16361_/A sky130_fd_sc_hd__nor2_1
X_13544_ _17895_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13544_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19051_ _19049_/Y _19050_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25704_/D sky130_fd_sc_hd__a21oi_1
X_16263_ _16263_/A _16263_/B vssd1 vssd1 vccd1 vccd1 _16269_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_153_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13475_ hold668/A vssd1 vssd1 vccd1 vccd1 _17832_/A sky130_fd_sc_hd__inv_2
X_18002_ _18529_/A _18002_/B _18083_/C vssd1 vssd1 vccd1 vccd1 _18003_/C sky130_fd_sc_hd__nand3_1
X_15214_ _15214_/A _15214_/B vssd1 vssd1 vccd1 vccd1 _15268_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_164_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16194_ _16194_/A vssd1 vssd1 vccd1 vccd1 _16208_/B sky130_fd_sc_hd__inv_2
XFILLER_0_153_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15145_ _15145_/A _15145_/B vssd1 vssd1 vccd1 vccd1 _15162_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_26_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15076_ _15076_/A _15076_/B vssd1 vssd1 vccd1 vccd1 _15077_/B sky130_fd_sc_hd__nand2_1
X_19953_ _19975_/A _19953_/B vssd1 vssd1 vccd1 vccd1 _19953_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_121_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14027_ _25799_/Q vssd1 vssd1 vccd1 vccd1 _18173_/B sky130_fd_sc_hd__inv_2
X_18904_ _18902_/Y _18903_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25689_/D sky130_fd_sc_hd__a21oi_1
X_19884_ _20828_/A _22640_/B _25642_/Q vssd1 vssd1 vccd1 vccd1 _20833_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18835_ _20720_/B _22566_/A vssd1 vssd1 vccd1 vccd1 _20711_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_101_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15978_ _15978_/A _15978_/B vssd1 vssd1 vccd1 vccd1 _15987_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_179_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18766_ _20597_/B _19802_/A vssd1 vssd1 vccd1 vccd1 _18767_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_93_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14929_ _14926_/X _14927_/Y _14928_/X vssd1 vssd1 vccd1 vccd1 _25415_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17717_ _17717_/A _17750_/B vssd1 vssd1 vccd1 vccd1 _17764_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_136_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18697_ _18899_/A _18988_/A vssd1 vssd1 vccd1 vccd1 _18698_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17648_ _17648_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _17648_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17579_ _22786_/A vssd1 vssd1 vccd1 vccd1 _18393_/C sky130_fd_sc_hd__buf_8
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19318_ _20779_/A _21764_/B _25602_/Q vssd1 vssd1 vccd1 vccd1 _20784_/C sky130_fd_sc_hd__nand3_1
X_20590_ _20590_/A _22224_/B _20590_/C vssd1 vssd1 vccd1 vccd1 _20593_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19249_ _26222_/Q hold533/X vssd1 vssd1 vccd1 vccd1 _19249_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_61_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22260_ _22561_/A _22260_/B vssd1 vssd1 vccd1 vccd1 _22260_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_26_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21211_ _21211_/A _21211_/B vssd1 vssd1 vccd1 vccd1 _21214_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_143_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22191_ _17992_/A _25788_/Q _22189_/Y _22190_/Y vssd1 vssd1 vccd1 vccd1 _22192_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21142_ _21561_/C _21613_/B vssd1 vssd1 vccd1 vccd1 _21144_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25950_ _26023_/CLK _25950_/D vssd1 vssd1 vccd1 vccd1 _25950_/Q sky130_fd_sc_hd__dfxtp_1
X_21073_ _21071_/Y _21072_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _21073_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24901_ _15866_/B _15881_/B _24945_/S vssd1 vssd1 vccd1 vccd1 _24901_/X sky130_fd_sc_hd__mux2_1
X_20024_ _20024_/A _20024_/B vssd1 vssd1 vccd1 vccd1 _20025_/B sky130_fd_sc_hd__nand2_1
X_25881_ _25901_/CLK _25881_/D vssd1 vssd1 vccd1 vccd1 _25881_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24832_ _26338_/Q hold2702/X _24835_/S vssd1 vssd1 vccd1 vccd1 _24832_/X sky130_fd_sc_hd__mux2_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24763_ _26315_/Q hold2589/X _24817_/S vssd1 vssd1 vccd1 vccd1 _24763_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_179_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21975_ _19402_/A _21974_/A _21974_/Y vssd1 vssd1 vccd1 vccd1 _21977_/A sky130_fd_sc_hd__o21ai_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23714_ hold2018/X _25977_/Q _23754_/S vssd1 vssd1 vccd1 vccd1 _23714_/X sky130_fd_sc_hd__mux2_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20926_ _20926_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _20931_/A sky130_fd_sc_hd__nand2_1
X_24694_ _24694_/A vssd1 vssd1 vccd1 vccd1 _26293_/D sky130_fd_sc_hd__clkbuf_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23645_ _23645_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23646_/A sky130_fd_sc_hd__and2_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20857_ _20860_/A _20860_/C vssd1 vssd1 vccd1 vccd1 _20858_/A sky130_fd_sc_hd__nand2_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23576_ _23573_/Y _23575_/Y _24946_/A vssd1 vssd1 vccd1 vccd1 _23576_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_107_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20788_ _20788_/A _20788_/B vssd1 vssd1 vccd1 vccd1 _21419_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_187_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25315_ _26263_/CLK hold226/X vssd1 vssd1 vccd1 vccd1 hold224/A sky130_fd_sc_hd__dfxtp_1
X_22527_ _15173_/B _22387_/B _14273_/X vssd1 vssd1 vccd1 vccd1 _22527_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26295_ _26296_/CLK _26295_/D vssd1 vssd1 vccd1 vccd1 _26295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25246_ _26339_/CLK hold828/X vssd1 vssd1 vccd1 vccd1 hold827/A sky130_fd_sc_hd__dfxtp_1
X_13260_ _26307_/Q _19458_/A vssd1 vssd1 vccd1 vccd1 _14584_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_150_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22458_ _22458_/A _22900_/B vssd1 vssd1 vccd1 vccd1 _22458_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_32_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21409_ _21636_/A _21409_/B _21408_/X vssd1 vssd1 vccd1 vccd1 _21410_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_121_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13191_ _26168_/Q _13065_/X _13190_/X vssd1 vssd1 vccd1 vccd1 _13191_/X sky130_fd_sc_hd__a21o_1
X_25177_ _25773_/CLK hold673/X vssd1 vssd1 vccd1 vccd1 hold671/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22389_ _22389_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _22389_/X sky130_fd_sc_hd__and2_1
XFILLER_0_60_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24128_ _24128_/A vssd1 vssd1 vccd1 vccd1 _26109_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16950_ _16948_/Y _16949_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _16950_/Y sky130_fd_sc_hd__a21oi_1
X_24059_ hold2239/X hold2096/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24060_/A sky130_fd_sc_hd__mux2_1
X_15901_ _15901_/A _16697_/B _15909_/A vssd1 vssd1 vccd1 vccd1 _15901_/Y sky130_fd_sc_hd__nand3_1
X_16881_ _16935_/A _16886_/B vssd1 vssd1 vccd1 vccd1 _16883_/B sky130_fd_sc_hd__nand2_1
X_15832_ _15830_/Y _15789_/B _15831_/Y vssd1 vssd1 vccd1 vccd1 _15832_/Y sky130_fd_sc_hd__o21ai_1
X_18620_ _18620_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18620_/Y sky130_fd_sc_hd__nand2_1
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _15763_/A _15764_/A _15764_/B vssd1 vssd1 vccd1 vccd1 _15824_/B sky130_fd_sc_hd__and3_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ _18551_/A _18551_/B _18551_/C vssd1 vssd1 vccd1 vccd1 _22210_/A sky130_fd_sc_hd__nand3_2
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _12930_/X _12973_/X _12917_/X _12974_/X vssd1 vssd1 vccd1 vccd1 _12975_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _14893_/A _14714_/B vssd1 vssd1 vccd1 vccd1 _21797_/A sky130_fd_sc_hd__nand2_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17502_ _17502_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17502_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_99_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18482_ _20055_/B _19602_/A vssd1 vssd1 vccd1 vccd1 _18483_/B sky130_fd_sc_hd__nand2_1
X_15694_ _15694_/A _15695_/B vssd1 vssd1 vccd1 vccd1 _15825_/A sky130_fd_sc_hd__and2_1
XFILLER_0_59_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _17601_/A _17651_/B vssd1 vssd1 vccd1 vccd1 _17434_/B sky130_fd_sc_hd__xnor2_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14645_ _14645_/A hold152/X vssd1 vssd1 vccd1 vccd1 hold153/A sky130_fd_sc_hd__nand2_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17364_ _17362_/X _17241_/X _17363_/X vssd1 vssd1 vccd1 vccd1 _17365_/A sky130_fd_sc_hd__a21o_1
X_14576_ _14585_/A hold35/X vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16315_ _16473_/A hold958/X vssd1 vssd1 vccd1 vccd1 _16315_/Y sky130_fd_sc_hd__nand2_1
X_19103_ output8/A _21203_/A vssd1 vssd1 vccd1 vccd1 _20986_/A sky130_fd_sc_hd__nor2_8
X_13527_ _13583_/A _13527_/B vssd1 vssd1 vccd1 vccd1 _13527_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_67_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17295_ _17506_/A _17295_/B vssd1 vssd1 vccd1 vccd1 _17295_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_55_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19034_ _19032_/X _18879_/X _19033_/X vssd1 vssd1 vccd1 vccd1 _19035_/A sky130_fd_sc_hd__a21o_1
X_16246_ _16246_/A _16270_/B vssd1 vssd1 vccd1 vccd1 _16252_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_179_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13458_ _26340_/Q _25709_/Q vssd1 vssd1 vccd1 vccd1 _14687_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_180_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16177_ hold860/X vssd1 vssd1 vccd1 vccd1 _16177_/Y sky130_fd_sc_hd__inv_2
X_13389_ _13389_/A vssd1 vssd1 vccd1 vccd1 _19758_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15128_ _15112_/X _15162_/B _16698_/A vssd1 vssd1 vccd1 vccd1 _15128_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15059_ _15059_/A _15059_/B vssd1 vssd1 vccd1 vccd1 _15067_/B sky130_fd_sc_hd__nand2_2
X_19936_ _19936_/A _19980_/B _19936_/C vssd1 vssd1 vccd1 vccd1 _19936_/X sky130_fd_sc_hd__and3_1
XFILLER_0_177_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19867_ _26266_/Q hold617/X vssd1 vssd1 vccd1 vccd1 _19867_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_128_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18818_ _18818_/A _18818_/B vssd1 vssd1 vccd1 vccd1 _18818_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19798_ _26261_/Q _19134_/X hold404/X vssd1 vssd1 vccd1 vccd1 _19798_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_179_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18749_ _18792_/A _18753_/B vssd1 vssd1 vccd1 vccd1 _18751_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_144_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21760_ _21760_/A _22145_/B vssd1 vssd1 vccd1 vccd1 _21760_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_176_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20711_ _20711_/A _22564_/B vssd1 vssd1 vccd1 vccd1 _20712_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_187_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21691_ _21691_/A _21691_/B _21691_/C vssd1 vssd1 vccd1 vccd1 _21695_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_136_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23430_ _23424_/X _23429_/X _24867_/S vssd1 vssd1 vccd1 vccd1 _23430_/X sky130_fd_sc_hd__mux2_1
X_20642_ _20642_/A _20642_/B vssd1 vssd1 vccd1 vccd1 _20644_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_74_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23361_ _23361_/A _23377_/B _23366_/A vssd1 vssd1 vccd1 vccd1 _23361_/X sky130_fd_sc_hd__and3_1
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20573_ _21319_/C _21596_/A vssd1 vssd1 vccd1 vccd1 _20574_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_2_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25100_ _26184_/CLK _25100_/D vssd1 vssd1 vccd1 vccd1 _25100_/Q sky130_fd_sc_hd__dfxtp_1
X_22312_ _25856_/Q _22313_/A vssd1 vssd1 vccd1 vccd1 _22314_/A sky130_fd_sc_hd__or2_1
X_26080_ _26080_/CLK _26080_/D vssd1 vssd1 vccd1 vccd1 _26080_/Q sky130_fd_sc_hd__dfxtp_1
X_23292_ _23292_/A vssd1 vssd1 vccd1 vccd1 _23298_/B sky130_fd_sc_hd__inv_2
XFILLER_0_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25031_ _26117_/CLK _25031_/D vssd1 vssd1 vccd1 vccd1 _25031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22243_ _22243_/A _22243_/B vssd1 vssd1 vccd1 vccd1 _22874_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_108_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22174_ _22680_/A vssd1 vssd1 vccd1 vccd1 _22387_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21125_ _21125_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _21125_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25933_ _25933_/CLK _25933_/D vssd1 vssd1 vccd1 vccd1 _25933_/Q sky130_fd_sc_hd__dfxtp_1
X_21056_ _21564_/B vssd1 vssd1 vccd1 vccd1 _21561_/C sky130_fd_sc_hd__inv_2
XFILLER_0_100_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20007_ _20006_/B _20007_/B _20007_/C vssd1 vssd1 vccd1 vccd1 _20008_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_185_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25864_ _25864_/CLK _25864_/D vssd1 vssd1 vccd1 vccd1 _25864_/Q sky130_fd_sc_hd__dfxtp_4
X_24815_ _24815_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24816_/A sky130_fd_sc_hd__and2_1
XFILLER_0_97_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25795_ _26287_/CLK _25795_/D vssd1 vssd1 vccd1 vccd1 _25795_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12760_ _26087_/Q _12748_/X _12759_/X vssd1 vssd1 vccd1 vccd1 _12760_/X sky130_fd_sc_hd__a21o_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24746_ _24746_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24747_/A sky130_fd_sc_hd__and2_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21958_ _21958_/A _21958_/B vssd1 vssd1 vccd1 vccd1 _21960_/A sky130_fd_sc_hd__xor2_4
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20909_ _20909_/A _20909_/B vssd1 vssd1 vccd1 vccd1 _20913_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12691_ _12713_/B _12691_/B _24989_/Q vssd1 vssd1 vccd1 vccd1 _12696_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_139_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24677_ hold2485/X _26288_/Q _24740_/S vssd1 vssd1 vccd1 vccd1 _24677_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21889_ _21889_/A _21889_/B vssd1 vssd1 vccd1 vccd1 _21891_/A sky130_fd_sc_hd__xor2_4
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14428_/Y hold240/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold241/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_166_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23628_ hold2101/X hold1947/X _23677_/S vssd1 vssd1 vccd1 vccd1 _23629_/A sky130_fd_sc_hd__mux2_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14361_ _14361_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14361_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_182_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23559_ _24922_/S hold287/A _23558_/X vssd1 vssd1 vccd1 vccd1 _23559_/Y sky130_fd_sc_hd__o21ai_1
X_16100_ _16098_/X _16099_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _16100_/X sky130_fd_sc_hd__a21o_1
X_13312_ _26187_/Q _13239_/X _13311_/X vssd1 vssd1 vccd1 vccd1 _13312_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17080_ _17272_/A _17080_/B vssd1 vssd1 vccd1 vccd1 _17080_/Y sky130_fd_sc_hd__nand2_1
X_14292_ _14292_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14292_/Y sky130_fd_sc_hd__nand2_1
X_26278_ _26279_/CLK _26278_/D vssd1 vssd1 vccd1 vccd1 _26278_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_135_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16031_ _16031_/A _16031_/B vssd1 vssd1 vccd1 vccd1 _16040_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13243_ _13220_/X _14575_/A _13242_/X _19416_/A vssd1 vssd1 vccd1 vccd1 _13243_/X
+ sky130_fd_sc_hd__a22o_1
X_25229_ _26313_/CLK hold571/X vssd1 vssd1 vccd1 vccd1 hold569/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13174_ hold979/X _13320_/B vssd1 vssd1 vccd1 vccd1 _13174_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17982_ _20547_/B _19230_/A vssd1 vssd1 vccd1 vccd1 _17983_/B sky130_fd_sc_hd__nand2_1
X_19721_ _19719_/X _19720_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19721_/Y sky130_fd_sc_hd__a21oi_1
X_16933_ _16977_/A _16933_/B vssd1 vssd1 vccd1 vccd1 _16933_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19652_ _19723_/A _19652_/B vssd1 vssd1 vccd1 vccd1 _19652_/Y sky130_fd_sc_hd__nand2_1
X_16864_ _16864_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16864_/Y sky130_fd_sc_hd__nand2_1
X_18603_ _19687_/A vssd1 vssd1 vccd1 vccd1 _22297_/B sky130_fd_sc_hd__inv_4
X_15815_ _15816_/B _15816_/A vssd1 vssd1 vccd1 vccd1 _15817_/A sky130_fd_sc_hd__nor2_1
X_16795_ _16796_/B _16796_/A vssd1 vssd1 vccd1 vccd1 _16795_/X sky130_fd_sc_hd__or2_1
X_19583_ _19581_/Y _19582_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19583_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15746_ _15746_/A _15746_/B vssd1 vssd1 vccd1 vccd1 _15764_/B sky130_fd_sc_hd__nor2_1
X_18534_ _18534_/A _18534_/B vssd1 vssd1 vccd1 vccd1 _18534_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_172_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ _26125_/Q _12907_/X _12957_/X vssd1 vssd1 vccd1 vccd1 _12958_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15677_ _15692_/B _15678_/A vssd1 vssd1 vccd1 vccd1 _15677_/X sky130_fd_sc_hd__or2_1
X_18465_ _18792_/A _18469_/B vssd1 vssd1 vccd1 vccd1 _18467_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_158_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12889_ _17373_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12889_/X sky130_fd_sc_hd__or2_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17416_ _17416_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17416_/Y sky130_fd_sc_hd__nand2_1
X_14628_ _14626_/Y hold150/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold151/A sky130_fd_sc_hd__a21oi_1
X_18396_ _18641_/A _19289_/A vssd1 vssd1 vccd1 vccd1 _18396_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_173_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17347_ _17345_/Y _17346_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _17347_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14559_ _14557_/Y hold72/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17278_ _20829_/B _25898_/Q _25834_/Q vssd1 vssd1 vccd1 vccd1 _17279_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16229_ _16238_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16229_/Y sky130_fd_sc_hd__nand2_1
X_19017_ _19017_/A _19017_/B vssd1 vssd1 vccd1 vccd1 _19018_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2704 _26302_/Q vssd1 vssd1 vccd1 vccd1 hold2704/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2715 _26220_/Q vssd1 vssd1 vccd1 vccd1 hold2715/X sky130_fd_sc_hd__dlygate4sd3_1
X_19919_ _19916_/Y _19917_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _19919_/Y sky130_fd_sc_hd__a21oi_1
Xhold2726 _26214_/Q vssd1 vssd1 vccd1 vccd1 hold2726/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2737 _26213_/Q vssd1 vssd1 vccd1 vccd1 hold2737/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2748 _25910_/Q vssd1 vssd1 vccd1 vccd1 _23232_/A sky130_fd_sc_hd__clkbuf_4
Xhold2759 _25902_/Q vssd1 vssd1 vccd1 vccd1 hold2759/X sky130_fd_sc_hd__dlygate4sd3_1
X_22930_ _26068_/Q vssd1 vssd1 vccd1 vccd1 _22931_/A sky130_fd_sc_hd__inv_2
XFILLER_0_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22861_ _23010_/A _22861_/B vssd1 vssd1 vccd1 vccd1 _22862_/A sky130_fd_sc_hd__xor2_1
X_24600_ hold2329/X _26263_/Q _24664_/S vssd1 vssd1 vccd1 vccd1 _24600_/X sky130_fd_sc_hd__mux2_1
X_21812_ _21812_/A _21812_/B vssd1 vssd1 vccd1 vccd1 _21812_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25580_ _25878_/CLK _25580_/D vssd1 vssd1 vccd1 vccd1 _25580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22792_ _22792_/A _23104_/B vssd1 vssd1 vccd1 vccd1 _22793_/B sky130_fd_sc_hd__nand2_1
X_24531_ _24531_/A vssd1 vssd1 vccd1 vccd1 _26240_/D sky130_fd_sc_hd__clkbuf_1
X_21743_ _21743_/A _22561_/B vssd1 vssd1 vccd1 vccd1 _21744_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_176_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24462_ _24462_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24463_/A sky130_fd_sc_hd__and2_1
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21674_ _21676_/A _21677_/B vssd1 vssd1 vccd1 vccd1 _21675_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26201_ _26202_/CLK _26201_/D vssd1 vssd1 vccd1 vccd1 _26201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23413_ hold254/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23413_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20625_ _20625_/A _20625_/B vssd1 vssd1 vccd1 vccd1 _20628_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_50_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24393_ _24393_/A vssd1 vssd1 vccd1 vccd1 _26195_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26132_ _26136_/CLK _26132_/D vssd1 vssd1 vccd1 vccd1 _26132_/Q sky130_fd_sc_hd__dfxtp_1
X_23344_ _23344_/A vssd1 vssd1 vccd1 vccd1 _25931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20556_ _21319_/C vssd1 vssd1 vccd1 vccd1 _21322_/B sky130_fd_sc_hd__inv_2
XFILLER_0_22_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26063_ _26064_/CLK _26063_/D vssd1 vssd1 vccd1 vccd1 _26063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23275_ _23275_/A _23275_/B vssd1 vssd1 vccd1 vccd1 _23276_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20487_ _20487_/A _20487_/B _20487_/C vssd1 vssd1 vccd1 vccd1 _20488_/B sky130_fd_sc_hd__nand3_1
X_25014_ _26096_/CLK _25014_/D vssd1 vssd1 vccd1 vccd1 _25014_/Q sky130_fd_sc_hd__dfxtp_1
X_22226_ _22227_/A _22227_/C _23138_/A vssd1 vssd1 vccd1 vccd1 _22226_/X sky130_fd_sc_hd__a21o_1
X_22157_ _22157_/A _22824_/A vssd1 vssd1 vccd1 vccd1 _22168_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21108_ _21108_/A _21108_/B vssd1 vssd1 vccd1 vccd1 _21110_/A sky130_fd_sc_hd__nand2_1
X_22088_ _22561_/A _22088_/B vssd1 vssd1 vccd1 vccd1 _22088_/Y sky130_fd_sc_hd__nand2_1
X_13930_ hold537/X _13929_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold538/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25916_ _26341_/CLK _25916_/D vssd1 vssd1 vccd1 vccd1 _25916_/Q sky130_fd_sc_hd__dfxtp_1
X_21039_ _26305_/Q _20731_/X hold482/X vssd1 vssd1 vccd1 vccd1 _21042_/B sky130_fd_sc_hd__a21oi_1
X_25847_ _26208_/CLK _25847_/D vssd1 vssd1 vccd1 vccd1 _25847_/Q sky130_fd_sc_hd__dfxtp_4
X_13861_ hold807/X _13860_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold808/A sky130_fd_sc_hd__a21oi_1
X_15600_ _15621_/A _16532_/B vssd1 vssd1 vccd1 vccd1 _15603_/A sky130_fd_sc_hd__nor2_1
X_12812_ _12746_/X _12810_/X _14910_/B _12811_/X vssd1 vssd1 vccd1 vccd1 _12812_/X
+ sky130_fd_sc_hd__o211a_1
X_16580_ _16580_/A _16596_/A vssd1 vssd1 vccd1 vccd1 _16581_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25778_ _25779_/CLK _25778_/D vssd1 vssd1 vccd1 vccd1 _25778_/Q sky130_fd_sc_hd__dfxtp_1
X_13792_ _13880_/A hold733/X vssd1 vssd1 vccd1 vccd1 hold734/A sky130_fd_sc_hd__nand2_1
X_15531_ _15531_/A _15531_/B vssd1 vssd1 vccd1 vccd1 _15550_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_69_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _12723_/X _12724_/X _12726_/Y _12730_/Y _14260_/A vssd1 vssd1 vccd1 vccd1
+ _12743_/X sky130_fd_sc_hd__a41o_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24729_ _24729_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24730_/A sky130_fd_sc_hd__and2_1
XFILLER_0_9_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ _18248_/Y _17528_/X _18249_/X vssd1 vssd1 vccd1 vccd1 _18251_/A sky130_fd_sc_hd__a21o_1
X_15462_ _15463_/B _15463_/A vssd1 vssd1 vccd1 vccd1 _15462_/X sky130_fd_sc_hd__or2_1
X_12674_ _12674_/A _12674_/B vssd1 vssd1 vccd1 vccd1 _12676_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_167_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _17199_/X _23187_/B _17200_/X vssd1 vssd1 vccd1 vccd1 _17202_/A sky130_fd_sc_hd__a21o_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14413_ _14413_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14413_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_65_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18181_ _18252_/A _18181_/B vssd1 vssd1 vccd1 vccd1 _18181_/Y sky130_fd_sc_hd__nand2_1
X_15393_ _15391_/X _15392_/Y _15090_/X vssd1 vssd1 vccd1 vccd1 _25451_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17132_ _19729_/A _17132_/B vssd1 vssd1 vccd1 vccd1 _17548_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_108_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14344_ _14344_/A hold338/X vssd1 vssd1 vccd1 vccd1 hold339/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17063_ _17063_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17063_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14275_ _14277_/B _14277_/C vssd1 vssd1 vccd1 vccd1 _14275_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_123_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16014_ _16014_/A _16027_/A vssd1 vssd1 vccd1 vccd1 _16016_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_122_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13226_ _13207_/X _13224_/X _13192_/X _13225_/X vssd1 vssd1 vccd1 vccd1 _13226_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _13109_/X _13155_/X _13096_/X _13156_/X vssd1 vssd1 vccd1 vccd1 _13157_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965_ _17965_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _17965_/Y sky130_fd_sc_hd__nand2_1
X_13088_ _26278_/Q _25647_/Q vssd1 vssd1 vccd1 vccd1 _14494_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_97_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19704_ _19720_/B _19793_/B vssd1 vssd1 vccd1 vccd1 _19706_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16916_ _23053_/B _13468_/X _16774_/Y vssd1 vssd1 vccd1 vccd1 _16916_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17896_ _17896_/A _17896_/B _17896_/C vssd1 vssd1 vccd1 vccd1 _22133_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_189_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19635_ _19635_/A _19635_/B vssd1 vssd1 vccd1 vccd1 _19635_/Y sky130_fd_sc_hd__nand2_1
X_16847_ _16848_/B _16848_/A vssd1 vssd1 vccd1 vccd1 _16847_/X sky130_fd_sc_hd__or2_1
XFILLER_0_189_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19566_ _19564_/X _19565_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19566_/Y sky130_fd_sc_hd__a21oi_1
X_16778_ _16776_/Y _15290_/A _16777_/Y vssd1 vssd1 vccd1 vccd1 _16778_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18517_ _18517_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18517_/Y sky130_fd_sc_hd__nand2_1
X_15729_ _15729_/A vssd1 vssd1 vccd1 vccd1 _16946_/A sky130_fd_sc_hd__inv_2
XFILLER_0_158_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19497_ _19487_/X _19495_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19497_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18448_ _18954_/A _25748_/Q vssd1 vssd1 vccd1 vccd1 _18450_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_173_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18379_ _21981_/B _25617_/Q vssd1 vssd1 vccd1 vccd1 _18381_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_172_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20410_ _20410_/A _20410_/B vssd1 vssd1 vccd1 vccd1 _21531_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21390_ _26320_/Q _21228_/X hold748/X vssd1 vssd1 vccd1 vccd1 _21393_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20341_ _26285_/Q _20078_/X hold389/X vssd1 vssd1 vccd1 vccd1 _20344_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23060_ _23188_/A _23060_/B vssd1 vssd1 vccd1 vccd1 _23060_/X sky130_fd_sc_hd__or2_1
X_20272_ _20272_/A _22297_/B vssd1 vssd1 vccd1 vccd1 _20273_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22011_ _22011_/A _22011_/B vssd1 vssd1 vccd1 vccd1 _22012_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2501 _12672_/X vssd1 vssd1 vccd1 vccd1 _12673_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2512 _26105_/Q vssd1 vssd1 vccd1 vccd1 hold2512/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2523 _26081_/Q vssd1 vssd1 vccd1 vccd1 hold2523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2534 _26083_/Q vssd1 vssd1 vccd1 vccd1 hold2534/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1800 _23956_/X vssd1 vssd1 vccd1 vccd1 _23957_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2545 _25682_/Q vssd1 vssd1 vccd1 vccd1 _13295_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1811 _25839_/Q vssd1 vssd1 vccd1 vccd1 _21793_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2556 _24489_/X vssd1 vssd1 vccd1 vccd1 _24490_/A sky130_fd_sc_hd__dlygate4sd3_1
X_23962_ hold2183/X _26056_/Q _24001_/S vssd1 vssd1 vccd1 vccd1 _23962_/X sky130_fd_sc_hd__mux2_1
Xhold1822 _14902_/Y vssd1 vssd1 vccd1 vccd1 _14905_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2567 _26249_/Q vssd1 vssd1 vccd1 vccd1 hold2567/X sky130_fd_sc_hd__buf_1
Xhold1833 _24089_/X vssd1 vssd1 vccd1 vccd1 _24090_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2578 _26299_/Q vssd1 vssd1 vccd1 vccd1 hold2578/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1844 _21863_/Y vssd1 vssd1 vccd1 vccd1 _25841_/D sky130_fd_sc_hd__dlygate4sd3_1
X_25701_ _26335_/CLK _25701_/D vssd1 vssd1 vccd1 vccd1 _25701_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2589 _26316_/Q vssd1 vssd1 vccd1 vccd1 hold2589/X sky130_fd_sc_hd__dlygate4sd3_1
X_22913_ _26067_/Q vssd1 vssd1 vccd1 vccd1 _22914_/A sky130_fd_sc_hd__inv_2
Xhold1855 _21966_/Y vssd1 vssd1 vccd1 vccd1 _25844_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1866 _25631_/Q vssd1 vssd1 vccd1 vccd1 _17553_/B sky130_fd_sc_hd__dlygate4sd3_1
X_23893_ _23893_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23894_/A sky130_fd_sc_hd__and2_1
Xhold1877 _17533_/Y vssd1 vssd1 vccd1 vccd1 _25628_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1888 _25999_/Q vssd1 vssd1 vccd1 vccd1 _14859_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1899 _25705_/Q vssd1 vssd1 vccd1 vccd1 _19057_/B sky130_fd_sc_hd__dlygate4sd3_1
X_25632_ _25716_/CLK _25632_/D vssd1 vssd1 vccd1 vccd1 _25632_/Q sky130_fd_sc_hd__dfxtp_4
X_22844_ _22844_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22844_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_116_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25563_ _26066_/CLK _25563_/D vssd1 vssd1 vccd1 vccd1 _25563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22775_ _22775_/A _23088_/B vssd1 vssd1 vccd1 vccd1 _22776_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_93_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24514_ hold2683/X hold2380/X _24587_/S vssd1 vssd1 vccd1 vccd1 _24515_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21726_ _21721_/X _14270_/A _21722_/Y _14703_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _21727_/A sky130_fd_sc_hd__a32o_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25494_ _25495_/CLK hold765/X vssd1 vssd1 vccd1 vccd1 hold763/A sky130_fd_sc_hd__dfxtp_1
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24445_ _24445_/A vssd1 vssd1 vccd1 vccd1 _26212_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21657_ _21708_/B _21661_/B vssd1 vssd1 vccd1 vccd1 _21659_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_164_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20608_ _21612_/A vssd1 vssd1 vccd1 vccd1 _21611_/A sky130_fd_sc_hd__inv_2
X_24376_ _24560_/A vssd1 vssd1 vccd1 vccd1 _24465_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21588_ _21588_/A _22902_/B vssd1 vssd1 vccd1 vccd1 _21588_/Y sky130_fd_sc_hd__nand2_1
X_26115_ _26116_/CLK _26115_/D vssd1 vssd1 vccd1 vccd1 _26115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23327_ _23327_/A vssd1 vssd1 vccd1 vccd1 _23330_/B sky130_fd_sc_hd__inv_2
X_20539_ _20538_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20539_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_62_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26046_ _26046_/CLK _26046_/D vssd1 vssd1 vccd1 vccd1 _26046_/Q sky130_fd_sc_hd__dfxtp_1
X_14060_ _26307_/Q _13988_/X _13981_/X _14059_/Y vssd1 vssd1 vccd1 vccd1 _14061_/B
+ sky130_fd_sc_hd__a22o_1
X_23258_ _23258_/A _23278_/B vssd1 vssd1 vccd1 vccd1 _23267_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_120_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13011_ _17557_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13011_/X sky130_fd_sc_hd__or2_1
X_22209_ _18553_/A _25817_/Q _22207_/Y _22208_/Y vssd1 vssd1 vccd1 vccd1 _22210_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23189_ _15811_/B _22893_/A _22829_/A vssd1 vssd1 vccd1 vccd1 _23189_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14962_ _14962_/A _14962_/B vssd1 vssd1 vccd1 vccd1 _14962_/Y sky130_fd_sc_hd__nand2_1
X_17750_ _17750_/A _17750_/B vssd1 vssd1 vccd1 vccd1 _17924_/B sky130_fd_sc_hd__nand2_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
X_16701_ _16858_/A _22423_/B vssd1 vssd1 vccd1 vccd1 _16701_/Y sky130_fd_sc_hd__nand2_1
X_13913_ _25781_/Q vssd1 vssd1 vccd1 vccd1 _18124_/B sky130_fd_sc_hd__inv_2
X_14893_ _14893_/A _14893_/B vssd1 vssd1 vccd1 vccd1 _22387_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17681_ _17692_/A _17691_/B _17692_/B vssd1 vssd1 vccd1 vccd1 _17723_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19420_ _19421_/B _19421_/A vssd1 vssd1 vccd1 vccd1 _19420_/X sky130_fd_sc_hd__or2_1
X_16632_ _16649_/B _16610_/B _16631_/Y vssd1 vssd1 vccd1 vccd1 _16634_/A sky130_fd_sc_hd__o21ai_1
X_13844_ _13880_/A hold780/X vssd1 vssd1 vccd1 vccd1 hold781/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19351_ _19349_/X _19350_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19351_/Y sky130_fd_sc_hd__a21oi_1
X_16563_ _16563_/A vssd1 vssd1 vccd1 vccd1 _16575_/A sky130_fd_sc_hd__inv_2
X_13775_ _25759_/Q vssd1 vssd1 vccd1 vccd1 _18673_/B sky130_fd_sc_hd__inv_2
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18302_ _25869_/Q _21843_/A vssd1 vssd1 vccd1 vccd1 _18310_/A sky130_fd_sc_hd__or2_2
X_15514_ _15514_/A vssd1 vssd1 vccd1 vccd1 _16862_/A sky130_fd_sc_hd__inv_2
X_12726_ _14287_/A _12726_/B vssd1 vssd1 vccd1 vccd1 _12726_/Y sky130_fd_sc_hd__nand2_1
X_16494_ _16489_/B _16393_/B _16491_/X _16493_/X vssd1 vssd1 vccd1 vccd1 _16495_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19282_ _19274_/X _19281_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19282_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_183_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15445_ _15427_/A _15404_/A _15426_/A vssd1 vssd1 vccd1 vccd1 _15446_/B sky130_fd_sc_hd__a21oi_1
X_18233_ _18231_/Y _18232_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25656_/D sky130_fd_sc_hd__a21oi_1
X_12657_ _12657_/A _24836_/B _12664_/B vssd1 vssd1 vccd1 vccd1 _12658_/A sky130_fd_sc_hd__and3_1
XFILLER_0_38_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15376_ _15331_/X _15406_/B _15406_/C _15375_/X vssd1 vssd1 vccd1 vccd1 _15378_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_154_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18164_ _20936_/B _19388_/A vssd1 vssd1 vccd1 vccd1 _18165_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_108_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12588_ _12591_/A _24836_/B _12588_/C vssd1 vssd1 vccd1 vccd1 _12589_/A sky130_fd_sc_hd__and3_1
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17115_ _20547_/B _25852_/Q _25788_/Q vssd1 vssd1 vccd1 vccd1 _17116_/B sky130_fd_sc_hd__mux2_2
X_14327_ _14325_/Y hold333/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold334/A sky130_fd_sc_hd__a21oi_1
X_18095_ _18445_/A _18101_/B vssd1 vssd1 vccd1 vccd1 _18097_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold407 hold407/A vssd1 vssd1 vccd1 vccd1 hold407/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold418 hold418/A vssd1 vssd1 vccd1 vccd1 hold418/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17046_ _17044_/X _23187_/B _17045_/X vssd1 vssd1 vccd1 vccd1 _17047_/A sky130_fd_sc_hd__a21o_1
Xhold429 hold429/A vssd1 vssd1 vccd1 vccd1 hold429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14258_ _14264_/A _14258_/B vssd1 vssd1 vccd1 vccd1 _14258_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13209_ _26299_/Q _19345_/A vssd1 vssd1 vccd1 vccd1 _14560_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_111_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14189_ _25825_/Q vssd1 vssd1 vccd1 vccd1 _18714_/B sky130_fd_sc_hd__inv_2
XFILLER_0_21_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _18997_/A _18997_/B vssd1 vssd1 vccd1 vccd1 _18997_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_139_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 _25041_/Q vssd1 vssd1 vccd1 vccd1 _17479_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1118 _16880_/Y vssd1 vssd1 vccd1 vccd1 _25565_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17948_ _19317_/A vssd1 vssd1 vccd1 vccd1 _21764_/B sky130_fd_sc_hd__inv_2
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1129 _25108_/Q vssd1 vssd1 vccd1 vccd1 _18880_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17879_ _17881_/A vssd1 vssd1 vccd1 vccd1 _17880_/A sky130_fd_sc_hd__inv_2
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19618_ _20098_/A _19616_/Y _20102_/C vssd1 vssd1 vccd1 vccd1 _19706_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_136_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20890_ _20890_/A _20890_/B vssd1 vssd1 vccd1 vccd1 _21467_/B sky130_fd_sc_hd__nand2_4
X_19549_ _19565_/B _19635_/B vssd1 vssd1 vccd1 vccd1 _19551_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22560_ _22551_/Y _22559_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22560_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_152_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21511_ _21562_/A _21515_/A vssd1 vssd1 vccd1 vccd1 _21513_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_91_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22491_ _19802_/A _22490_/A _22490_/Y vssd1 vssd1 vccd1 vccd1 _22493_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_173_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24230_ _24230_/A vssd1 vssd1 vccd1 vccd1 _26142_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_173_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21442_ _21442_/A _21442_/B vssd1 vssd1 vccd1 vccd1 _21443_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_146_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24161_ _24161_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24162_/A sky130_fd_sc_hd__and2_1
X_21373_ _21373_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21378_/A sky130_fd_sc_hd__nand2_1
X_23112_ _23111_/A _22849_/X _23111_/B vssd1 vssd1 vccd1 vccd1 _23113_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20324_ _20324_/A _25885_/Q vssd1 vssd1 vccd1 vccd1 _20330_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24092_ hold2270/X hold2267/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24093_/A sky130_fd_sc_hd__mux2_1
Xhold930 hold930/A vssd1 vssd1 vccd1 vccd1 hold930/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold941 hold941/A vssd1 vssd1 vccd1 vccd1 hold941/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold952 hold952/A vssd1 vssd1 vccd1 vccd1 hold952/X sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_209_clk _26093_/CLK vssd1 vssd1 vccd1 vccd1 _25587_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold963 hold963/A vssd1 vssd1 vccd1 vccd1 hold963/X sky130_fd_sc_hd__dlygate4sd3_1
X_23043_ _23043_/A _23187_/B vssd1 vssd1 vccd1 vccd1 _23043_/Y sky130_fd_sc_hd__nand2_1
X_20255_ _20255_/A _20255_/B vssd1 vssd1 vccd1 vccd1 _21114_/C sky130_fd_sc_hd__nand2_4
Xhold974 hold974/A vssd1 vssd1 vccd1 vccd1 hold974/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 hold985/A vssd1 vssd1 vccd1 vccd1 hold985/X sky130_fd_sc_hd__buf_1
Xhold996 hold996/A vssd1 vssd1 vccd1 vccd1 hold996/X sky130_fd_sc_hd__dlygate4sd3_1
X_20186_ _20186_/A _20978_/C vssd1 vssd1 vccd1 vccd1 _20188_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_122_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2320 _25934_/Q vssd1 vssd1 vccd1 vccd1 _23354_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2331 _26191_/Q vssd1 vssd1 vccd1 vccd1 hold2331/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2342 _24966_/Q vssd1 vssd1 vccd1 vccd1 _12562_/A sky130_fd_sc_hd__buf_1
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24994_ _25422_/CLK _24994_/D vssd1 vssd1 vccd1 vccd1 _24994_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2353 _26199_/Q vssd1 vssd1 vccd1 vccd1 hold2353/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2364 _25416_/Q vssd1 vssd1 vccd1 vccd1 _14931_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2375 _15039_/Y vssd1 vssd1 vccd1 vccd1 hold2375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1630 _25588_/Q vssd1 vssd1 vccd1 vccd1 _17112_/B sky130_fd_sc_hd__clkbuf_2
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1641 _25810_/Q vssd1 vssd1 vccd1 vccd1 _21262_/B sky130_fd_sc_hd__dlygate4sd3_1
X_23945_ _23945_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23946_/A sky130_fd_sc_hd__and2_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2386 _25659_/Q vssd1 vssd1 vccd1 vccd1 _13152_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1652 _21607_/Y vssd1 vssd1 vccd1 vccd1 _25830_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2397 _26143_/Q vssd1 vssd1 vccd1 vccd1 hold2397/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1663 _25876_/Q vssd1 vssd1 vccd1 vccd1 _22789_/B sky130_fd_sc_hd__buf_1
XFILLER_0_93_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1674 _25586_/Q vssd1 vssd1 vccd1 vccd1 _17080_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1685 _25798_/Q vssd1 vssd1 vccd1 vccd1 _20933_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1696 _25886_/Q vssd1 vssd1 vccd1 vccd1 _22954_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23876_ _23876_/A vssd1 vssd1 vccd1 vccd1 _26029_/D sky130_fd_sc_hd__clkbuf_1
X_25615_ _26249_/CLK _25615_/D vssd1 vssd1 vccd1 vccd1 _25615_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22827_ _22827_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22827_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_39_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25546_ _26053_/CLK _25546_/D vssd1 vssd1 vccd1 vccd1 _25546_/Q sky130_fd_sc_hd__dfxtp_1
X_13560_ hold447/X _13558_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold448/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22758_ _23071_/B _22758_/B vssd1 vssd1 vccd1 vccd1 _22760_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12511_ hold410/A _24994_/Q hold997/A hold837/A vssd1 vssd1 vccd1 vccd1 _12514_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_48_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21709_ _21709_/A _21709_/B vssd1 vssd1 vccd1 vccd1 _21710_/C sky130_fd_sc_hd__nand2_1
X_25477_ _25913_/CLK hold694/X vssd1 vssd1 vccd1 vccd1 hold692/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13491_ hold414/X _13490_/Y _12558_/B vssd1 vssd1 vccd1 vccd1 hold415/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22689_ _22937_/A _22689_/B vssd1 vssd1 vccd1 vccd1 _22689_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15230_ _15230_/A vssd1 vssd1 vccd1 vccd1 _16754_/A sky130_fd_sc_hd__inv_2
X_24428_ _24428_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24429_/A sky130_fd_sc_hd__and2_1
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15161_ _15161_/A _15161_/B vssd1 vssd1 vccd1 vccd1 _15184_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_152_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24359_ _24835_/S vssd1 vssd1 vccd1 vccd1 _24433_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14112_ _14118_/A hold587/X vssd1 vssd1 vccd1 vccd1 hold588/A sky130_fd_sc_hd__nand2_1
XFILLER_0_132_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15092_ _15092_/A vssd1 vssd1 vccd1 vccd1 _15100_/B sky130_fd_sc_hd__inv_2
XFILLER_0_120_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26029_ _26032_/CLK _26029_/D vssd1 vssd1 vccd1 vccd1 _26029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14043_ _14061_/A _14043_/B vssd1 vssd1 vccd1 vccd1 _14043_/Y sky130_fd_sc_hd__nand2_1
X_18920_ _19026_/A _18920_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18920_/X sky130_fd_sc_hd__and3_1
X_18851_ _18851_/A _25832_/Q _18851_/C vssd1 vssd1 vccd1 vccd1 _20758_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_101_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17802_ _20396_/B _22078_/A vssd1 vssd1 vccd1 vccd1 _20389_/A sky130_fd_sc_hd__nand2_4
X_18782_ _18986_/A _19560_/A vssd1 vssd1 vccd1 vccd1 _18782_/Y sky130_fd_sc_hd__nand2_1
X_15994_ _22115_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _15996_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17733_ _17733_/A _17733_/B vssd1 vssd1 vccd1 vccd1 _17771_/C sky130_fd_sc_hd__nand2_2
X_14945_ _14945_/A _14945_/B vssd1 vssd1 vccd1 vccd1 _14946_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17664_ _17665_/B _17665_/A vssd1 vssd1 vccd1 vccd1 _20026_/A sky130_fd_sc_hd__or2_2
X_14876_ _14882_/B _22344_/A vssd1 vssd1 vccd1 vccd1 _22343_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19403_ _20964_/A _21972_/B _25608_/Q vssd1 vssd1 vccd1 vccd1 _20969_/C sky130_fd_sc_hd__nand3_1
X_16615_ hold887/X vssd1 vssd1 vccd1 vccd1 _24952_/A sky130_fd_sc_hd__inv_2
XFILLER_0_98_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13827_ _25767_/Q vssd1 vssd1 vccd1 vccd1 _18833_/B sky130_fd_sc_hd__inv_2
XFILLER_0_58_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17595_ _17624_/A _17595_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _17595_/X sky130_fd_sc_hd__and3_1
XFILLER_0_134_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19334_ _19350_/B _19421_/B vssd1 vssd1 vccd1 vccd1 _19336_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_187_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16546_ _16537_/B _16533_/Y _16525_/Y _16542_/A _16535_/B vssd1 vssd1 vccd1 vccd1
+ _16554_/B sky130_fd_sc_hd__o221a_1
XFILLER_0_134_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13758_ _13823_/A _13758_/B vssd1 vssd1 vccd1 vccd1 _13758_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12709_ _24989_/Q _24988_/Q vssd1 vssd1 vccd1 vccd1 _12713_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_39_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19265_ _19265_/A _19994_/B _19265_/C vssd1 vssd1 vccd1 vccd1 _19265_/X sky130_fd_sc_hd__and3_1
X_16477_ _16477_/A _16483_/B vssd1 vssd1 vccd1 vccd1 _16478_/A sky130_fd_sc_hd__nand2_1
X_13689_ _18387_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13689_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_156_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18216_ _20994_/B _19416_/A vssd1 vssd1 vccd1 vccd1 _18217_/B sky130_fd_sc_hd__nand2_1
X_15428_ _15414_/A _15403_/Y _15404_/A vssd1 vssd1 vccd1 vccd1 _15430_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_142_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19196_ _19191_/X _18879_/X _19195_/X vssd1 vssd1 vccd1 vccd1 _19198_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_171_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15359_ _15331_/X _15406_/B _15342_/B vssd1 vssd1 vccd1 vccd1 _15361_/A sky130_fd_sc_hd__a21o_1
X_18147_ _18252_/A _18147_/B vssd1 vssd1 vccd1 vccd1 _18147_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_81_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold204 hold204/A vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold215 hold215/A vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18078_ _22248_/B _25598_/Q vssd1 vssd1 vccd1 vccd1 _18080_/A sky130_fd_sc_hd__nand2_1
Xhold226 hold226/A vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold237 hold237/A vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 hold248/A vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 hold259/A vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
X_17029_ _17393_/A _17029_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17029_/X sky130_fd_sc_hd__and3_1
XFILLER_0_106_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20040_ _20040_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _20040_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21991_ _25845_/Q _25781_/Q vssd1 vssd1 vccd1 vccd1 _21992_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23730_ hold2161/X hold2244/X _23754_/S vssd1 vssd1 vccd1 vccd1 _23731_/A sky130_fd_sc_hd__mux2_1
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20942_ _20944_/B vssd1 vssd1 vccd1 vccd1 _20943_/B sky130_fd_sc_hd__inv_2
XFILLER_0_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23661_ _23661_/A vssd1 vssd1 vccd1 vccd1 _25959_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20873_ _20873_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _20878_/A sky130_fd_sc_hd__nand2_1
X_25400_ _25425_/CLK _25400_/D vssd1 vssd1 vccd1 vccd1 _25400_/Q sky130_fd_sc_hd__dfxtp_1
X_22612_ _22937_/A _22612_/B vssd1 vssd1 vccd1 vccd1 _22612_/Y sky130_fd_sc_hd__nand2_1
X_23592_ _23592_/A _24745_/A _23592_/C vssd1 vssd1 vccd1 vccd1 _23593_/B sky130_fd_sc_hd__and3_1
XFILLER_0_113_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25331_ _26283_/CLK hold91/X vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22543_ _22544_/B _22544_/A vssd1 vssd1 vccd1 vccd1 _22545_/A sky130_fd_sc_hd__or2_1
XFILLER_0_107_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25262_ _26219_/CLK hold157/X vssd1 vssd1 vccd1 vccd1 hold155/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22474_ _23152_/A _22474_/B vssd1 vssd1 vccd1 vccd1 _22475_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24213_ hold2001/X _26137_/Q _24279_/S vssd1 vssd1 vccd1 vccd1 _24213_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21425_ _21636_/A _21425_/B _21424_/X vssd1 vssd1 vccd1 vccd1 _21426_/B sky130_fd_sc_hd__or3b_1
X_25193_ _26251_/CLK hold727/X vssd1 vssd1 vccd1 vccd1 hold725/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24144_ _24144_/A vssd1 vssd1 vccd1 vccd1 _26114_/D sky130_fd_sc_hd__clkbuf_1
X_21356_ _21356_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21361_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20307_ _20660_/A _20307_/B vssd1 vssd1 vccd1 vccd1 _20307_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_130_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24075_ _24075_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24076_/A sky130_fd_sc_hd__and2_1
Xhold760 hold760/A vssd1 vssd1 vccd1 vccd1 hold760/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21287_ _21287_/A _21508_/B vssd1 vssd1 vccd1 vccd1 _21287_/Y sky130_fd_sc_hd__nand2_1
Xhold771 hold771/A vssd1 vssd1 vccd1 vccd1 hold771/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 hold782/A vssd1 vssd1 vccd1 vccd1 hold782/X sky130_fd_sc_hd__dlygate4sd3_1
X_23026_ _23026_/A _23026_/B vssd1 vssd1 vccd1 vccd1 _23027_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_102_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold793 hold793/A vssd1 vssd1 vccd1 vccd1 hold793/X sky130_fd_sc_hd__dlygate4sd3_1
X_20238_ _20238_/A _25883_/Q vssd1 vssd1 vccd1 vccd1 _20244_/A sky130_fd_sc_hd__nand2_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20169_ _20171_/B vssd1 vssd1 vccd1 vccd1 _20170_/B sky130_fd_sc_hd__inv_2
Xhold2150 _25937_/Q vssd1 vssd1 vccd1 vccd1 _23369_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2161 _25981_/Q vssd1 vssd1 vccd1 vccd1 hold2161/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_189_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2172 _25926_/Q vssd1 vssd1 vccd1 vccd1 _23316_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2183 _26055_/Q vssd1 vssd1 vccd1 vccd1 hold2183/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _12930_/X _12989_/X _12917_/X _12990_/X vssd1 vssd1 vccd1 vccd1 _12991_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2194 _25425_/Q vssd1 vssd1 vccd1 vccd1 _15006_/B sky130_fd_sc_hd__dlygate4sd3_1
X_24977_ _25420_/CLK _24977_/D vssd1 vssd1 vccd1 vccd1 _24977_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1460 _13334_/X vssd1 vssd1 vccd1 vccd1 _25107_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1471 _25398_/Q vssd1 vssd1 vccd1 vccd1 _14786_/B sky130_fd_sc_hd__clkbuf_2
X_14730_ _14730_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14730_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1482 _16779_/Y vssd1 vssd1 vccd1 vccd1 _25550_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23928_ _24047_/S vssd1 vssd1 vccd1 vccd1 _24001_/S sky130_fd_sc_hd__buf_12
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1493 _25101_/Q vssd1 vssd1 vccd1 vccd1 _18739_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _14688_/A hold392/X vssd1 vssd1 vccd1 vccd1 hold393/A sky130_fd_sc_hd__nand2_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23859_ hold1907/X _26024_/Q _23907_/S vssd1 vssd1 vccd1 vccd1 _23859_/X sky130_fd_sc_hd__mux2_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16400_ _16676_/A _15422_/A _16399_/Y vssd1 vssd1 vccd1 vccd1 _16402_/A sky130_fd_sc_hd__o21a_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13612_ _14262_/B vssd1 vssd1 vccd1 vccd1 _13612_/X sky130_fd_sc_hd__buf_12
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _14589_/Y hold186/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold187/A sky130_fd_sc_hd__a21oi_1
X_17380_ _19532_/A _17380_/B vssd1 vssd1 vccd1 vccd1 _17615_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_156_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16331_ _16331_/A _16331_/B vssd1 vssd1 vccd1 vccd1 _16332_/B sky130_fd_sc_hd__and2_1
XFILLER_0_137_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13543_ _25722_/Q vssd1 vssd1 vccd1 vccd1 _17895_/B sky130_fd_sc_hd__inv_2
XFILLER_0_94_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25529_ _25533_/CLK hold911/X vssd1 vssd1 vccd1 vccd1 hold910/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16262_ _16262_/A _16262_/B vssd1 vssd1 vccd1 vccd1 _16263_/B sky130_fd_sc_hd__nand2_1
X_19050_ _19186_/A _19050_/B vssd1 vssd1 vccd1 vccd1 _19050_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13474_ _13522_/A hold497/X vssd1 vssd1 vccd1 vccd1 hold498/A sky130_fd_sc_hd__nand2_1
XFILLER_0_137_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15213_ _16747_/A _15213_/B vssd1 vssd1 vccd1 vccd1 _15214_/B sky130_fd_sc_hd__and2_1
XFILLER_0_35_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18001_ _18528_/A _25731_/Q vssd1 vssd1 vccd1 vccd1 _18003_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_113_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16193_ _16195_/B _16195_/A vssd1 vssd1 vccd1 vccd1 _16194_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_180_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15144_ _16719_/A _15144_/B vssd1 vssd1 vccd1 vccd1 _15145_/B sky130_fd_sc_hd__and2_1
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15075_ _15076_/B _15076_/A vssd1 vssd1 vccd1 vccd1 _15077_/A sky130_fd_sc_hd__or2_1
XFILLER_0_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19952_ _19947_/X _19951_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19952_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14026_ _14118_/A hold437/X vssd1 vssd1 vccd1 vccd1 hold438/A sky130_fd_sc_hd__nand2_1
X_18903_ _18986_/A _19644_/A vssd1 vssd1 vccd1 vccd1 _18903_/Y sky130_fd_sc_hd__nand2_1
X_19883_ _19883_/A _19980_/B _19883_/C vssd1 vssd1 vccd1 vccd1 _19883_/X sky130_fd_sc_hd__and3_1
X_18834_ _18834_/A _18834_/B _18834_/C vssd1 vssd1 vccd1 vccd1 _22566_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18765_ _22488_/B _25636_/Q vssd1 vssd1 vccd1 vccd1 _18767_/A sky130_fd_sc_hd__nand2_1
X_15977_ _15978_/B _15978_/A vssd1 vssd1 vccd1 vccd1 _15979_/A sky130_fd_sc_hd__or2_1
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17716_ _17726_/A _17725_/B _17726_/C vssd1 vssd1 vccd1 vccd1 _17724_/A sky130_fd_sc_hd__nand3_1
X_14928_ _15464_/A vssd1 vssd1 vccd1 vccd1 _14928_/X sky130_fd_sc_hd__buf_6
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18696_ _18696_/A _20438_/A vssd1 vssd1 vccd1 vccd1 _18988_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_37_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17647_ _17645_/X _17528_/X _17646_/X vssd1 vssd1 vccd1 vccd1 _17648_/A sky130_fd_sc_hd__a21o_1
X_14859_ _14893_/A _14859_/B vssd1 vssd1 vccd1 vccd1 _22293_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_148_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17578_ _17578_/A _17578_/B vssd1 vssd1 vccd1 vccd1 _17578_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19317_ _19317_/A _20780_/B vssd1 vssd1 vccd1 vccd1 _19317_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16529_ _16529_/A _16686_/B _16537_/A vssd1 vssd1 vccd1 vccd1 _16529_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19248_ _19248_/A _19248_/B vssd1 vssd1 vccd1 vccd1 _19248_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_116_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19179_ _20389_/A _22076_/B _25592_/Q vssd1 vssd1 vccd1 vccd1 _20394_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21210_ _21210_/A _21981_/B vssd1 vssd1 vccd1 vccd1 _21211_/A sky130_fd_sc_hd__nand2_1
X_22190_ _25788_/Q _22190_/B vssd1 vssd1 vccd1 vccd1 _22190_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21141_ _21141_/A _21141_/B _21141_/C vssd1 vssd1 vccd1 vccd1 _21145_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21072_ _21235_/A _21072_/B vssd1 vssd1 vccd1 vccd1 _21072_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24900_ _15844_/B _15855_/B _24945_/S vssd1 vssd1 vccd1 vccd1 _24900_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20023_ _20023_/A _20023_/B vssd1 vssd1 vccd1 vccd1 _20024_/B sky130_fd_sc_hd__nand2_1
X_25880_ _25901_/CLK _25880_/D vssd1 vssd1 vccd1 vccd1 _25880_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_67_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24831_ _24831_/A vssd1 vssd1 vccd1 vccd1 _26338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24762_ _24762_/A vssd1 vssd1 vccd1 vccd1 _26315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21974_ _21974_/A _21974_/B vssd1 vssd1 vccd1 vccd1 _21974_/Y sky130_fd_sc_hd__nand2_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23713_ _23713_/A vssd1 vssd1 vccd1 vccd1 _25976_/D sky130_fd_sc_hd__clkbuf_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20925_ _20925_/A _20925_/B vssd1 vssd1 vccd1 vccd1 _20926_/A sky130_fd_sc_hd__nand2_1
X_24693_ _24693_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24694_/A sky130_fd_sc_hd__and2_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23644_ hold2118/X hold2086/X _23677_/S vssd1 vssd1 vccd1 vccd1 _23645_/A sky130_fd_sc_hd__mux2_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20856_ _20856_/A _20856_/B vssd1 vssd1 vccd1 vccd1 _20860_/A sky130_fd_sc_hd__nand2_1
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23575_ _24922_/S hold350/A _23574_/X vssd1 vssd1 vccd1 vccd1 _23575_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_181_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20787_ _20786_/B _20787_/B _20787_/C vssd1 vssd1 vccd1 vccd1 _20788_/B sky130_fd_sc_hd__nand3b_2
XFILLER_0_76_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25314_ _26263_/CLK hold55/X vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22526_ _22653_/A _22526_/B vssd1 vssd1 vccd1 vccd1 _22526_/X sky130_fd_sc_hd__or2_1
XFILLER_0_135_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26294_ _26296_/CLK _26294_/D vssd1 vssd1 vccd1 vccd1 _26294_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_134_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25245_ _25709_/CLK hold424/X vssd1 vssd1 vccd1 vccd1 hold422/A sky130_fd_sc_hd__dfxtp_1
X_22457_ _16715_/B _22421_/X _22449_/X _22450_/Y _22456_/X vssd1 vssd1 vccd1 vccd1
+ _22458_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_161_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21408_ _21407_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21408_/X
+ sky130_fd_sc_hd__a211o_1
X_13190_ _13049_/X _14551_/A _13067_/X _19303_/A vssd1 vssd1 vccd1 vccd1 _13190_/X
+ sky130_fd_sc_hd__a22o_1
X_25176_ _25773_/CLK hold502/X vssd1 vssd1 vccd1 vccd1 hold500/A sky130_fd_sc_hd__dfxtp_1
X_22388_ _22386_/X _15839_/B _22387_/Y _14900_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _22389_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_121_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24127_ _24127_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24128_/A sky130_fd_sc_hd__and2_1
XFILLER_0_32_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21339_ _21339_/A _21339_/B vssd1 vssd1 vccd1 vccd1 _21340_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_130_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24058_ _24058_/A vssd1 vssd1 vccd1 vccd1 _26086_/D sky130_fd_sc_hd__clkbuf_1
Xhold590 hold590/A vssd1 vssd1 vccd1 vccd1 hold590/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15900_ _15900_/A _15900_/B vssd1 vssd1 vccd1 vccd1 _15909_/A sky130_fd_sc_hd__nand2_1
X_23009_ _23009_/A _23009_/B vssd1 vssd1 vccd1 vccd1 _23010_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_159_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16880_ _16878_/Y _16879_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16880_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15831_ _15830_/A _15800_/B _15817_/A vssd1 vssd1 vccd1 vccd1 _15831_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ _18612_/A _18550_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18551_/C sky130_fd_sc_hd__nand3_1
X_15762_ _15762_/A _15762_/B vssd1 vssd1 vccd1 vccd1 _15786_/B sky130_fd_sc_hd__nand2_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ _17507_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12974_/X sky130_fd_sc_hd__or2_1
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1290 _25792_/Q vssd1 vssd1 vccd1 vccd1 _20738_/B sky130_fd_sc_hd__buf_1
X_17501_ _17499_/X _17241_/X _17500_/X vssd1 vssd1 vccd1 vccd1 _17502_/A sky130_fd_sc_hd__a21o_1
X_14713_ _14711_/Y _14712_/Y _14646_/X vssd1 vssd1 vccd1 vccd1 _14713_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18481_ _22120_/B _25622_/Q vssd1 vssd1 vccd1 vccd1 _18483_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_185_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15693_ _15693_/A _15693_/B _15693_/C vssd1 vssd1 vccd1 vccd1 _15695_/B sky130_fd_sc_hd__and3_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17432_ _19602_/A _17432_/B vssd1 vssd1 vccd1 vccd1 _17651_/B sky130_fd_sc_hd__xor2_4
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14644_ _14644_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14644_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_68_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17363_ _17393_/A _17363_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17363_/X sky130_fd_sc_hd__and3_1
X_14575_ _14575_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14575_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_172_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19102_ _26213_/Q hold452/X vssd1 vssd1 vccd1 vccd1 _19102_/Y sky130_fd_sc_hd__nand2_1
X_16314_ _16314_/A _16697_/B _16322_/A vssd1 vssd1 vccd1 vccd1 _16314_/Y sky130_fd_sc_hd__nand3_1
X_13526_ _26222_/Q _13426_/X _13468_/X _13525_/Y vssd1 vssd1 vccd1 vccd1 _13527_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17294_ _17556_/A _17637_/A vssd1 vssd1 vccd1 vccd1 _17295_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19033_ _19082_/A _19033_/B _22786_/A vssd1 vssd1 vccd1 vccd1 _19033_/X sky130_fd_sc_hd__and3_1
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16245_ _16245_/A _16245_/B vssd1 vssd1 vccd1 vccd1 _16270_/B sky130_fd_sc_hd__nor2_1
X_13457_ _13522_/A _13455_/X _23629_/B _13456_/X vssd1 vssd1 vccd1 vccd1 _13457_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16176_ _16174_/X hold755/X _16076_/X vssd1 vssd1 vccd1 vccd1 hold756/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13388_ _13315_/X _13386_/X _13300_/X _13387_/X vssd1 vssd1 vccd1 vccd1 _13388_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15127_ _16231_/A vssd1 vssd1 vccd1 vccd1 _16698_/A sky130_fd_sc_hd__buf_6
XFILLER_0_121_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15058_ _15058_/A _15058_/B vssd1 vssd1 vccd1 vccd1 _15059_/B sky130_fd_sc_hd__nand2_1
X_19935_ _26271_/Q _19134_/X hold626/X vssd1 vssd1 vccd1 vccd1 _19936_/C sky130_fd_sc_hd__a21o_1
X_14009_ _25796_/Q vssd1 vssd1 vccd1 vccd1 _18053_/B sky130_fd_sc_hd__inv_2
X_19866_ _19864_/Y _19865_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19866_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18817_ _18981_/A _19031_/A vssd1 vssd1 vccd1 vccd1 _18818_/B sky130_fd_sc_hd__xnor2_1
X_19797_ _19795_/Y _19796_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19797_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18748_ _25891_/Q _22462_/A vssd1 vssd1 vccd1 vccd1 _18756_/A sky130_fd_sc_hd__or2_2
XFILLER_0_78_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18679_ _19026_/A _18679_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18679_/X sky130_fd_sc_hd__and3_1
XFILLER_0_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20710_ _21387_/B vssd1 vssd1 vccd1 vccd1 _21384_/C sky130_fd_sc_hd__inv_2
XFILLER_0_77_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21690_ _21692_/A _21693_/B vssd1 vssd1 vccd1 vccd1 _21691_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_176_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20641_ _20643_/B vssd1 vssd1 vccd1 vccd1 _20642_/B sky130_fd_sc_hd__inv_2
XFILLER_0_175_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23360_ _23360_/A _23360_/B vssd1 vssd1 vccd1 vccd1 _23366_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_184_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20572_ _21322_/B _21595_/A vssd1 vssd1 vccd1 vccd1 _20574_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22311_ _19289_/A _22310_/A _22310_/Y vssd1 vssd1 vccd1 vccd1 _22313_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23291_ _23289_/X hold856/X _12702_/A vssd1 vssd1 vccd1 vccd1 hold857/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25030_ _26116_/CLK _25030_/D vssd1 vssd1 vccd1 vccd1 _25030_/Q sky130_fd_sc_hd__dfxtp_1
X_22242_ _22242_/A _22888_/B vssd1 vssd1 vccd1 vccd1 _22243_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22173_ _22653_/A _22173_/B vssd1 vssd1 vccd1 vccd1 _22173_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21124_ _21124_/A _21124_/B vssd1 vssd1 vccd1 vccd1 _21125_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25932_ _25939_/CLK _25932_/D vssd1 vssd1 vccd1 vccd1 _25932_/Q sky130_fd_sc_hd__dfxtp_1
X_21055_ _21055_/A _21055_/B vssd1 vssd1 vccd1 vccd1 _21564_/B sky130_fd_sc_hd__nand2_2
X_20006_ _20006_/A _20006_/B vssd1 vssd1 vccd1 vccd1 _20008_/A sky130_fd_sc_hd__nand2_1
X_25863_ _25864_/CLK _25863_/D vssd1 vssd1 vccd1 vccd1 _25863_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_185_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24814_ hold2684/X _26333_/Q _24817_/S vssd1 vssd1 vccd1 vccd1 _24814_/X sky130_fd_sc_hd__mux2_1
X_25794_ _25794_/CLK _25794_/D vssd1 vssd1 vccd1 vccd1 _25794_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24745_ _24745_/A vssd1 vssd1 vccd1 vccd1 _24833_/B sky130_fd_sc_hd__buf_8
X_21957_ _25844_/Q _25780_/Q vssd1 vssd1 vccd1 vccd1 _21958_/B sky130_fd_sc_hd__nor2_2
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ _20908_/A _21904_/B vssd1 vssd1 vccd1 vccd1 _20909_/A sky130_fd_sc_hd__nand2_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12690_ _12700_/B _12713_/B vssd1 vssd1 vccd1 vccd1 _12690_/Y sky130_fd_sc_hd__nand2_1
X_24676_ _24676_/A vssd1 vssd1 vccd1 vccd1 _26287_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21888_ _25842_/Q _25778_/Q vssd1 vssd1 vccd1 vccd1 _21889_/B sky130_fd_sc_hd__nor2_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23627_ _23627_/A vssd1 vssd1 vccd1 vccd1 _25948_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20839_ _21709_/B vssd1 vssd1 vccd1 vccd1 _21708_/B sky130_fd_sc_hd__inv_2
XFILLER_0_166_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14360_ _14358_/Y hold363/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold364/A sky130_fd_sc_hd__a21oi_1
X_23558_ hold173/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23558_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_147_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13311_ _13220_/X _14611_/A _13242_/X _19574_/A vssd1 vssd1 vccd1 vccd1 _13311_/X
+ sky130_fd_sc_hd__a22o_1
X_22509_ _22500_/Y _22508_/Y _23197_/A vssd1 vssd1 vccd1 vccd1 _22509_/X sky130_fd_sc_hd__a21o_1
X_14291_ _14287_/Y hold264/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold265/A sky130_fd_sc_hd__a21oi_1
X_26277_ _26279_/CLK _26277_/D vssd1 vssd1 vccd1 vccd1 _26277_/Q sky130_fd_sc_hd__dfxtp_2
X_23489_ _23486_/Y _23488_/Y _24858_/S vssd1 vssd1 vccd1 vccd1 _23489_/X sky130_fd_sc_hd__mux2_1
X_16030_ _16031_/B _16031_/A vssd1 vssd1 vccd1 vccd1 _16032_/A sky130_fd_sc_hd__or2_1
XFILLER_0_134_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13242_ _13242_/A vssd1 vssd1 vccd1 vccd1 _13242_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25228_ _25678_/CLK hold790/X vssd1 vssd1 vccd1 vccd1 hold789/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13173_ _26165_/Q _13065_/X _13172_/X vssd1 vssd1 vccd1 vccd1 _13173_/X sky130_fd_sc_hd__a21o_1
X_25159_ _25743_/CLK hold418/X vssd1 vssd1 vccd1 vccd1 hold416/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17981_ _22190_/B _25596_/Q vssd1 vssd1 vccd1 vccd1 _17983_/A sky130_fd_sc_hd__nand2_1
X_19720_ _19720_/A _19720_/B vssd1 vssd1 vccd1 vccd1 _19720_/Y sky130_fd_sc_hd__nand2_1
X_16932_ _16932_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16932_/Y sky130_fd_sc_hd__nand2_1
X_19651_ _19643_/X _19650_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19651_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16863_ _16861_/X _16711_/X _16862_/Y _25884_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16864_/A sky130_fd_sc_hd__a32o_1
X_18602_ _18600_/Y _18601_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25674_/D sky130_fd_sc_hd__a21oi_1
X_15814_ _16691_/A _16711_/A vssd1 vssd1 vccd1 vccd1 _15816_/A sky130_fd_sc_hd__nand2_1
X_19582_ _19723_/A _19582_/B vssd1 vssd1 vccd1 vccd1 _19582_/Y sky130_fd_sc_hd__nand2_1
X_16794_ _16935_/A _16799_/B vssd1 vssd1 vccd1 vccd1 _16796_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_172_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18533_ _18738_/A _18878_/A vssd1 vssd1 vccd1 vccd1 _18534_/B sky130_fd_sc_hd__xnor2_1
X_15745_ _15745_/A _16953_/A vssd1 vssd1 vccd1 vccd1 _15746_/B sky130_fd_sc_hd__nor2_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _12891_/X _14416_/A _12909_/X _25622_/Q vssd1 vssd1 vccd1 vccd1 _12957_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18464_ _25877_/Q _22094_/A vssd1 vssd1 vccd1 vccd1 _18472_/A sky130_fd_sc_hd__or2_2
X_15676_ _15662_/A _15658_/A _15657_/B vssd1 vssd1 vccd1 vccd1 _15676_/X sky130_fd_sc_hd__a21o_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _26112_/Q _12748_/X _12887_/X vssd1 vssd1 vccd1 vccd1 _12888_/X sky130_fd_sc_hd__a21o_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _17413_/X _17241_/X _17414_/X vssd1 vssd1 vccd1 vccd1 _17416_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_184_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14627_ _14645_/A hold149/X vssd1 vssd1 vccd1 vccd1 hold150/A sky130_fd_sc_hd__nand2_1
XFILLER_0_157_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18395_ _18395_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18395_/Y sky130_fd_sc_hd__nand2_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17346_ _17467_/A _17346_/B vssd1 vssd1 vccd1 vccd1 _17346_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14558_ _14585_/A hold71/X vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__nand2_1
XFILLER_0_172_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13509_ hold740/X _13508_/Y _12558_/B vssd1 vssd1 vccd1 vccd1 hold741/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17277_ _25642_/Q vssd1 vssd1 vccd1 vccd1 _20829_/B sky130_fd_sc_hd__inv_2
XFILLER_0_71_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14489_ _14525_/A hold80/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__nand2_1
XFILLER_0_126_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19016_ _19014_/Y _19015_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25699_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16228_ _16246_/A _16228_/B vssd1 vssd1 vccd1 vccd1 _16238_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_180_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16159_ _16272_/A vssd1 vssd1 vccd1 vccd1 _16160_/B sky130_fd_sc_hd__inv_2
XFILLER_0_141_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2705 _26270_/Q vssd1 vssd1 vccd1 vccd1 hold2705/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2716 _26340_/Q vssd1 vssd1 vccd1 vccd1 hold2716/X sky130_fd_sc_hd__dlygate4sd3_1
X_19918_ _21099_/A vssd1 vssd1 vccd1 vccd1 _19918_/X sky130_fd_sc_hd__buf_8
XFILLER_0_43_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2727 _26254_/Q vssd1 vssd1 vccd1 vccd1 hold2727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2738 _26261_/Q vssd1 vssd1 vccd1 vccd1 hold2738/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2749 _25453_/Q vssd1 vssd1 vccd1 vccd1 _15416_/A sky130_fd_sc_hd__dlygate4sd3_1
X_19849_ _19849_/A _19849_/B vssd1 vssd1 vccd1 vccd1 _19849_/Y sky130_fd_sc_hd__nand2_1
X_22860_ _22860_/A _22860_/B vssd1 vssd1 vccd1 vccd1 _22861_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21811_ _18290_/A _25804_/Q _21809_/Y _21810_/Y vssd1 vssd1 vccd1 vccd1 _21812_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22791_ _23103_/B _22791_/B vssd1 vssd1 vccd1 vccd1 _22793_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24530_ _24530_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24531_/A sky130_fd_sc_hd__and2_1
XFILLER_0_176_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21742_ _22561_/B _21743_/A vssd1 vssd1 vccd1 vccd1 _21744_/A sky130_fd_sc_hd__or2_1
XFILLER_0_148_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24461_ hold2606/X _26218_/Q _24510_/S vssd1 vssd1 vccd1 vccd1 _24461_/X sky130_fd_sc_hd__mux2_1
X_21673_ _21676_/B _21677_/A vssd1 vssd1 vccd1 vccd1 _21675_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_148_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26200_ _26200_/CLK _26200_/D vssd1 vssd1 vccd1 vccd1 _26200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23412_ _23409_/Y _23411_/Y _24858_/S vssd1 vssd1 vccd1 vccd1 _23412_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_149_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20624_ _20624_/A _22248_/B vssd1 vssd1 vccd1 vccd1 _20625_/A sky130_fd_sc_hd__nand2_1
X_24392_ _24392_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24393_/A sky130_fd_sc_hd__and2_1
XFILLER_0_74_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26131_ _26135_/CLK _26131_/D vssd1 vssd1 vccd1 vccd1 _26131_/Q sky130_fd_sc_hd__dfxtp_1
X_23343_ _23343_/A _23377_/B _23347_/A vssd1 vssd1 vccd1 vccd1 _23344_/A sky130_fd_sc_hd__and3_1
XFILLER_0_62_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20555_ _20555_/A _20555_/B vssd1 vssd1 vccd1 vccd1 _21319_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_73_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26062_ _26065_/CLK _26062_/D vssd1 vssd1 vccd1 vccd1 _26062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23274_ _23272_/X hold830/X _12702_/A vssd1 vssd1 vccd1 vccd1 hold831/A sky130_fd_sc_hd__a21oi_1
X_20486_ _20486_/A _20486_/B vssd1 vssd1 vccd1 vccd1 _20488_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25013_ _25594_/CLK hold978/X vssd1 vssd1 vccd1 vccd1 hold977/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22225_ _22225_/A _22225_/B vssd1 vssd1 vccd1 vccd1 _23138_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_120_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22156_ _22823_/B vssd1 vssd1 vccd1 vccd1 _22824_/A sky130_fd_sc_hd__inv_2
XFILLER_0_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21107_ _21109_/C vssd1 vssd1 vccd1 vccd1 _21108_/B sky130_fd_sc_hd__inv_2
XFILLER_0_100_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22087_ _22586_/A vssd1 vssd1 vccd1 vccd1 _22561_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25915_ _26341_/CLK hold877/X vssd1 vssd1 vccd1 vccd1 hold875/A sky130_fd_sc_hd__dfxtp_1
X_21038_ _21038_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _21043_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25846_ _26336_/CLK _25846_/D vssd1 vssd1 vccd1 vccd1 _25846_/Q sky130_fd_sc_hd__dfxtp_4
X_13860_ _13941_/A _13860_/B vssd1 vssd1 vccd1 vccd1 _13860_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12811_ _17187_/B _14264_/A vssd1 vssd1 vccd1 vccd1 _12811_/X sky130_fd_sc_hd__or2_1
X_22989_ _22987_/X _22988_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _22989_/Y sky130_fd_sc_hd__a21oi_1
X_25777_ _26281_/CLK _25777_/D vssd1 vssd1 vccd1 vccd1 _25777_/Q sky130_fd_sc_hd__dfxtp_1
X_13791_ hold522/X _13790_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold523/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15530_ _15530_/A _16869_/A vssd1 vssd1 vccd1 vccd1 _15531_/B sky130_fd_sc_hd__nor2_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24728_ hold2610/X hold1959/X _24740_/S vssd1 vssd1 vccd1 vccd1 _24729_/A sky130_fd_sc_hd__mux2_1
X_12742_ _14125_/A vssd1 vssd1 vccd1 vccd1 _14260_/A sky130_fd_sc_hd__buf_12
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _12673_/A vssd1 vssd1 vccd1 vccd1 _24986_/D sky130_fd_sc_hd__clkbuf_1
X_15461_ _15447_/B _15466_/B _15442_/B vssd1 vssd1 vccd1 vccd1 _15461_/X sky130_fd_sc_hd__a21o_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_190_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _26284_/CLK sky130_fd_sc_hd__clkbuf_16
X_24659_ _24659_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24660_/A sky130_fd_sc_hd__and2_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17200_ _17393_/A _17200_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17200_/X sky130_fd_sc_hd__and3_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _14409_/Y hold408/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold409/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_182_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18180_ _18180_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _18180_/Y sky130_fd_sc_hd__nand2_1
X_15392_ _15392_/A _15405_/A vssd1 vssd1 vccd1 vccd1 _15392_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_64_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17131_ _20401_/B _25887_/Q _25823_/Q vssd1 vssd1 vccd1 vccd1 _17132_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_52_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26329_ _26330_/CLK _26329_/D vssd1 vssd1 vccd1 vccd1 _26329_/Q sky130_fd_sc_hd__dfxtp_2
X_14343_ _14343_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14343_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_64_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14274_ _23199_/C _14273_/X _12527_/A _14277_/A _14277_/B vssd1 vssd1 vccd1 vccd1
+ _14274_/X sky130_fd_sc_hd__o32a_1
X_17062_ _17060_/X _23187_/B _17061_/X vssd1 vssd1 vccd1 vccd1 _17063_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_162_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16013_ _16028_/B _16013_/B vssd1 vssd1 vccd1 vccd1 _16027_/B sky130_fd_sc_hd__nand2_1
X_13225_ _18515_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13225_/X sky130_fd_sc_hd__or2_1
XFILLER_0_100_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13156_ _18293_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13156_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17964_ _17962_/X _17528_/X _17963_/X vssd1 vssd1 vccd1 vccd1 _17965_/A sky130_fd_sc_hd__a21o_1
X_13087_ _13018_/X _13085_/X _13005_/X _13086_/X vssd1 vssd1 vccd1 vccd1 _13087_/X
+ sky130_fd_sc_hd__o211a_1
X_19703_ _20321_/A _19701_/Y _20326_/C vssd1 vssd1 vccd1 vccd1 _19793_/B sky130_fd_sc_hd__o21a_2
X_16915_ _16913_/Y _16914_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16915_/Y sky130_fd_sc_hd__a21oi_1
X_17895_ _18529_/A _17895_/B _18083_/C vssd1 vssd1 vccd1 vccd1 _17896_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19634_ _19635_/B _19635_/A vssd1 vssd1 vccd1 vccd1 _19634_/X sky130_fd_sc_hd__or2_1
X_16846_ _16935_/A _16851_/B vssd1 vssd1 vccd1 vccd1 _16848_/B sky130_fd_sc_hd__nand2_1
X_19565_ _19565_/A _19565_/B vssd1 vssd1 vccd1 vccd1 _19565_/Y sky130_fd_sc_hd__nand2_1
X_16777_ _15287_/A _16776_/Y _15621_/A vssd1 vssd1 vccd1 vccd1 _16777_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13989_ _25793_/Q vssd1 vssd1 vccd1 vccd1 _17909_/B sky130_fd_sc_hd__inv_2
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18516_ _18514_/X _18269_/X _18515_/X vssd1 vssd1 vccd1 vccd1 _18517_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_87_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15728_ hold883/X vssd1 vssd1 vccd1 vccd1 _15730_/A sky130_fd_sc_hd__inv_2
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19496_ _22902_/B vssd1 vssd1 vccd1 vccd1 _19496_/X sky130_fd_sc_hd__buf_8
XFILLER_0_87_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18447_ _18447_/A _25812_/Q _18447_/C vssd1 vssd1 vccd1 vccd1 _21296_/B sky130_fd_sc_hd__nand3_1
X_15659_ _15693_/C _15626_/B _15641_/A vssd1 vssd1 vccd1 vccd1 _15659_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_158_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_181_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _25796_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_185_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18378_ _19532_/A vssd1 vssd1 vccd1 vccd1 _21981_/B sky130_fd_sc_hd__inv_2
XFILLER_0_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17329_ _19458_/A _17329_/B vssd1 vssd1 vccd1 vccd1 _17578_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_172_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20340_ _20340_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20345_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_113_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20271_ _20269_/Y _20270_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _20271_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22010_ _22011_/B _22011_/A vssd1 vssd1 vccd1 vccd1 _22012_/A sky130_fd_sc_hd__or2_1
XFILLER_0_105_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2502 _25691_/Q vssd1 vssd1 vccd1 vccd1 _13353_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2513 _25698_/Q vssd1 vssd1 vccd1 vccd1 _13395_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2524 _24041_/X vssd1 vssd1 vccd1 vccd1 _24042_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2535 _24044_/X vssd1 vssd1 vccd1 vccd1 _24045_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2546 _25916_/Q vssd1 vssd1 vccd1 vccd1 _23269_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1801 _25626_/Q vssd1 vssd1 vccd1 vccd1 _17517_/B sky130_fd_sc_hd__dlygate4sd3_1
X_23961_ _23961_/A vssd1 vssd1 vccd1 vccd1 _26055_/D sky130_fd_sc_hd__clkbuf_1
Xhold1812 _21794_/Y vssd1 vssd1 vccd1 vccd1 _25839_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2557 _26239_/Q vssd1 vssd1 vccd1 vccd1 hold2557/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1823 _14905_/X vssd1 vssd1 vccd1 vccd1 _14906_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2568 _24559_/X vssd1 vssd1 vccd1 vccd1 _24561_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1834 _25623_/Q vssd1 vssd1 vccd1 vccd1 _17496_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2579 _24713_/X vssd1 vssd1 vccd1 vccd1 _24714_/A sky130_fd_sc_hd__dlygate4sd3_1
X_25700_ _26334_/CLK _25700_/D vssd1 vssd1 vccd1 vccd1 _25700_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1845 _25634_/Q vssd1 vssd1 vccd1 vccd1 _17575_/B sky130_fd_sc_hd__dlygate4sd3_1
X_22912_ _15509_/B _22680_/X _22829_/X vssd1 vssd1 vccd1 vccd1 _22912_/Y sky130_fd_sc_hd__a21oi_1
Xhold1856 _25853_/Q vssd1 vssd1 vccd1 vccd1 _22230_/B sky130_fd_sc_hd__dlygate4sd3_1
X_23892_ hold2080/X _26035_/Q _23907_/S vssd1 vssd1 vccd1 vccd1 _23892_/X sky130_fd_sc_hd__mux2_1
Xhold1867 _17554_/Y vssd1 vssd1 vccd1 vccd1 _25631_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1878 _25847_/Q vssd1 vssd1 vccd1 vccd1 _22058_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1889 _23785_/X vssd1 vssd1 vccd1 vccd1 _23786_/A sky130_fd_sc_hd__dlygate4sd3_1
X_22843_ _22994_/A _22843_/B vssd1 vssd1 vccd1 vccd1 _22844_/A sky130_fd_sc_hd__xor2_1
X_25631_ _25716_/CLK _25631_/D vssd1 vssd1 vccd1 vccd1 _25631_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_116_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25562_ _25878_/CLK _25562_/D vssd1 vssd1 vccd1 vccd1 _25562_/Q sky130_fd_sc_hd__dfxtp_1
X_22774_ _23087_/B _22774_/B vssd1 vssd1 vccd1 vccd1 _22776_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21725_ _21725_/A vssd1 vssd1 vccd1 vccd1 _21725_/X sky130_fd_sc_hd__buf_8
X_24513_ _24835_/S vssd1 vssd1 vccd1 vccd1 _24587_/S sky130_fd_sc_hd__buf_12
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25493_ _25495_/CLK hold550/X vssd1 vssd1 vccd1 vccd1 hold548/A sky130_fd_sc_hd__dfxtp_1
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_172_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _25727_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_176_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24444_ _24444_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24445_/A sky130_fd_sc_hd__and2_1
X_21656_ _21654_/Y _21655_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21656_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20607_ _21338_/B _21612_/A vssd1 vssd1 vccd1 vccd1 _20610_/A sky130_fd_sc_hd__nand2_1
X_24375_ hold2325/X hold2090/X _24433_/S vssd1 vssd1 vccd1 vccd1 _24377_/A sky130_fd_sc_hd__mux2_1
X_21587_ _21587_/A _21587_/B vssd1 vssd1 vccd1 vccd1 _21588_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_117_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23326_ _23326_/A vssd1 vssd1 vccd1 vccd1 _25927_/D sky130_fd_sc_hd__clkbuf_1
X_26114_ _26116_/CLK _26114_/D vssd1 vssd1 vccd1 vccd1 _26114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20538_ _26290_/Q hold728/X vssd1 vssd1 vccd1 vccd1 _20538_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_22_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23257_ _23275_/B vssd1 vssd1 vccd1 vccd1 _23258_/A sky130_fd_sc_hd__inv_2
X_26045_ _26046_/CLK _26045_/D vssd1 vssd1 vccd1 vccd1 _26045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20469_ _20472_/A _20472_/C vssd1 vssd1 vccd1 vccd1 _20470_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ _26135_/Q _12907_/X _13009_/X vssd1 vssd1 vccd1 vccd1 _13010_/X sky130_fd_sc_hd__a21o_1
X_22208_ _25817_/Q _22208_/B vssd1 vssd1 vccd1 vccd1 _22208_/Y sky130_fd_sc_hd__nor2_1
X_23188_ _23188_/A _23188_/B vssd1 vssd1 vccd1 vccd1 _23188_/X sky130_fd_sc_hd__or2_1
X_22139_ _22139_/A _23090_/A _22139_/C vssd1 vssd1 vccd1 vccd1 _22139_/Y sky130_fd_sc_hd__nand3_1
X_14961_ _14962_/B _14962_/A vssd1 vssd1 vccd1 vccd1 _14963_/A sky130_fd_sc_hd__or2_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
X_16700_ _16773_/A vssd1 vssd1 vccd1 vccd1 _16858_/A sky130_fd_sc_hd__clkbuf_8
X_13912_ _14000_/A hold736/X vssd1 vssd1 vccd1 vccd1 hold737/A sky130_fd_sc_hd__nand2_1
X_17680_ _17688_/A _25905_/Q _17707_/B vssd1 vssd1 vccd1 vccd1 _17692_/B sky130_fd_sc_hd__nand3_1
X_14892_ _14890_/Y _14891_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14892_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16631_ _16629_/A _16607_/A _16618_/B vssd1 vssd1 vccd1 vccd1 _16631_/Y sky130_fd_sc_hd__a21oi_1
X_25829_ _25864_/CLK _25829_/D vssd1 vssd1 vccd1 vccd1 _25829_/Q sky130_fd_sc_hd__dfxtp_4
X_13843_ hold813/X _13842_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold814/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19350_ _19350_/A _19350_/B vssd1 vssd1 vccd1 vccd1 _19350_/Y sky130_fd_sc_hd__nand2_1
X_16562_ _16562_/A _16562_/B vssd1 vssd1 vccd1 vccd1 _16563_/A sky130_fd_sc_hd__nor2_1
X_13774_ _13880_/A hold713/X vssd1 vssd1 vccd1 vccd1 _13774_/Y sky130_fd_sc_hd__nand2_1
X_18301_ _18301_/A _18301_/B vssd1 vssd1 vccd1 vccd1 _21843_/A sky130_fd_sc_hd__nand2_1
X_15513_ hold878/X vssd1 vssd1 vccd1 vccd1 _15515_/A sky130_fd_sc_hd__inv_2
XFILLER_0_57_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19281_ _19279_/X _19280_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19281_/Y sky130_fd_sc_hd__a21oi_1
X_12725_ _26213_/Q _25582_/Q vssd1 vssd1 vccd1 vccd1 _14287_/A sky130_fd_sc_hd__xor2_1
X_16493_ _16486_/B _16479_/A _16468_/B _16478_/A _16492_/X vssd1 vssd1 vccd1 vccd1
+ _16493_/X sky130_fd_sc_hd__o311a_1
Xclkbuf_leaf_163_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _26298_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18232_ _18252_/A _18232_/B vssd1 vssd1 vccd1 vccd1 _18232_/Y sky130_fd_sc_hd__nand2_1
X_15444_ _15467_/B _15414_/A vssd1 vssd1 vccd1 vccd1 _15446_/A sky130_fd_sc_hd__or2b_1
X_12656_ _12656_/A _12656_/B vssd1 vssd1 vccd1 vccd1 _12664_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18163_ _21938_/B _25607_/Q vssd1 vssd1 vccd1 vccd1 _18165_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15375_ _15406_/C _15342_/B _15357_/A vssd1 vssd1 vccd1 vccd1 _15375_/X sky130_fd_sc_hd__a21o_1
X_12587_ _12587_/A _23923_/B vssd1 vssd1 vccd1 vccd1 _12588_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17114_ _25596_/Q vssd1 vssd1 vccd1 vccd1 _20547_/B sky130_fd_sc_hd__inv_2
XFILLER_0_80_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14326_ _14344_/A hold332/X vssd1 vssd1 vccd1 vccd1 hold333/A sky130_fd_sc_hd__nand2_1
XFILLER_0_123_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18094_ _25861_/Q _21868_/A vssd1 vssd1 vccd1 vccd1 _18104_/A sky130_fd_sc_hd__or2_2
XFILLER_0_64_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold408 hold408/A vssd1 vssd1 vccd1 vccd1 hold408/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17045_ _17393_/A _17045_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17045_/X sky130_fd_sc_hd__and3_1
Xhold419 hold419/A vssd1 vssd1 vccd1 vccd1 hold419/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_14257_ _26339_/Q _13518_/B _14170_/X _14256_/Y vssd1 vssd1 vccd1 vccd1 _14258_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13208_ _13208_/A vssd1 vssd1 vccd1 vccd1 _19345_/A sky130_fd_sc_hd__buf_4
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14188_ _14236_/A hold422/X vssd1 vssd1 vccd1 vccd1 hold423/A sky130_fd_sc_hd__nand2_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13139_ _18229_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13139_/X sky130_fd_sc_hd__or2_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ _18996_/A _19066_/B vssd1 vssd1 vccd1 vccd1 _18997_/B sky130_fd_sc_hd__xnor2_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ _17947_/A _20506_/A vssd1 vssd1 vccd1 vccd1 _19059_/A sky130_fd_sc_hd__xor2_4
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1108 _12955_/X vssd1 vssd1 vccd1 vccd1 _25041_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1119 _25734_/Q vssd1 vssd1 vccd1 vccd1 _19467_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17878_ _17878_/A _17878_/B vssd1 vssd1 vccd1 vccd1 _17881_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_136_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16829_ _16935_/A _16834_/B vssd1 vssd1 vccd1 vccd1 _16831_/B sky130_fd_sc_hd__nand2_1
X_19617_ _20098_/A _22149_/B _25623_/Q vssd1 vssd1 vccd1 vccd1 _20102_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_177_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19548_ _21237_/A _19546_/Y _21241_/C vssd1 vssd1 vccd1 vccd1 _19635_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_48_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19479_ _19477_/X _19478_/Y _19146_/X vssd1 vssd1 vccd1 vccd1 _19479_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_154_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _26305_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_146_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21510_ _21508_/Y _21509_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21510_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22490_ _22490_/A _22490_/B vssd1 vssd1 vccd1 vccd1 _22490_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_118_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21441_ _21636_/A _21441_/B _21440_/X vssd1 vssd1 vccd1 vccd1 _21442_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24160_ hold2324/X hold2233/X _24203_/S vssd1 vssd1 vccd1 vccd1 _24161_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_71_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21372_ _21372_/A _21372_/B vssd1 vssd1 vccd1 vccd1 _21373_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23111_ _23111_/A _23111_/B _23191_/C vssd1 vssd1 vccd1 vccd1 _23113_/A sky130_fd_sc_hd__or3_1
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20323_ _20326_/A _20326_/C vssd1 vssd1 vccd1 vccd1 _20324_/A sky130_fd_sc_hd__nand2_1
X_24091_ _24091_/A vssd1 vssd1 vccd1 vccd1 _26097_/D sky130_fd_sc_hd__clkbuf_1
Xhold920 hold920/A vssd1 vssd1 vccd1 vccd1 hold920/X sky130_fd_sc_hd__buf_1
XFILLER_0_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold931 hold931/A vssd1 vssd1 vccd1 vccd1 hold931/X sky130_fd_sc_hd__buf_1
XFILLER_0_101_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold942 hold942/A vssd1 vssd1 vccd1 vccd1 hold942/X sky130_fd_sc_hd__buf_1
X_23042_ _23042_/A _23042_/B vssd1 vssd1 vccd1 vccd1 _23043_/A sky130_fd_sc_hd__xor2_2
Xhold953 hold953/A vssd1 vssd1 vccd1 vccd1 hold953/X sky130_fd_sc_hd__dlygate4sd3_1
X_20254_ _20254_/A _20254_/B _20254_/C vssd1 vssd1 vccd1 vccd1 _20255_/B sky130_fd_sc_hd__nand3_1
Xhold964 hold964/A vssd1 vssd1 vccd1 vccd1 hold964/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 hold975/A vssd1 vssd1 vccd1 vccd1 hold975/X sky130_fd_sc_hd__buf_1
XFILLER_0_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold986 hold986/A vssd1 vssd1 vccd1 vccd1 hold986/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 hold997/A vssd1 vssd1 vccd1 vccd1 hold997/X sky130_fd_sc_hd__buf_1
X_20185_ _20187_/A _20187_/B vssd1 vssd1 vccd1 vccd1 _20186_/A sky130_fd_sc_hd__nand2_1
Xhold2310 _26198_/Q vssd1 vssd1 vccd1 vccd1 hold2310/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2321 _26200_/Q vssd1 vssd1 vccd1 vccd1 hold2321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2332 _26179_/Q vssd1 vssd1 vccd1 vccd1 hold2332/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2343 _26024_/Q vssd1 vssd1 vccd1 vccd1 hold2343/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24993_ _25491_/CLK hold838/X vssd1 vssd1 vccd1 vccd1 hold837/A sky130_fd_sc_hd__dfxtp_1
Xhold2354 _26127_/Q vssd1 vssd1 vccd1 vccd1 hold2354/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1620 _25618_/Q vssd1 vssd1 vccd1 vccd1 _17460_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2365 _25678_/Q vssd1 vssd1 vccd1 vccd1 _13271_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2376 _15040_/Y vssd1 vssd1 vccd1 vccd1 _25428_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1631 _17113_/Y vssd1 vssd1 vccd1 vccd1 _25588_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23944_ hold2469/X hold2401/X _24001_/S vssd1 vssd1 vccd1 vccd1 _23945_/A sky130_fd_sc_hd__mux2_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1642 _21263_/Y vssd1 vssd1 vccd1 vccd1 _25810_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2387 _25686_/Q vssd1 vssd1 vccd1 vccd1 _13322_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2398 _25450_/Q vssd1 vssd1 vccd1 vccd1 _15363_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1653 _25782_/Q vssd1 vssd1 vccd1 vccd1 _20347_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1664 _22790_/Y vssd1 vssd1 vccd1 vccd1 _25876_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1675 _17081_/Y vssd1 vssd1 vccd1 vccd1 _25586_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1686 _20934_/Y vssd1 vssd1 vccd1 vccd1 _25798_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23875_ _23875_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23876_/A sky130_fd_sc_hd__and2_1
Xhold1697 _22955_/Y vssd1 vssd1 vccd1 vccd1 _25886_/D sky130_fd_sc_hd__dlygate4sd3_1
X_25614_ _26117_/CLK _25614_/D vssd1 vssd1 vccd1 vccd1 _25614_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_67_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22826_ _22977_/A _22826_/B vssd1 vssd1 vccd1 vccd1 _22827_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25545_ _26053_/CLK _25545_/D vssd1 vssd1 vccd1 vccd1 _25545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22757_ _22755_/X _22756_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22757_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_145_clk clkbuf_4_11__f_clk/X vssd1 vssd1 vccd1 vccd1 _26313_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_149_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12510_ _24991_/Q _24990_/Q _24989_/Q _24988_/Q vssd1 vssd1 vccd1 vccd1 _12514_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_0_94_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13490_ _13583_/A _13490_/B vssd1 vssd1 vccd1 vccd1 _13490_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21708_ _21708_/A _21708_/B vssd1 vssd1 vccd1 vccd1 _21710_/A sky130_fd_sc_hd__nand2_1
X_25476_ _25913_/CLK hold508/X vssd1 vssd1 vccd1 vccd1 hold506/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22688_ _22677_/Y _22687_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22688_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24427_ hold2344/X hold2089/X _24433_/S vssd1 vssd1 vccd1 vccd1 _24428_/A sky130_fd_sc_hd__mux2_1
X_21639_ _22058_/A _21639_/B vssd1 vssd1 vccd1 vccd1 _21639_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15160_ _15160_/A _16726_/A vssd1 vssd1 vccd1 vccd1 _15161_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24358_ _24358_/A vssd1 vssd1 vccd1 vccd1 _26184_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14111_ hold528/X _14110_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold529/A sky130_fd_sc_hd__a21oi_1
X_23309_ _23317_/A vssd1 vssd1 vccd1 vccd1 _23314_/A sky130_fd_sc_hd__inv_2
X_15091_ _15088_/X hold2148/X _15090_/X vssd1 vssd1 vccd1 vccd1 _15091_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24289_ _24289_/A vssd1 vssd1 vccd1 vccd1 _26161_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26028_ _26032_/CLK _26028_/D vssd1 vssd1 vccd1 vccd1 _26028_/Q sky130_fd_sc_hd__dfxtp_1
X_14042_ _26304_/Q _13988_/X _13981_/X _14041_/Y vssd1 vssd1 vccd1 vccd1 _14043_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18850_ _18952_/A _25768_/Q _18952_/C vssd1 vssd1 vccd1 vccd1 _18851_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17801_ _17801_/A _17801_/B _17801_/C vssd1 vssd1 vccd1 vccd1 _22078_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_98_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18781_ _18781_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18781_/Y sky130_fd_sc_hd__nand2_1
X_15993_ hold798/X vssd1 vssd1 vccd1 vccd1 _15996_/B sky130_fd_sc_hd__inv_2
XFILLER_0_101_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17732_ _17734_/B vssd1 vssd1 vccd1 vccd1 _17733_/B sky130_fd_sc_hd__inv_2
X_14944_ _14945_/B _14945_/A vssd1 vssd1 vccd1 vccd1 _14946_/A sky130_fd_sc_hd__or2_1
X_17663_ _25902_/Q _25710_/Q vssd1 vssd1 vccd1 vccd1 _17665_/A sky130_fd_sc_hd__xor2_1
X_14875_ _15839_/A _14875_/B vssd1 vssd1 vccd1 vccd1 _22344_/A sky130_fd_sc_hd__nand2_1
X_19402_ _19402_/A _20965_/B vssd1 vssd1 vccd1 vccd1 _19402_/Y sky130_fd_sc_hd__nor2_1
X_16614_ _16612_/X _16613_/Y _16594_/X vssd1 vssd1 vccd1 vccd1 hold872/A sky130_fd_sc_hd__a21oi_1
X_13826_ _13944_/A vssd1 vssd1 vccd1 vccd1 _13941_/A sky130_fd_sc_hd__buf_8
X_17594_ _17594_/A _17594_/B vssd1 vssd1 vccd1 vccd1 _17594_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19333_ _20817_/A _19331_/Y _20822_/C vssd1 vssd1 vccd1 vccd1 _19421_/B sky130_fd_sc_hd__o21a_2
X_16545_ _16599_/A _16545_/B vssd1 vssd1 vccd1 vccd1 _16554_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_175_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_136_clk clkbuf_leaf_82_clk/A vssd1 vssd1 vccd1 vccd1 _25827_/CLK sky130_fd_sc_hd__clkbuf_16
X_13757_ _26259_/Q _13612_/X _13605_/X _13756_/Y vssd1 vssd1 vccd1 vccd1 _13758_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12708_ hold997/X hold837/X vssd1 vssd1 vccd1 vccd1 _12714_/A sky130_fd_sc_hd__nand2_1
X_19264_ _26223_/Q _19483_/A hold509/X vssd1 vssd1 vccd1 vccd1 _19265_/C sky130_fd_sc_hd__a21o_1
X_16476_ _16483_/B _16477_/A vssd1 vssd1 vccd1 vccd1 _16479_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_155_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13688_ _25745_/Q vssd1 vssd1 vccd1 vccd1 _18387_/B sky130_fd_sc_hd__inv_2
XFILLER_0_85_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18215_ _22006_/B _25609_/Q vssd1 vssd1 vccd1 vccd1 _18217_/A sky130_fd_sc_hd__nand2_1
X_15427_ _15427_/A vssd1 vssd1 vccd1 vccd1 _15443_/B sky130_fd_sc_hd__inv_2
X_12639_ _12654_/A _12654_/C vssd1 vssd1 vccd1 vccd1 _12639_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_115_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19195_ _19195_/A _19994_/B _19195_/C vssd1 vssd1 vccd1 vccd1 _19195_/X sky130_fd_sc_hd__and3_1
XFILLER_0_155_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18146_ _18146_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _18146_/Y sky130_fd_sc_hd__nand2_1
X_15358_ _15406_/C vssd1 vssd1 vccd1 vccd1 _15361_/B sky130_fd_sc_hd__inv_2
XFILLER_0_171_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14309_ _14307_/Y hold279/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold280/A sky130_fd_sc_hd__a21oi_1
Xhold205 hold205/A vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
X_18077_ _19257_/A vssd1 vssd1 vccd1 vccd1 _22248_/B sky130_fd_sc_hd__inv_2
X_15289_ _15290_/B _15290_/A vssd1 vssd1 vccd1 vccd1 _15291_/A sky130_fd_sc_hd__nor2_1
Xhold216 hold216/A vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 hold227/A vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 hold238/A vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17028_ _17616_/A _17028_/B vssd1 vssd1 vccd1 vccd1 _17028_/X sky130_fd_sc_hd__xor2_1
Xhold249 hold249/A vssd1 vssd1 vccd1 vccd1 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ _18986_/A _19715_/A vssd1 vssd1 vccd1 vccd1 _18979_/Y sky130_fd_sc_hd__nand2_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21990_ _22245_/A _23168_/A vssd1 vssd1 vccd1 vccd1 _21996_/B sky130_fd_sc_hd__nand2_1
X_20941_ _20944_/A _20944_/C vssd1 vssd1 vccd1 vccd1 _20943_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23660_ _23660_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23661_/A sky130_fd_sc_hd__and2_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20872_ _20872_/A _20872_/B vssd1 vssd1 vccd1 vccd1 _20873_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_138_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22611_ _22602_/Y _22610_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22611_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23591_ hold875/X _24871_/B vssd1 vssd1 vccd1 vccd1 _23592_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_159_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_127_clk clkbuf_4_14__f_clk/X vssd1 vssd1 vccd1 vccd1 _25708_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22542_ _19830_/A _22541_/A _22541_/Y vssd1 vssd1 vccd1 vccd1 _22544_/A sky130_fd_sc_hd__o21ai_1
X_25330_ _25650_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22473_ _22473_/A _22473_/B vssd1 vssd1 vccd1 vccd1 _22474_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_17_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25261_ _26122_/CLK hold265/X vssd1 vssd1 vccd1 vccd1 hold263/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24212_ _24212_/A vssd1 vssd1 vccd1 vccd1 _26136_/D sky130_fd_sc_hd__clkbuf_1
X_21424_ _21423_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21424_/X
+ sky130_fd_sc_hd__a211o_1
X_25192_ _26275_/CLK hold808/X vssd1 vssd1 vccd1 vccd1 hold806/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24143_ _24143_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24144_/A sky130_fd_sc_hd__and2_1
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21355_ _21355_/A _21355_/B vssd1 vssd1 vccd1 vccd1 _21356_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_170_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20306_ _20306_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _20306_/Y sky130_fd_sc_hd__nand2_1
X_24074_ hold2164/X hold2255/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24075_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_102_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21286_ _21286_/A _21286_/B vssd1 vssd1 vccd1 vccd1 _21287_/A sky130_fd_sc_hd__nand2_1
Xhold750 hold750/A vssd1 vssd1 vccd1 vccd1 hold750/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 hold761/A vssd1 vssd1 vccd1 vccd1 hold761/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 hold772/A vssd1 vssd1 vccd1 vccd1 hold772/X sky130_fd_sc_hd__dlygate4sd3_1
X_23025_ _23025_/A _23025_/B vssd1 vssd1 vccd1 vccd1 _23026_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold783 hold783/A vssd1 vssd1 vccd1 vccd1 hold783/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20237_ _20240_/A _20240_/C vssd1 vssd1 vccd1 vccd1 _20238_/A sky130_fd_sc_hd__nand2_1
Xhold794 hold794/A vssd1 vssd1 vccd1 vccd1 hold794/X sky130_fd_sc_hd__dlygate4sd3_1
X_20168_ _20171_/A _20171_/C vssd1 vssd1 vccd1 vccd1 _20170_/A sky130_fd_sc_hd__nand2_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2140 _25944_/Q vssd1 vssd1 vccd1 vccd1 hold2140/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2151 _23372_/Y vssd1 vssd1 vccd1 vccd1 _23373_/C sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2162 _23727_/X vssd1 vssd1 vccd1 vccd1 _23728_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2173 _23320_/Y vssd1 vssd1 vccd1 vccd1 _23321_/C sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24976_ _25420_/CLK _24976_/D vssd1 vssd1 vccd1 vccd1 _24976_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _17529_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _12990_/X sky130_fd_sc_hd__or2_1
X_20099_ _20099_/A _20099_/B vssd1 vssd1 vccd1 vccd1 _20102_/B sky130_fd_sc_hd__nand2_1
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2184 _23962_/X vssd1 vssd1 vccd1 vccd1 _23963_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2195 _15005_/X vssd1 vssd1 vccd1 vccd1 _15007_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1450 _14823_/Y vssd1 vssd1 vccd1 vccd1 _25402_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1461 _25737_/Q vssd1 vssd1 vccd1 vccd1 _19512_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1472 _14787_/Y vssd1 vssd1 vccd1 vccd1 _25398_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23927_ _23927_/A vssd1 vssd1 vccd1 vccd1 _24047_/S sky130_fd_sc_hd__buf_8
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1483 _25771_/Q vssd1 vssd1 vccd1 vccd1 _19975_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1494 _13294_/X vssd1 vssd1 vccd1 vccd1 _25101_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _14660_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _14660_/Y sky130_fd_sc_hd__nand2_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23858_ _23858_/A vssd1 vssd1 vccd1 vccd1 _26023_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _13642_/A hold599/X vssd1 vssd1 vccd1 vccd1 hold600/A sky130_fd_sc_hd__nand2_1
XFILLER_0_95_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22809_ _22809_/A _22809_/B vssd1 vssd1 vccd1 vccd1 _22810_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_184_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_118_clk clkbuf_4_14__f_clk/X vssd1 vssd1 vccd1 vccd1 _26202_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14591_ _14645_/A hold185/X vssd1 vssd1 vccd1 vccd1 hold186/A sky130_fd_sc_hd__nand2_1
X_23789_ _23789_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23790_/A sky130_fd_sc_hd__and2_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16330_ _16331_/B _16331_/A vssd1 vssd1 vccd1 vccd1 _16332_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25528_ _25533_/CLK hold905/X vssd1 vssd1 vccd1 vccd1 hold904/A sky130_fd_sc_hd__dfxtp_1
X_13542_ _13642_/A hold419/X vssd1 vssd1 vccd1 vccd1 hold420/A sky130_fd_sc_hd__nand2_1
XFILLER_0_137_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16261_ _16262_/B _16262_/A vssd1 vssd1 vccd1 vccd1 _16263_/A sky130_fd_sc_hd__or2_1
XFILLER_0_153_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25459_ _26064_/CLK _25459_/D vssd1 vssd1 vccd1 vccd1 _25459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13473_ hold453/X _13472_/Y _12558_/B vssd1 vssd1 vccd1 vccd1 hold454/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18000_ _18000_/A _25795_/Q _18000_/C vssd1 vssd1 vccd1 vccd1 _20824_/B sky130_fd_sc_hd__nand3_1
X_15212_ _15213_/B _16747_/A vssd1 vssd1 vccd1 vccd1 _15214_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_106_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16192_ _22501_/B _16369_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _16195_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_164_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15143_ _15144_/B _16719_/A vssd1 vssd1 vccd1 vccd1 _15145_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_152_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15074_ _15072_/X hold2305/X _14928_/X vssd1 vssd1 vccd1 vccd1 _15074_/Y sky130_fd_sc_hd__a21oi_1
X_19951_ _19949_/X _19950_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19951_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14025_ hold636/X _14024_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold637/A sky130_fd_sc_hd__a21oi_1
X_18902_ _18902_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18902_/Y sky130_fd_sc_hd__nand2_1
X_19882_ _26267_/Q _19134_/X hold944/X vssd1 vssd1 vccd1 vccd1 _19883_/C sky130_fd_sc_hd__a21o_1
X_18833_ _18955_/A _18833_/B _18894_/C vssd1 vssd1 vccd1 vccd1 _18834_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_184_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18764_ _19802_/A vssd1 vssd1 vccd1 vccd1 _22488_/B sky130_fd_sc_hd__inv_2
X_15976_ _16000_/B _16000_/A _15953_/B _15975_/Y vssd1 vssd1 vccd1 vccd1 _15978_/A
+ sky130_fd_sc_hd__o31ai_1
XFILLER_0_175_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17715_ _17719_/A _17719_/B _25905_/Q vssd1 vssd1 vccd1 vccd1 _17726_/C sky130_fd_sc_hd__nand3_1
X_14927_ _14927_/A _14927_/B vssd1 vssd1 vccd1 vccd1 _14927_/Y sky130_fd_sc_hd__nand2_1
X_18695_ _20447_/B _22393_/A vssd1 vssd1 vccd1 vccd1 _20438_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17646_ _18535_/A _17646_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _17646_/X sky130_fd_sc_hd__and3_1
X_14858_ _14900_/A _14860_/A vssd1 vssd1 vccd1 vccd1 _14858_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13809_ _18773_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13809_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_109_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _25425_/CLK sky130_fd_sc_hd__clkbuf_16
X_17577_ _17577_/A _17629_/A vssd1 vssd1 vccd1 vccd1 _17578_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14789_ _14795_/B _22061_/A vssd1 vssd1 vccd1 vccd1 _22060_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19316_ _19313_/Y _19316_/B _19980_/B vssd1 vssd1 vccd1 vccd1 _19316_/X sky130_fd_sc_hd__and3b_1
X_16528_ _16528_/A _16541_/A vssd1 vssd1 vccd1 vccd1 _16537_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19247_ _19261_/A _19336_/B vssd1 vssd1 vccd1 vccd1 _19248_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16459_ _16457_/X _16458_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 hold936/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19178_ _19177_/A _19176_/Y _20214_/C vssd1 vssd1 vccd1 vccd1 _19989_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_182_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18129_ _19373_/A vssd1 vssd1 vccd1 vccd1 _21904_/B sky130_fd_sc_hd__inv_2
XFILLER_0_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21140_ _21613_/B _21564_/B vssd1 vssd1 vccd1 vccd1 _21141_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_44_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21071_ _21071_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _21071_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_158_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20022_ _21369_/A _21677_/A vssd1 vssd1 vccd1 vccd1 _20028_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24830_ _24830_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24831_/A sky130_fd_sc_hd__and2_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24761_ _24761_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24762_/A sky130_fd_sc_hd__and2_1
XFILLER_0_179_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21973_ _18205_/A _25800_/Q _21971_/Y _21972_/Y vssd1 vssd1 vccd1 vccd1 _21974_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23712_ _23712_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23713_/A sky130_fd_sc_hd__and2_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20924_ _20924_/A _21432_/C _20924_/C vssd1 vssd1 vccd1 vccd1 _20925_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_179_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24692_ hold2744/X hold2638/X _24740_/S vssd1 vssd1 vccd1 vccd1 _24693_/A sky130_fd_sc_hd__mux2_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23643_ _23643_/A vssd1 vssd1 vccd1 vccd1 _25953_/D sky130_fd_sc_hd__clkbuf_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20855_ _20855_/A _21835_/B vssd1 vssd1 vccd1 vccd1 _20856_/A sky130_fd_sc_hd__nand2_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23574_ hold146/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23574_/X sky130_fd_sc_hd__or2b_1
X_20786_ _20786_/A _20786_/B vssd1 vssd1 vccd1 vccd1 _20788_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25313_ _26142_/CLK hold343/X vssd1 vssd1 vccd1 vccd1 hold341/A sky130_fd_sc_hd__dfxtp_1
X_22525_ _22525_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _22525_/Y sky130_fd_sc_hd__nand2_1
X_26293_ _26296_/CLK _26293_/D vssd1 vssd1 vccd1 vccd1 _26293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25244_ _25709_/CLK hold824/X vssd1 vssd1 vccd1 vccd1 hold823/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22456_ _22456_/A _23001_/B _22456_/C vssd1 vssd1 vccd1 vccd1 _22456_/X sky130_fd_sc_hd__and3_1
XFILLER_0_162_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21407_ _26321_/Q hold434/X vssd1 vssd1 vccd1 vccd1 _21407_/Y sky130_fd_sc_hd__nand2_1
X_22387_ _22387_/A _22387_/B vssd1 vssd1 vccd1 vccd1 _22387_/Y sky130_fd_sc_hd__nand2_1
X_25175_ _25756_/CLK hold526/X vssd1 vssd1 vccd1 vccd1 hold524/A sky130_fd_sc_hd__dfxtp_1
X_24126_ hold2279/X hold2257/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24127_/A sky130_fd_sc_hd__mux2_1
X_21338_ _21338_/A _21338_/B _21338_/C vssd1 vssd1 vccd1 vccd1 _21339_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_102_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24057_ _24057_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24058_/A sky130_fd_sc_hd__and2_1
X_21269_ _21271_/B _21271_/C vssd1 vssd1 vccd1 vccd1 _21270_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold580 hold580/A vssd1 vssd1 vccd1 vccd1 hold580/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 hold591/A vssd1 vssd1 vccd1 vccd1 hold591/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23008_ _23154_/A _23008_/B vssd1 vssd1 vccd1 vccd1 _23009_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15830_ _15830_/A _15830_/B vssd1 vssd1 vccd1 vccd1 _15830_/Y sky130_fd_sc_hd__nand2_1
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _16960_/A _15761_/B vssd1 vssd1 vccd1 vccd1 _15762_/B sky130_fd_sc_hd__nand2_1
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24959_ _24959_/A _24959_/B _24959_/C vssd1 vssd1 vccd1 vccd1 _24959_/X sky130_fd_sc_hd__and3_1
X_12973_ _26128_/Q _12907_/X _12972_/X vssd1 vssd1 vccd1 vccd1 _12973_/X sky130_fd_sc_hd__a21o_1
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1280 _25084_/Q vssd1 vssd1 vccd1 vccd1 _18393_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17500_ _17624_/A _17500_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17500_/X sky130_fd_sc_hd__and3_1
XFILLER_0_87_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _14900_/A _14712_/B vssd1 vssd1 vccd1 vccd1 _14712_/Y sky130_fd_sc_hd__nand2_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1291 _20739_/Y vssd1 vssd1 vccd1 vccd1 _25792_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18480_ _19602_/A vssd1 vssd1 vccd1 vccd1 _22120_/B sky130_fd_sc_hd__inv_2
X_15692_ _15692_/A _15692_/B vssd1 vssd1 vccd1 vccd1 _15693_/A sky130_fd_sc_hd__nor2_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _20055_/B _25878_/Q _25814_/Q vssd1 vssd1 vccd1 vccd1 _17432_/B sky130_fd_sc_hd__mux2_2
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14643_ _14641_/Y hold468/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold469/A sky130_fd_sc_hd__a21oi_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17362_ _17630_/A _17362_/B vssd1 vssd1 vccd1 vccd1 _17362_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_184_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14574_ _14572_/Y hold177/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold178/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19101_ _19990_/A _19101_/B vssd1 vssd1 vccd1 vccd1 _19101_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_94_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16313_ _16313_/A _16313_/B vssd1 vssd1 vccd1 vccd1 _16322_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_126_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13525_ _18186_/B _13638_/B vssd1 vssd1 vccd1 vccd1 _13525_/Y sky130_fd_sc_hd__nor2_1
X_17293_ _25707_/Q _17293_/B vssd1 vssd1 vccd1 vccd1 _17637_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_165_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19032_ _19032_/A _19032_/B vssd1 vssd1 vccd1 vccd1 _19032_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_42_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16244_ _16237_/A _16223_/A _16236_/B vssd1 vssd1 vccd1 vccd1 _16252_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13456_ _19075_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13456_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16175_ _16212_/A hold754/X vssd1 vssd1 vccd1 vccd1 hold755/A sky130_fd_sc_hd__nand2_1
X_13387_ _18990_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13387_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15126_ _16660_/B vssd1 vssd1 vccd1 vccd1 _16231_/A sky130_fd_sc_hd__inv_6
XFILLER_0_142_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15057_ _15058_/B _15058_/A vssd1 vssd1 vccd1 vccd1 _15059_/A sky130_fd_sc_hd__or2_1
X_19934_ _19933_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19936_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_120_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14008_ _14118_/A hold578/X vssd1 vssd1 vccd1 vccd1 hold579/A sky130_fd_sc_hd__nand2_1
X_19865_ _19975_/A _19865_/B vssd1 vssd1 vccd1 vccd1 _19865_/Y sky130_fd_sc_hd__nand2_1
X_18816_ _18816_/A _20672_/A vssd1 vssd1 vccd1 vccd1 _19031_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19796_ _19975_/A _19796_/B vssd1 vssd1 vccd1 vccd1 _19796_/Y sky130_fd_sc_hd__nand2_1
X_15959_ _22035_/B hold929/X _16691_/B vssd1 vssd1 vccd1 vccd1 _15960_/B sky130_fd_sc_hd__nand3_1
X_18747_ _18747_/A _18747_/B vssd1 vssd1 vccd1 vccd1 _22462_/A sky130_fd_sc_hd__nand2_1
X_18678_ _18678_/A _18678_/B vssd1 vssd1 vccd1 vccd1 _18678_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_77_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17629_ _17629_/A _17629_/B vssd1 vssd1 vccd1 vccd1 _17630_/B sky130_fd_sc_hd__xnor2_1
X_20640_ _20643_/A _20643_/C vssd1 vssd1 vccd1 vccd1 _20642_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_86_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20571_ _20571_/A _20571_/B _21249_/C vssd1 vssd1 vccd1 vccd1 _20575_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_160_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22310_ _22310_/A _22310_/B vssd1 vssd1 vccd1 vccd1 _22310_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23290_ _23290_/A hold855/X vssd1 vssd1 vccd1 vccd1 hold856/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22241_ _25882_/Q _22242_/A vssd1 vssd1 vccd1 vccd1 _22243_/A sky130_fd_sc_hd__or2_1
XFILLER_0_6_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22172_ _22170_/Y _22171_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _22172_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21123_ _21636_/A _21123_/B _21122_/X vssd1 vssd1 vccd1 vccd1 _21124_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_2_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25931_ _25939_/CLK _25931_/D vssd1 vssd1 vccd1 vccd1 _25931_/Q sky130_fd_sc_hd__dfxtp_1
X_21054_ _21053_/B _21054_/B _21054_/C vssd1 vssd1 vccd1 vccd1 _21055_/B sky130_fd_sc_hd__nand3b_1
X_20005_ _20007_/B _20007_/C vssd1 vssd1 vccd1 vccd1 _20006_/A sky130_fd_sc_hd__nand2_1
X_25862_ _25864_/CLK _25862_/D vssd1 vssd1 vccd1 vccd1 _25862_/Q sky130_fd_sc_hd__dfxtp_4
X_24813_ _24813_/A vssd1 vssd1 vccd1 vccd1 _26332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25793_ _25793_/CLK _25793_/D vssd1 vssd1 vccd1 vccd1 _25793_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24744_ hold2625/X hold2604/X _24817_/S vssd1 vssd1 vccd1 vccd1 _24746_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21956_ _22216_/A _23152_/A vssd1 vssd1 vccd1 vccd1 _21962_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _20905_/Y _20906_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _20907_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_179_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24675_ _24675_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24676_/A sky130_fd_sc_hd__and2_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21887_ _22157_/A _23120_/A vssd1 vssd1 vccd1 vccd1 _21893_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23626_ _23626_/A _23629_/B vssd1 vssd1 vccd1 vccd1 _23627_/A sky130_fd_sc_hd__and2_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20838_ _21432_/C _21709_/B vssd1 vssd1 vccd1 vccd1 _20841_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_154_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23557_ _24922_/S hold467/A _23556_/X vssd1 vssd1 vccd1 vccd1 _23557_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_181_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20769_ _22704_/A vssd1 vssd1 vccd1 vccd1 _21281_/B sky130_fd_sc_hd__buf_6
XFILLER_0_181_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13310_ _26315_/Q _19574_/A vssd1 vssd1 vccd1 vccd1 _14611_/A sky130_fd_sc_hd__xor2_1
X_22508_ _22508_/A _22900_/B vssd1 vssd1 vccd1 vccd1 _22508_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_162_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14290_ _14344_/A hold263/X vssd1 vssd1 vccd1 vccd1 hold264/A sky130_fd_sc_hd__nand2_1
X_26276_ _26279_/CLK _26276_/D vssd1 vssd1 vccd1 vccd1 _26276_/Q sky130_fd_sc_hd__dfxtp_2
X_23488_ _24940_/S hold248/A _23487_/X vssd1 vssd1 vccd1 vccd1 _23488_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13241_ _26304_/Q _19416_/A vssd1 vssd1 vccd1 vccd1 _14575_/A sky130_fd_sc_hd__xor2_1
X_25227_ _25678_/CLK hold490/X vssd1 vssd1 vccd1 vccd1 hold488/A sky130_fd_sc_hd__dfxtp_1
X_22439_ _19774_/A _22438_/A _22438_/Y vssd1 vssd1 vccd1 vccd1 _22441_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_165_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13172_ _13049_/X _14542_/A _13067_/X _19257_/A vssd1 vssd1 vccd1 vccd1 _13172_/X
+ sky130_fd_sc_hd__a22o_1
X_25158_ _26248_/CLK hold598/X vssd1 vssd1 vccd1 vccd1 hold596/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24109_ _24109_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24110_/A sky130_fd_sc_hd__and2_1
X_17980_ _19230_/A vssd1 vssd1 vccd1 vccd1 _22190_/B sky130_fd_sc_hd__inv_2
X_25089_ _26301_/CLK _25089_/D vssd1 vssd1 vccd1 vccd1 _25089_/Q sky130_fd_sc_hd__dfxtp_1
X_16931_ _16929_/X _16711_/X _16930_/Y _25894_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16932_/A sky130_fd_sc_hd__a32o_1
X_16862_ _16862_/A _16862_/B vssd1 vssd1 vccd1 vccd1 _16862_/Y sky130_fd_sc_hd__nand2_1
X_19650_ _19648_/X _19649_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19650_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15813_ _15813_/A vssd1 vssd1 vccd1 vccd1 _16691_/A sky130_fd_sc_hd__inv_2
X_18601_ _18641_/A _19430_/A vssd1 vssd1 vccd1 vccd1 _18601_/Y sky130_fd_sc_hd__nand2_1
X_19581_ _19573_/X _19580_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19581_/Y sky130_fd_sc_hd__o21ai_1
X_16793_ _22680_/A vssd1 vssd1 vccd1 vccd1 _16935_/A sky130_fd_sc_hd__buf_6
XFILLER_0_99_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18532_ _18532_/A _20131_/A vssd1 vssd1 vccd1 vccd1 _18878_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15744_ _15744_/A vssd1 vssd1 vccd1 vccd1 _16953_/A sky130_fd_sc_hd__inv_2
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12956_ _26253_/Q _25622_/Q vssd1 vssd1 vccd1 vccd1 _14416_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_158_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _18463_/A _18463_/B vssd1 vssd1 vccd1 vccd1 _22094_/A sky130_fd_sc_hd__nand2_1
X_15675_ _15675_/A vssd1 vssd1 vccd1 vccd1 _15692_/B sky130_fd_sc_hd__inv_2
XFILLER_0_75_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _12726_/B _14373_/A _12752_/X _25609_/Q vssd1 vssd1 vccd1 vccd1 _12887_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _17624_/A _17414_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17414_/X sky130_fd_sc_hd__and3_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _14626_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14626_/Y sky130_fd_sc_hd__nand2_1
X_18394_ _18392_/X _18269_/X _18393_/X vssd1 vssd1 vccd1 vccd1 _18395_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _17345_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17345_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_56_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _14557_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14557_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13508_ _13583_/A _13508_/B vssd1 vssd1 vccd1 vccd1 _13508_/Y sky130_fd_sc_hd__nand2_1
X_17276_ _19402_/A _17276_/B vssd1 vssd1 vccd1 vccd1 _17549_/A sky130_fd_sc_hd__xor2_4
X_14488_ _14488_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14488_/Y sky130_fd_sc_hd__nand2_1
X_19015_ _19186_/A _19788_/A vssd1 vssd1 vccd1 vccd1 _19015_/Y sky130_fd_sc_hd__nand2_1
X_16227_ _16227_/A _16227_/B vssd1 vssd1 vccd1 vccd1 _16246_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_125_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13439_ _13220_/A _14675_/A _13242_/A _25705_/Q vssd1 vssd1 vccd1 vccd1 _13439_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16158_ _16158_/A _16158_/B vssd1 vssd1 vccd1 vccd1 _16272_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_144_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15109_ _15084_/B _15106_/B _15107_/A _15086_/X _15101_/A vssd1 vssd1 vccd1 vccd1
+ _15111_/A sky130_fd_sc_hd__o221a_1
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16089_ _16089_/A _16697_/B _16097_/A vssd1 vssd1 vccd1 vccd1 _16089_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_11_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2706 _24978_/Q vssd1 vssd1 vccd1 vccd1 _12621_/A sky130_fd_sc_hd__dlygate4sd3_1
X_19917_ _19975_/A _19917_/B vssd1 vssd1 vccd1 vccd1 _19917_/Y sky130_fd_sc_hd__nand2_1
Xhold2717 _25439_/Q vssd1 vssd1 vccd1 vccd1 _15169_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2728 _24572_/X vssd1 vssd1 vccd1 vccd1 _24573_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2739 _26260_/Q vssd1 vssd1 vccd1 vccd1 hold2739/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19848_ _19849_/B _19849_/A vssd1 vssd1 vccd1 vccd1 _19848_/X sky130_fd_sc_hd__or2_1
XFILLER_0_177_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19779_ _19779_/A _19779_/B vssd1 vssd1 vccd1 vccd1 _19779_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21810_ _25804_/Q _21810_/B vssd1 vssd1 vccd1 vccd1 _21810_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22790_ _22788_/X _22789_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22790_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21741_ _19430_/A _21740_/A _21740_/Y vssd1 vssd1 vccd1 vccd1 _21743_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24460_ _24460_/A vssd1 vssd1 vccd1 vccd1 _26217_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21672_ _21670_/Y _21671_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21672_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23411_ _24940_/S hold338/A _23410_/X vssd1 vssd1 vccd1 vccd1 _23411_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20623_ _20621_/Y _20622_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _20623_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24391_ hold2294/X _26195_/Q _24433_/S vssd1 vssd1 vccd1 vccd1 _24391_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_31_clk _25759_/CLK vssd1 vssd1 vccd1 vccd1 _26080_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26130_ _26130_/CLK _26130_/D vssd1 vssd1 vccd1 vccd1 hold899/A sky130_fd_sc_hd__dfxtp_1
X_23342_ _23342_/A _23342_/B vssd1 vssd1 vccd1 vccd1 _23347_/A sky130_fd_sc_hd__nand2_1
X_20554_ _20553_/B _20554_/B _20554_/C vssd1 vssd1 vccd1 vccd1 _20555_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26061_ _26065_/CLK _26061_/D vssd1 vssd1 vccd1 vccd1 _26061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23273_ _23273_/A hold829/X vssd1 vssd1 vccd1 vccd1 hold830/A sky130_fd_sc_hd__nand2_1
X_20485_ _20487_/B vssd1 vssd1 vccd1 vccd1 _20486_/B sky130_fd_sc_hd__inv_2
XFILLER_0_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25012_ _26096_/CLK _25012_/D vssd1 vssd1 vccd1 vccd1 _25012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22224_ _22224_/A _22224_/B vssd1 vssd1 vccd1 vccd1 _22225_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22155_ _22155_/A _22155_/B vssd1 vssd1 vccd1 vccd1 _22823_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_100_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21106_ _21109_/A _21109_/B vssd1 vssd1 vccd1 vccd1 _21108_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_160_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22086_ _22063_/X _22085_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _22086_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_98_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _25483_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25914_ _26341_/CLK _25914_/D vssd1 vssd1 vccd1 vccd1 _25914_/Q sky130_fd_sc_hd__dfxtp_1
X_21037_ _21037_/A _21037_/B vssd1 vssd1 vccd1 vccd1 _21038_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_121_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25845_ _26208_/CLK _25845_/D vssd1 vssd1 vccd1 vccd1 _25845_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_92_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12810_ _26097_/Q _12748_/X _12809_/X vssd1 vssd1 vccd1 vccd1 _12810_/X sky130_fd_sc_hd__a21o_1
X_25776_ _26251_/CLK _25776_/D vssd1 vssd1 vccd1 vccd1 _25776_/Q sky130_fd_sc_hd__dfxtp_1
X_13790_ _13823_/A _13790_/B vssd1 vssd1 vccd1 vccd1 _13790_/Y sky130_fd_sc_hd__nand2_1
X_22988_ _23197_/A _22988_/B vssd1 vssd1 vccd1 vccd1 _22988_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_186_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24727_ _24727_/A vssd1 vssd1 vccd1 vccd1 _26304_/D sky130_fd_sc_hd__clkbuf_1
X_12741_ _14064_/A vssd1 vssd1 vccd1 vccd1 _14125_/A sky130_fd_sc_hd__inv_6
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21939_ _18175_/A _25799_/Q _21937_/Y _21938_/Y vssd1 vssd1 vccd1 vccd1 _21940_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _15466_/A vssd1 vssd1 vccd1 vccd1 _15463_/B sky130_fd_sc_hd__inv_2
XFILLER_0_155_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _12672_/A _24836_/B _12681_/B vssd1 vssd1 vccd1 vccd1 _12672_/X sky130_fd_sc_hd__and3_1
X_24658_ hold2628/X _26282_/Q _24664_/S vssd1 vssd1 vccd1 vccd1 _24658_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14411_ _14465_/A hold407/X vssd1 vssd1 vccd1 vccd1 hold408/A sky130_fd_sc_hd__nand2_1
X_23609_ _23609_/A vssd1 vssd1 vccd1 vccd1 _25942_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15391_ _15405_/A _15392_/A vssd1 vssd1 vccd1 vccd1 _15391_/X sky130_fd_sc_hd__or2_1
XFILLER_0_38_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24589_ _24589_/A vssd1 vssd1 vccd1 vccd1 _26259_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_22_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _26281_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_170_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17130_ _25631_/Q vssd1 vssd1 vccd1 vccd1 _20401_/B sky130_fd_sc_hd__inv_2
X_26328_ _26330_/CLK _26328_/D vssd1 vssd1 vccd1 vccd1 _26328_/Q sky130_fd_sc_hd__dfxtp_2
X_14342_ _14340_/Y hold117/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold118/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17061_ _17393_/A hold988/X _19994_/B vssd1 vssd1 vccd1 vccd1 _17061_/X sky130_fd_sc_hd__and3_1
X_14273_ _22829_/A vssd1 vssd1 vccd1 vccd1 _14273_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_80_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26259_ _26273_/CLK _26259_/D vssd1 vssd1 vccd1 vccd1 _26259_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16012_ _22144_/B _16691_/B _16018_/B vssd1 vssd1 vccd1 vccd1 _16013_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_150_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13224_ _26173_/Q _13065_/X _13223_/X vssd1 vssd1 vccd1 vccd1 _13224_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_123_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13155_ _26162_/Q _13065_/X _13154_/X vssd1 vssd1 vccd1 vccd1 _13155_/X sky130_fd_sc_hd__a21o_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17963_ _18535_/A _17963_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _17963_/X sky130_fd_sc_hd__and3_1
X_13086_ _17819_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13086_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_89_clk clkbuf_leaf_95_clk/A vssd1 vssd1 vccd1 vccd1 _25510_/CLK sky130_fd_sc_hd__clkbuf_16
X_19702_ _20321_/A _22327_/B _25629_/Q vssd1 vssd1 vccd1 vccd1 _20326_/C sky130_fd_sc_hd__nand3_1
X_16914_ _16977_/A _16914_/B vssd1 vssd1 vccd1 vccd1 _16914_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17894_ _18528_/A _25722_/Q vssd1 vssd1 vccd1 vccd1 _17896_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19633_ _19649_/B _19720_/B vssd1 vssd1 vccd1 vccd1 _19635_/A sky130_fd_sc_hd__xnor2_1
X_16845_ _22866_/B _16773_/A _16841_/Y _16844_/Y _12702_/A vssd1 vssd1 vccd1 vccd1
+ _16845_/Y sky130_fd_sc_hd__a221oi_1
X_16776_ _16980_/A _16776_/B vssd1 vssd1 vccd1 vccd1 _16776_/Y sky130_fd_sc_hd__nand2_1
X_19564_ _19565_/B _19565_/A vssd1 vssd1 vccd1 vccd1 _19564_/X sky130_fd_sc_hd__or2_1
XFILLER_0_88_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13988_ _14120_/A vssd1 vssd1 vccd1 vccd1 _13988_/X sky130_fd_sc_hd__clkbuf_16
X_15727_ hold883/X _15729_/A vssd1 vssd1 vccd1 vccd1 _15731_/A sky130_fd_sc_hd__nor2_1
X_18515_ _18535_/A _18515_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18515_/X sky130_fd_sc_hd__and3_1
XFILLER_0_186_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12939_ _17457_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12939_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19495_ _19492_/X _19493_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19495_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15658_ _15658_/A vssd1 vssd1 vccd1 vccd1 _15692_/A sky130_fd_sc_hd__inv_2
XFILLER_0_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18446_ _18446_/A _25748_/Q _21716_/A vssd1 vssd1 vccd1 vccd1 _18447_/C sky130_fd_sc_hd__nand3_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14609_ _14645_/A hold23/X vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__nand2_1
XFILLER_0_139_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18377_ _18375_/Y _18376_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25663_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15589_ _15589_/A _16890_/A vssd1 vssd1 vccd1 vccd1 _15590_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _26146_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17328_ _21075_/B _25868_/Q _25804_/Q vssd1 vssd1 vccd1 vccd1 _17329_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_16_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17259_ _17272_/A _17259_/B vssd1 vssd1 vccd1 vccd1 _17259_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20270_ _20660_/A _20270_/B vssd1 vssd1 vccd1 vccd1 _20270_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_113_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2503 _18945_/Y vssd1 vssd1 vccd1 vccd1 _25691_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2514 _26196_/Q vssd1 vssd1 vccd1 vccd1 hold2514/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2525 _25438_/Q vssd1 vssd1 vccd1 vccd1 _15158_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2536 _24985_/Q vssd1 vssd1 vccd1 vccd1 _12671_/C sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2547 _23273_/A vssd1 vssd1 vccd1 vccd1 _23270_/C sky130_fd_sc_hd__dlygate4sd3_1
X_23960_ _23960_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23961_/A sky130_fd_sc_hd__and2_1
Xhold1802 _17518_/Y vssd1 vssd1 vccd1 vccd1 _25626_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1813 _25629_/Q vssd1 vssd1 vccd1 vccd1 _17539_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2558 _24529_/X vssd1 vssd1 vccd1 vccd1 _24530_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2569 _25463_/Q vssd1 vssd1 vccd1 vccd1 _15602_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1824 _25592_/Q vssd1 vssd1 vccd1 vccd1 _17164_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22911_ _23188_/A _22911_/B vssd1 vssd1 vccd1 vccd1 _22911_/X sky130_fd_sc_hd__or2_1
Xhold1835 _25843_/Q vssd1 vssd1 vccd1 vccd1 _21931_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1846 _17576_/Y vssd1 vssd1 vccd1 vccd1 _25634_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23891_ _23891_/A vssd1 vssd1 vccd1 vccd1 _26034_/D sky130_fd_sc_hd__clkbuf_1
Xhold1857 _22231_/Y vssd1 vssd1 vccd1 vccd1 _25853_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1868 _25632_/Q vssd1 vssd1 vccd1 vccd1 _17560_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1879 _22059_/Y vssd1 vssd1 vccd1 vccd1 _25847_/D sky130_fd_sc_hd__dlygate4sd3_1
X_25630_ _25716_/CLK _25630_/D vssd1 vssd1 vccd1 vccd1 _25630_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_155_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22842_ _22842_/A _22842_/B vssd1 vssd1 vccd1 vccd1 _22843_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_155_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25561_ _25878_/CLK _25561_/D vssd1 vssd1 vccd1 vccd1 _25561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22773_ _22771_/X _22772_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22773_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24512_ _24512_/A vssd1 vssd1 vccd1 vccd1 _26234_/D sky130_fd_sc_hd__clkbuf_1
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21724_ _23193_/B _22421_/A vssd1 vssd1 vccd1 vccd1 _21725_/A sky130_fd_sc_hd__or2_1
XFILLER_0_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25492_ _25925_/CLK hold802/X vssd1 vssd1 vccd1 vccd1 hold800/A sky130_fd_sc_hd__dfxtp_1
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24443_ _26211_/Q hold1997/X _24510_/S vssd1 vssd1 vccd1 vccd1 _24443_/X sky130_fd_sc_hd__mux2_1
X_21655_ _22058_/A _21655_/B vssd1 vssd1 vccd1 vccd1 _21655_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_87_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20606_ _20606_/A _20606_/B vssd1 vssd1 vccd1 vccd1 _21612_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_35_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24374_ _24374_/A vssd1 vssd1 vccd1 vccd1 _26189_/D sky130_fd_sc_hd__clkbuf_1
X_21586_ _21636_/A _21586_/B _21585_/X vssd1 vssd1 vccd1 vccd1 _21587_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_35_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26113_ _26116_/CLK _26113_/D vssd1 vssd1 vccd1 vccd1 _26113_/Q sky130_fd_sc_hd__dfxtp_1
X_23325_ _23325_/A _23377_/B _23330_/A vssd1 vssd1 vccd1 vccd1 _23325_/X sky130_fd_sc_hd__and3_1
X_20537_ _26290_/Q _20078_/X hold728/X vssd1 vssd1 vccd1 vccd1 _20540_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26044_ _26079_/CLK _26044_/D vssd1 vssd1 vccd1 vccd1 _26044_/Q sky130_fd_sc_hd__dfxtp_1
X_23256_ _23256_/A _23256_/B vssd1 vssd1 vccd1 vccd1 _23275_/B sky130_fd_sc_hd__nand2_1
X_20468_ _20468_/A _20468_/B vssd1 vssd1 vccd1 vccd1 _20472_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22207_ _22207_/A _25881_/Q vssd1 vssd1 vccd1 vccd1 _22207_/Y sky130_fd_sc_hd__nand2_1
X_23187_ _23187_/A _23187_/B vssd1 vssd1 vccd1 vccd1 _23187_/Y sky130_fd_sc_hd__nand2_1
X_20399_ _21222_/C vssd1 vssd1 vccd1 vccd1 _21225_/B sky130_fd_sc_hd__inv_2
X_22138_ _22139_/A _22139_/C _23090_/A vssd1 vssd1 vccd1 vccd1 _22138_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_24_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14960_ _14958_/X hold2207/X _14928_/X vssd1 vssd1 vccd1 vccd1 _14960_/Y sky130_fd_sc_hd__a21oi_1
X_22069_ _22789_/B _22070_/A vssd1 vssd1 vccd1 vccd1 _22071_/A sky130_fd_sc_hd__or2_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ hold684/X _13910_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold685/A sky130_fd_sc_hd__a21oi_1
X_14891_ _14900_/A _14891_/B vssd1 vssd1 vccd1 vccd1 _14891_/Y sky130_fd_sc_hd__nand2_1
X_16630_ _16630_/A vssd1 vssd1 vccd1 vccd1 _16649_/B sky130_fd_sc_hd__inv_2
X_25828_ _25838_/CLK _25828_/D vssd1 vssd1 vccd1 vccd1 _25828_/Q sky130_fd_sc_hd__dfxtp_2
X_13842_ _13941_/A _13842_/B vssd1 vssd1 vccd1 vccd1 _13842_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_187_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16561_ _16561_/A hold910/X _16691_/B vssd1 vssd1 vccd1 vccd1 _16562_/B sky130_fd_sc_hd__and3_1
X_25759_ _25759_/CLK _25759_/D vssd1 vssd1 vccd1 vccd1 _25759_/Q sky130_fd_sc_hd__dfxtp_1
X_13773_ hold405/X _13772_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold406/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15512_ hold878/X _15514_/A vssd1 vssd1 vccd1 vccd1 _15516_/A sky130_fd_sc_hd__nor2_1
X_18300_ _21102_/B _19473_/A vssd1 vssd1 vccd1 vccd1 _18301_/B sky130_fd_sc_hd__nand2_1
X_19280_ _19280_/A _19280_/B vssd1 vssd1 vccd1 vccd1 _19280_/Y sky130_fd_sc_hd__nand2_1
X_12724_ _25582_/Q _12724_/B vssd1 vssd1 vccd1 vccd1 _12724_/X sky130_fd_sc_hd__or2_1
X_16492_ _16492_/A _16492_/B vssd1 vssd1 vccd1 vccd1 _16492_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18231_ _18231_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18231_/Y sky130_fd_sc_hd__nand2_1
X_15443_ _15443_/A _15443_/B vssd1 vssd1 vccd1 vccd1 _15467_/B sky130_fd_sc_hd__or2_1
XFILLER_0_154_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12655_ _12656_/B _12656_/A vssd1 vssd1 vccd1 vccd1 _12657_/A sky130_fd_sc_hd__or2_1
XFILLER_0_127_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18162_ _19388_/A vssd1 vssd1 vccd1 vccd1 _21938_/B sky130_fd_sc_hd__inv_2
X_15374_ _15374_/A _15374_/B vssd1 vssd1 vccd1 vccd1 _15405_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_170_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12586_ _23923_/B _12587_/A vssd1 vssd1 vccd1 vccd1 _12591_/A sky130_fd_sc_hd__or2_1
XFILLER_0_167_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17113_ _17111_/Y _17112_/Y _16941_/X vssd1 vssd1 vccd1 vccd1 _17113_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14325_ _14325_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14325_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_151_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18093_ _18093_/A _18093_/B vssd1 vssd1 vccd1 vccd1 _21868_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_151_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17044_ _17623_/A _17044_/B vssd1 vssd1 vccd1 vccd1 _17044_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_52_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold409 hold409/A vssd1 vssd1 vccd1 vccd1 hold409/X sky130_fd_sc_hd__dlygate4sd3_1
X_14256_ _18936_/B _14262_/B vssd1 vssd1 vccd1 vccd1 _14256_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_150_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13207_ _14260_/A vssd1 vssd1 vccd1 vccd1 _13207_/X sky130_fd_sc_hd__buf_4
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14187_ _14182_/Y _14186_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold824/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _14064_/A vssd1 vssd1 vccd1 vccd1 _13320_/B sky130_fd_sc_hd__buf_6
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _18992_/Y _18994_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25696_/D sky130_fd_sc_hd__a21oi_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17946_ _20513_/B _22162_/A vssd1 vssd1 vccd1 vccd1 _20506_/A sky130_fd_sc_hd__nand2_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _26146_/Q _13065_/X _13068_/X vssd1 vssd1 vccd1 vccd1 _13069_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_2_clk _26093_/CLK vssd1 vssd1 vccd1 vccd1 _26122_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1109 _25060_/Q vssd1 vssd1 vccd1 vccd1 _17617_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17877_ _17877_/A _17877_/B vssd1 vssd1 vccd1 vccd1 _17878_/B sky130_fd_sc_hd__nand2_1
X_19616_ _19616_/A _20099_/B vssd1 vssd1 vccd1 vccd1 _19616_/Y sky130_fd_sc_hd__nor2_1
X_16828_ _16826_/Y _16827_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16828_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19547_ _21237_/A _22015_/B _25618_/Q vssd1 vssd1 vccd1 vccd1 _21241_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_177_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16759_ _16980_/A _16764_/B vssd1 vssd1 vccd1 vccd1 _16761_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_76_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19478_ _19478_/A _19478_/B vssd1 vssd1 vccd1 vccd1 _19478_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_119_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18429_ _18793_/A _18429_/B _18894_/C vssd1 vssd1 vccd1 vccd1 _18430_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21440_ _21439_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21440_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21371_ _21371_/A _21371_/B _21371_/C vssd1 vssd1 vccd1 vccd1 _21372_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_185_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23110_ _26079_/Q vssd1 vssd1 vccd1 vccd1 _23111_/A sky130_fd_sc_hd__inv_2
X_20322_ _20322_/A _20322_/B vssd1 vssd1 vccd1 vccd1 _20326_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24090_ _24090_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24091_/A sky130_fd_sc_hd__and2_1
Xhold910 hold910/A vssd1 vssd1 vccd1 vccd1 hold910/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 hold921/A vssd1 vssd1 vccd1 vccd1 hold921/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 hold932/A vssd1 vssd1 vccd1 vccd1 hold932/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold943 hold943/A vssd1 vssd1 vccd1 vccd1 hold943/X sky130_fd_sc_hd__dlygate4sd3_1
X_23041_ _23041_/A _23041_/B vssd1 vssd1 vccd1 vccd1 _23042_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_12_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20253_ _20254_/A _20254_/C _20254_/B vssd1 vssd1 vccd1 vccd1 _20255_/A sky130_fd_sc_hd__a21o_1
Xhold954 hold954/A vssd1 vssd1 vccd1 vccd1 hold954/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 hold965/A vssd1 vssd1 vccd1 vccd1 hold965/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 hold976/A vssd1 vssd1 vccd1 vccd1 hold976/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 hold987/A vssd1 vssd1 vccd1 vccd1 hold987/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold998 hold998/A vssd1 vssd1 vccd1 vccd1 hold998/X sky130_fd_sc_hd__dlygate4sd3_1
X_20184_ _21434_/A _21059_/C vssd1 vssd1 vccd1 vccd1 _20187_/B sky130_fd_sc_hd__nand2_1
Xhold2300 _15430_/Y vssd1 vssd1 vccd1 vccd1 hold2300/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2311 _24403_/X vssd1 vssd1 vccd1 vccd1 _24404_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2322 _26185_/Q vssd1 vssd1 vccd1 vccd1 hold2322/X sky130_fd_sc_hd__dlygate4sd3_1
X_24992_ _25491_/CLK hold998/X vssd1 vssd1 vccd1 vccd1 hold997/A sky130_fd_sc_hd__dfxtp_1
Xhold2333 _24341_/X vssd1 vssd1 vccd1 vccd1 _24342_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2344 _26206_/Q vssd1 vssd1 vccd1 vccd1 hold2344/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1610 _25827_/Q vssd1 vssd1 vccd1 vccd1 _21557_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2355 _24181_/X vssd1 vssd1 vccd1 vccd1 _24182_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2366 _26336_/Q vssd1 vssd1 vccd1 vccd1 hold2366/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1621 _17461_/Y vssd1 vssd1 vccd1 vccd1 _25618_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23943_ _23943_/A vssd1 vssd1 vccd1 vccd1 _26049_/D sky130_fd_sc_hd__clkbuf_1
Xhold1632 _25645_/Q vssd1 vssd1 vccd1 vccd1 _17656_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2377 _25658_/Q vssd1 vssd1 vccd1 vccd1 _13146_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2388 _25669_/Q vssd1 vssd1 vccd1 vccd1 _13214_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1643 hold2754/X vssd1 vssd1 vccd1 vccd1 _18147_/B sky130_fd_sc_hd__clkbuf_2
Xhold2399 _15378_/Y vssd1 vssd1 vccd1 vccd1 hold2399/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1654 _20348_/Y vssd1 vssd1 vccd1 vccd1 _25782_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1665 _25764_/Q vssd1 vssd1 vccd1 vccd1 _19891_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1676 _25885_/Q vssd1 vssd1 vccd1 vccd1 _22937_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23874_ hold2130/X hold2240/X _23907_/S vssd1 vssd1 vccd1 vccd1 _23875_/A sky130_fd_sc_hd__mux2_1
Xhold1687 _25641_/Q vssd1 vssd1 vccd1 vccd1 _17627_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1698 _25609_/Q vssd1 vssd1 vccd1 vccd1 _17376_/B sky130_fd_sc_hd__dlygate4sd3_1
X_25613_ _26117_/CLK _25613_/D vssd1 vssd1 vccd1 vccd1 _25613_/Q sky130_fd_sc_hd__dfxtp_2
X_22825_ _22825_/A _22825_/B vssd1 vssd1 vccd1 vccd1 _22826_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25544_ _26047_/CLK _25544_/D vssd1 vssd1 vccd1 vccd1 _25544_/Q sky130_fd_sc_hd__dfxtp_1
X_22756_ _22937_/A _22756_/B vssd1 vssd1 vccd1 vccd1 _22756_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21707_ _21707_/A _21707_/B _21707_/C vssd1 vssd1 vccd1 vccd1 _21711_/A sky130_fd_sc_hd__nand3_1
X_25475_ _25535_/CLK _25475_/D vssd1 vssd1 vccd1 vccd1 _25475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22687_ _22687_/A _22900_/B vssd1 vssd1 vccd1 vccd1 _22687_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_81_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24426_ _24426_/A vssd1 vssd1 vccd1 vccd1 _26206_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21638_ _21638_/A _22902_/B vssd1 vssd1 vccd1 vccd1 _21638_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_180_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24357_ _24357_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24358_/A sky130_fd_sc_hd__and2_1
X_21569_ _21568_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21569_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14110_ _14180_/A _14110_/B vssd1 vssd1 vccd1 vccd1 _14110_/Y sky130_fd_sc_hd__nand2_1
X_23308_ _23310_/B _23310_/A vssd1 vssd1 vccd1 vccd1 _23317_/A sky130_fd_sc_hd__nor2_1
X_15090_ _15464_/A vssd1 vssd1 vccd1 vccd1 _15090_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24288_ _24288_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24289_/A sky130_fd_sc_hd__and2_1
XFILLER_0_132_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26027_ _26042_/CLK _26027_/D vssd1 vssd1 vccd1 vccd1 _26027_/Q sky130_fd_sc_hd__dfxtp_1
X_14041_ _18224_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14041_/Y sky130_fd_sc_hd__nor2_1
X_23239_ _23237_/X hold2678/X _12702_/A vssd1 vssd1 vccd1 vccd1 _23239_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17800_ _18529_/A _17800_/B _18083_/C vssd1 vssd1 vccd1 vccd1 _17801_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_24_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15992_ _15990_/X hold772/X _15805_/X vssd1 vssd1 vccd1 vccd1 hold773/A sky130_fd_sc_hd__a21oi_1
X_18780_ _18778_/X _18269_/X _18779_/X vssd1 vssd1 vccd1 vccd1 _18781_/A sky130_fd_sc_hd__a21o_1
X_14943_ _14941_/X hold2204/X _14928_/X vssd1 vssd1 vccd1 vccd1 _14943_/Y sky130_fd_sc_hd__a21oi_1
X_17731_ _17764_/B _17699_/B _17699_/A vssd1 vssd1 vccd1 vccd1 _17734_/B sky130_fd_sc_hd__a21boi_1
X_14874_ _14872_/Y _14873_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14874_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17662_ _17662_/A _17662_/B _20025_/A vssd1 vssd1 vccd1 vccd1 _17667_/A sky130_fd_sc_hd__and3_2
X_19401_ _19398_/Y _19401_/B _19980_/B vssd1 vssd1 vccd1 vccd1 _19401_/X sky130_fd_sc_hd__and3b_1
X_16613_ _16698_/A hold871/X vssd1 vssd1 vccd1 vccd1 _16613_/Y sky130_fd_sc_hd__nand2_1
X_13825_ _13880_/A hold659/X vssd1 vssd1 vccd1 vccd1 hold660/A sky130_fd_sc_hd__nand2_1
X_17593_ _17593_/A _17644_/A vssd1 vssd1 vccd1 vccd1 _17594_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16544_ _16598_/B vssd1 vssd1 vccd1 vccd1 _16545_/B sky130_fd_sc_hd__inv_2
X_19332_ _20817_/A _21801_/B _25603_/Q vssd1 vssd1 vccd1 vccd1 _20822_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_168_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13756_ _18612_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13756_/Y sky130_fd_sc_hd__nor2_1
X_12707_ hold2010/X _12707_/B vssd1 vssd1 vccd1 vccd1 _12707_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_35_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16475_ _16676_/A _16475_/B vssd1 vssd1 vccd1 vccd1 _16477_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19263_ _19262_/Y _21228_/A _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _19265_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13687_ _13760_/A hold401/X vssd1 vssd1 vccd1 vccd1 hold402/A sky130_fd_sc_hd__nand2_1
X_15426_ _15426_/A _15426_/B vssd1 vssd1 vccd1 vccd1 _15427_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_54_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18214_ _19416_/A vssd1 vssd1 vccd1 vccd1 _22006_/B sky130_fd_sc_hd__inv_2
XFILLER_0_182_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12638_ _12654_/C _12654_/A vssd1 vssd1 vccd1 vccd1 _12640_/A sky130_fd_sc_hd__or2_1
XFILLER_0_26_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19194_ _26218_/Q _19483_/A hold530/X vssd1 vssd1 vccd1 vccd1 _19195_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15357_ _15357_/A _15357_/B vssd1 vssd1 vccd1 vccd1 _15406_/C sky130_fd_sc_hd__nor2_1
X_18145_ _18143_/X _17528_/X _18144_/X vssd1 vssd1 vccd1 vccd1 _18146_/A sky130_fd_sc_hd__a21o_1
X_12569_ _12575_/A vssd1 vssd1 vccd1 vccd1 _12574_/A sky130_fd_sc_hd__inv_2
XFILLER_0_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14308_ _14344_/A hold278/X vssd1 vssd1 vccd1 vccd1 hold279/A sky130_fd_sc_hd__nand2_1
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18076_ _18076_/A _20247_/A vssd1 vssd1 vccd1 vccd1 _19060_/A sky130_fd_sc_hd__xnor2_4
X_15288_ _16294_/A _16711_/A vssd1 vssd1 vccd1 vccd1 _15290_/A sky130_fd_sc_hd__nand2_1
Xhold206 hold206/A vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 hold217/A vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 hold228/A vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
X_17027_ _17413_/A _17498_/A vssd1 vssd1 vccd1 vccd1 _17028_/B sky130_fd_sc_hd__xnor2_1
X_14239_ _26336_/Q _13518_/B _14170_/X _14238_/Y vssd1 vssd1 vccd1 vccd1 _14240_/B
+ sky130_fd_sc_hd__a22o_1
Xhold239 hold239/A vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18978_ _18978_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _18978_/Y sky130_fd_sc_hd__nand2_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _17931_/A vssd1 vssd1 vccd1 vccd1 _17930_/A sky130_fd_sc_hd__inv_2
X_20940_ _20940_/A _21943_/B _20940_/C vssd1 vssd1 vccd1 vccd1 _20944_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_117_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20871_ _20871_/A _21400_/C _20871_/C vssd1 vssd1 vccd1 vccd1 _20872_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_152_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22610_ _22610_/A _22900_/B vssd1 vssd1 vccd1 vccd1 _22610_/Y sky130_fd_sc_hd__nand2_1
X_23590_ _23590_/A _23590_/B vssd1 vssd1 vccd1 vccd1 _23592_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_14_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22541_ _22541_/A _22541_/B vssd1 vssd1 vccd1 vccd1 _22541_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_76_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25260_ _26046_/CLK _25260_/D vssd1 vssd1 vccd1 vccd1 _25260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22472_ _22875_/A _23024_/B vssd1 vssd1 vccd1 vccd1 _22473_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24211_ _24211_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24212_/A sky130_fd_sc_hd__and2_1
XFILLER_0_162_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21423_ _26322_/Q hold825/X vssd1 vssd1 vccd1 vccd1 _21423_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25191_ _25770_/CLK hold682/X vssd1 vssd1 vccd1 vccd1 hold680/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24142_ hold2336/X hold2323/X _24203_/S vssd1 vssd1 vccd1 vccd1 _24143_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21354_ _21354_/A _21354_/B _21354_/C vssd1 vssd1 vccd1 vccd1 _21355_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_124_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20305_ _20305_/A _20305_/B vssd1 vssd1 vccd1 vccd1 _20306_/A sky130_fd_sc_hd__nand2_1
X_24073_ _24073_/A vssd1 vssd1 vccd1 vccd1 _26091_/D sky130_fd_sc_hd__clkbuf_1
Xhold740 hold740/A vssd1 vssd1 vccd1 vccd1 hold740/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21285_ _21636_/A _21285_/B _21284_/X vssd1 vssd1 vccd1 vccd1 _21286_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold751 hold751/A vssd1 vssd1 vccd1 vccd1 hold751/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 hold762/A vssd1 vssd1 vccd1 vccd1 hold762/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 hold773/A vssd1 vssd1 vccd1 vccd1 hold773/X sky130_fd_sc_hd__dlygate4sd3_1
X_23024_ _23170_/A _23024_/B vssd1 vssd1 vccd1 vccd1 _23025_/B sky130_fd_sc_hd__nand2_1
X_20236_ _20236_/A _20236_/B vssd1 vssd1 vccd1 vccd1 _20240_/A sky130_fd_sc_hd__nand2_1
Xhold784 hold784/A vssd1 vssd1 vccd1 vccd1 hold784/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 hold795/A vssd1 vssd1 vccd1 vccd1 hold795/X sky130_fd_sc_hd__dlygate4sd3_1
X_20167_ _20167_/A _20167_/B _20167_/C vssd1 vssd1 vccd1 vccd1 _20171_/C sky130_fd_sc_hd__nand3_1
Xhold2130 _26028_/Q vssd1 vssd1 vccd1 vccd1 hold2130/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2141 _23616_/X vssd1 vssd1 vccd1 vccd1 _23617_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2152 _23373_/X vssd1 vssd1 vccd1 vccd1 _23374_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24975_ _25420_/CLK hold870/X vssd1 vssd1 vccd1 vccd1 hold868/A sky130_fd_sc_hd__dfxtp_1
Xhold2163 _25969_/Q vssd1 vssd1 vccd1 vccd1 hold2163/X sky130_fd_sc_hd__dlygate4sd3_1
X_20098_ _20098_/A _22149_/B vssd1 vssd1 vccd1 vccd1 _20099_/A sky130_fd_sc_hd__nand2_1
Xhold2174 _23321_/X vssd1 vssd1 vccd1 vccd1 _23322_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2185 _26095_/Q vssd1 vssd1 vccd1 vccd1 hold2185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1440 _13028_/X vssd1 vssd1 vccd1 vccd1 _25055_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1451 _25057_/Q vssd1 vssd1 vccd1 vccd1 _17595_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2196 _15015_/A vssd1 vssd1 vccd1 vccd1 _15010_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23926_ _23598_/B _23924_/Y _23925_/X _12515_/X vssd1 vssd1 vccd1 vccd1 _23927_/A
+ sky130_fd_sc_hd__a211o_2
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1462 _19513_/Y vssd1 vssd1 vccd1 vccd1 _25737_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1473 _25092_/Q vssd1 vssd1 vccd1 vccd1 _18557_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1484 _19976_/Y vssd1 vssd1 vccd1 vccd1 _25771_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1495 _25053_/Q vssd1 vssd1 vccd1 vccd1 _17564_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23857_ _23857_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23858_/A sky130_fd_sc_hd__and2_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ hold642/X _13609_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold643/A sky130_fd_sc_hd__a21oi_1
X_22808_ _22808_/A _23120_/B vssd1 vssd1 vccd1 vccd1 _22809_/B sky130_fd_sc_hd__nand2_1
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _14590_/A vssd1 vssd1 vccd1 vccd1 _14645_/A sky130_fd_sc_hd__clkbuf_8
X_23788_ _14866_/B _14875_/B _23831_/S vssd1 vssd1 vccd1 vccd1 _23789_/A sky130_fd_sc_hd__mux2_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25527_ _25533_/CLK _25527_/D vssd1 vssd1 vccd1 vccd1 _25527_/Q sky130_fd_sc_hd__dfxtp_1
X_13541_ hold459/X _13540_/Y _12558_/B vssd1 vssd1 vccd1 vccd1 hold460/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22739_ _22730_/Y _22738_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22739_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_55_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16260_ _16260_/A _16401_/C vssd1 vssd1 vccd1 vccd1 _16262_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_165_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25458_ _26064_/CLK hold879/X vssd1 vssd1 vccd1 vccd1 hold878/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ _13583_/A _13472_/B vssd1 vssd1 vccd1 vccd1 _13472_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ _16235_/A _16711_/A vssd1 vssd1 vccd1 vccd1 _16747_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_164_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24409_ hold2321/X hold2276/X _24433_/S vssd1 vssd1 vccd1 vccd1 _24410_/A sky130_fd_sc_hd__mux2_1
X_16191_ hold882/X vssd1 vssd1 vccd1 vccd1 _16195_/B sky130_fd_sc_hd__inv_2
XFILLER_0_152_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25389_ _25859_/CLK _25389_/D vssd1 vssd1 vccd1 vccd1 _25389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15142_ _16179_/A _16711_/A vssd1 vssd1 vccd1 vccd1 _16719_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_164_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15073_ _15073_/A _15085_/A vssd1 vssd1 vccd1 vccd1 _15073_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_132_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19950_ _19950_/A _19950_/B vssd1 vssd1 vccd1 vccd1 _19950_/Y sky130_fd_sc_hd__nand2_1
X_14024_ _14061_/A _14024_/B vssd1 vssd1 vccd1 vccd1 _14024_/Y sky130_fd_sc_hd__nand2_1
X_18901_ _18899_/X _18879_/X _18900_/X vssd1 vssd1 vccd1 vccd1 _18902_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19881_ _19880_/Y _19130_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19883_/A
+ sky130_fd_sc_hd__a211o_1
X_18832_ _18954_/A _25767_/Q vssd1 vssd1 vccd1 vccd1 _18834_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18763_ _18761_/Y _18762_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25682_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15975_ _15975_/A vssd1 vssd1 vccd1 vccd1 _15975_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_175_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17714_ _17722_/A _17717_/A _17750_/B vssd1 vssd1 vccd1 vccd1 _17726_/A sky130_fd_sc_hd__nand3_1
X_14926_ _14927_/B _14927_/A vssd1 vssd1 vccd1 vccd1 _14926_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18694_ _18694_/A _18694_/B _18694_/C vssd1 vssd1 vccd1 vccd1 _22393_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17645_ _17645_/A _17645_/B vssd1 vssd1 vccd1 vccd1 _17645_/X sky130_fd_sc_hd__xor2_1
X_14857_ _14850_/Y _14856_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14857_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ _25764_/Q vssd1 vssd1 vccd1 vccd1 _18773_/B sky130_fd_sc_hd__inv_2
XFILLER_0_187_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14788_ _15839_/A _14788_/B vssd1 vssd1 vccd1 vccd1 _22061_/A sky130_fd_sc_hd__nand2_1
X_17576_ _17574_/Y _17575_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _17576_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19315_ _19314_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19316_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16527_ _16541_/A _16528_/A vssd1 vssd1 vccd1 vccd1 _16529_/A sky130_fd_sc_hd__or2_1
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13739_ _26256_/Q _13612_/X _13605_/X _13738_/Y vssd1 vssd1 vccd1 vccd1 _13740_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19246_ _20585_/A _19244_/Y _20590_/C vssd1 vssd1 vccd1 vccd1 _19336_/B sky130_fd_sc_hd__o21a_2
X_16458_ _16473_/A hold935/X vssd1 vssd1 vccd1 vccd1 _16458_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15409_ _15389_/A _15372_/A _15388_/A vssd1 vssd1 vccd1 vccd1 _15409_/X sky130_fd_sc_hd__a21o_1
X_16389_ _16389_/A vssd1 vssd1 vccd1 vccd1 _16404_/B sky130_fd_sc_hd__inv_2
XFILLER_0_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19177_ _19177_/A _21924_/A _25587_/Q vssd1 vssd1 vccd1 vccd1 _20214_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_143_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18128_ _19017_/A vssd1 vssd1 vccd1 vccd1 _19067_/A sky130_fd_sc_hd__inv_2
XFILLER_0_171_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18059_ _18057_/X _17528_/X _18058_/X vssd1 vssd1 vccd1 vccd1 _18060_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_1_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21070_ _21070_/A _21070_/B vssd1 vssd1 vccd1 vccd1 _21071_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_112_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20021_ _21370_/A vssd1 vssd1 vccd1 vccd1 _21369_/A sky130_fd_sc_hd__inv_2
XFILLER_0_158_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24760_ _26314_/Q hold2644/X _24817_/S vssd1 vssd1 vccd1 vccd1 _24760_/X sky130_fd_sc_hd__mux2_1
X_21972_ _25800_/Q _21972_/B vssd1 vssd1 vccd1 vccd1 _21972_/Y sky130_fd_sc_hd__nor2_1
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23711_ hold2045/X hold2018/X _23754_/S vssd1 vssd1 vccd1 vccd1 _23712_/A sky130_fd_sc_hd__mux2_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20923_ _21709_/A _21483_/B vssd1 vssd1 vccd1 vccd1 _20924_/C sky130_fd_sc_hd__nand2_1
X_24691_ _24691_/A vssd1 vssd1 vccd1 vccd1 _26292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23642_ _23642_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23643_/A sky130_fd_sc_hd__and2_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20854_ _20852_/Y _20853_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _20854_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_166_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23573_ _24922_/S hold317/A _23572_/X vssd1 vssd1 vccd1 vccd1 _23573_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20785_ _20787_/B _20787_/C vssd1 vssd1 vccd1 vccd1 _20786_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25312_ _26139_/CLK hold58/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22524_ _23184_/A _22524_/B vssd1 vssd1 vccd1 vccd1 _22525_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_91_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26292_ _26292_/CLK _26292_/D vssd1 vssd1 vccd1 vccd1 _26292_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_161_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25243_ _25709_/CLK hold700/X vssd1 vssd1 vccd1 vccd1 hold698/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22455_ _22453_/A _22454_/X _22453_/B vssd1 vssd1 vccd1 vccd1 _22456_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21406_ _26321_/Q _21228_/X hold434/X vssd1 vssd1 vccd1 vccd1 _21409_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_162_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25174_ _25174_/CLK hold586/X vssd1 vssd1 vccd1 vccd1 hold584/A sky130_fd_sc_hd__dfxtp_1
X_22386_ _22653_/A _22386_/B vssd1 vssd1 vccd1 vccd1 _22386_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24125_ _24125_/A vssd1 vssd1 vccd1 vccd1 _26108_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21337_ _21691_/C _21386_/A vssd1 vssd1 vccd1 vccd1 _21338_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_130_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24056_ hold2277/X hold2239/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24057_/A sky130_fd_sc_hd__mux2_1
Xhold570 hold570/A vssd1 vssd1 vccd1 vccd1 hold570/X sky130_fd_sc_hd__dlygate4sd3_1
X_21268_ _25875_/Q _21268_/B _21268_/C vssd1 vssd1 vccd1 vccd1 _21271_/C sky130_fd_sc_hd__nand3b_1
Xhold581 hold581/A vssd1 vssd1 vccd1 vccd1 hold581/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 hold592/A vssd1 vssd1 vccd1 vccd1 hold592/X sky130_fd_sc_hd__dlygate4sd3_1
X_23007_ _23007_/A _23007_/B vssd1 vssd1 vccd1 vccd1 _23009_/A sky130_fd_sc_hd__nand2_1
X_20219_ _21086_/C vssd1 vssd1 vccd1 vccd1 _21089_/B sky130_fd_sc_hd__inv_2
XFILLER_0_60_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21199_ _21199_/A _21199_/B vssd1 vssd1 vccd1 vccd1 _21200_/A sky130_fd_sc_hd__nand2_1
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15760_ _15760_/A vssd1 vssd1 vccd1 vccd1 _15762_/A sky130_fd_sc_hd__inv_2
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24958_ _24958_/A _24958_/B vssd1 vssd1 vccd1 vccd1 _24958_/Y sky130_fd_sc_hd__nand2_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _12891_/X _14425_/A _12909_/X _25625_/Q vssd1 vssd1 vccd1 vccd1 _12972_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1270 _25039_/Q vssd1 vssd1 vccd1 vccd1 _17464_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ _14711_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14711_/Y sky130_fd_sc_hd__nand2_1
Xhold1281 _13187_/X vssd1 vssd1 vccd1 vccd1 _25084_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15691_ _15691_/A _15691_/B vssd1 vssd1 vccd1 vccd1 _15718_/A sky130_fd_sc_hd__nand2_1
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23909_ _23909_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23910_/A sky130_fd_sc_hd__and2_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1292 _25018_/Q vssd1 vssd1 vccd1 vccd1 _17242_/B sky130_fd_sc_hd__dlygate4sd3_1
X_24889_ _24889_/A _24957_/S vssd1 vssd1 vccd1 vccd1 _24889_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_169_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _14645_/A hold467/X vssd1 vssd1 vccd1 vccd1 hold468/A sky130_fd_sc_hd__nand2_1
X_17430_ _25622_/Q vssd1 vssd1 vccd1 vccd1 _20055_/B sky130_fd_sc_hd__inv_2
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17361_ _17549_/A _17601_/A vssd1 vssd1 vccd1 vccd1 _17362_/B sky130_fd_sc_hd__xnor2_1
X_14573_ _14585_/A hold176/X vssd1 vssd1 vccd1 vccd1 hold177/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19100_ _19950_/B _19211_/B vssd1 vssd1 vccd1 vccd1 _19101_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16312_ _16313_/B _16313_/A vssd1 vssd1 vccd1 vccd1 _16314_/A sky130_fd_sc_hd__or2_1
XFILLER_0_138_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13524_ _14120_/A vssd1 vssd1 vccd1 vccd1 _13638_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17292_ _20000_/B _25899_/Q _25835_/Q vssd1 vssd1 vccd1 vccd1 _17293_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_153_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16243_ _16241_/X _16242_/Y _16076_/X vssd1 vssd1 vccd1 vccd1 _25505_/D sky130_fd_sc_hd__a21oi_1
X_19031_ _19031_/A _19081_/A vssd1 vssd1 vccd1 vccd1 _19032_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13455_ _26211_/Q _13426_/X _13454_/X vssd1 vssd1 vccd1 vccd1 _13455_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_180_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16174_ _16171_/A _16171_/B _16189_/B _16173_/Y vssd1 vssd1 vccd1 vccd1 _16174_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13386_ _26199_/Q _13239_/X _13385_/X vssd1 vssd1 vccd1 vccd1 _13386_/X sky130_fd_sc_hd__a21o_1
X_15125_ _14266_/A _12527_/A _22829_/A vssd1 vssd1 vccd1 vccd1 _16660_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15056_ _15054_/X _15055_/Y _14928_/X vssd1 vssd1 vccd1 vccd1 _25430_/D sky130_fd_sc_hd__a21oi_1
X_19933_ _26271_/Q hold626/X vssd1 vssd1 vccd1 vccd1 _19933_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_107_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14007_ _14125_/A vssd1 vssd1 vccd1 vccd1 _14118_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19864_ _19857_/X _19863_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19864_/Y sky130_fd_sc_hd__o21ai_1
X_18815_ _20681_/B _22541_/A vssd1 vssd1 vccd1 vccd1 _20672_/A sky130_fd_sc_hd__nand2_2
X_19795_ _19787_/X _19794_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19795_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_170_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18746_ _20558_/B _19788_/A vssd1 vssd1 vccd1 vccd1 _18747_/B sky130_fd_sc_hd__nand2_1
X_15958_ _22035_/B _16691_/B hold929/X vssd1 vssd1 vccd1 vccd1 _15960_/A sky130_fd_sc_hd__a21o_1
X_14909_ _14909_/A _14909_/B vssd1 vssd1 vccd1 vccd1 _14917_/A sky130_fd_sc_hd__nand2_1
X_18677_ _18878_/A _18981_/A vssd1 vssd1 vccd1 vccd1 _18678_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15889_ _21864_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _15891_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17628_ _17626_/Y _17627_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _25641_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17559_ _17559_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17559_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_50_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20570_ _21595_/A _21319_/C vssd1 vssd1 vccd1 vccd1 _20571_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_34_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19229_ _19227_/Y hold938/X _19086_/X vssd1 vssd1 vccd1 vccd1 hold939/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22240_ _19659_/A _22239_/A _22239_/Y vssd1 vssd1 vccd1 vccd1 _22242_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22171_ _22561_/A _22171_/B vssd1 vssd1 vccd1 vccd1 _22171_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_48_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21122_ _21121_/Y _20192_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21122_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_160_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25930_ _25939_/CLK _25930_/D vssd1 vssd1 vccd1 vccd1 _25930_/Q sky130_fd_sc_hd__dfxtp_1
X_21053_ _21053_/A _21053_/B vssd1 vssd1 vccd1 vccd1 _21055_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20004_ _20004_/A _25899_/Q _20004_/C vssd1 vssd1 vccd1 vccd1 _20007_/C sky130_fd_sc_hd__nand3_1
X_25861_ _25865_/CLK _25861_/D vssd1 vssd1 vccd1 vccd1 _25861_/Q sky130_fd_sc_hd__dfxtp_2
X_24812_ _24812_/A _24833_/B vssd1 vssd1 vccd1 vccd1 _24813_/A sky130_fd_sc_hd__and2_1
X_25792_ _25793_/CLK _25792_/D vssd1 vssd1 vccd1 vccd1 _25792_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_154_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24743_ _24743_/A vssd1 vssd1 vccd1 vccd1 _24817_/S sky130_fd_sc_hd__clkbuf_16
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21955_ _22703_/A vssd1 vssd1 vccd1 vccd1 _22216_/A sky130_fd_sc_hd__inv_2
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20906_ _21235_/A _20906_/B vssd1 vssd1 vccd1 vccd1 _20906_/Y sky130_fd_sc_hd__nand2_1
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24674_ hold2591/X hold2485/X _24740_/S vssd1 vssd1 vccd1 vccd1 _24675_/A sky130_fd_sc_hd__mux2_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21886_ _22651_/A vssd1 vssd1 vccd1 vccd1 _22157_/A sky130_fd_sc_hd__inv_2
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23625_ _25947_/Q hold2101/X _23677_/S vssd1 vssd1 vccd1 vccd1 _23625_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_65_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20837_ _20837_/A _20837_/B vssd1 vssd1 vccd1 vccd1 _21709_/B sky130_fd_sc_hd__nand2_8
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23556_ hold152/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23556_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20768_ _20768_/A _20768_/B vssd1 vssd1 vccd1 vccd1 _20770_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22507_ _16729_/B _22421_/X _22501_/X _22502_/Y _22506_/X vssd1 vssd1 vccd1 vccd1
+ _22508_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_174_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26275_ _26275_/CLK _26275_/D vssd1 vssd1 vccd1 vccd1 _26275_/Q sky130_fd_sc_hd__dfxtp_1
X_23487_ hold134/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23487_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_165_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20699_ _21235_/A _20699_/B vssd1 vssd1 vccd1 vccd1 _20699_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_107_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13240_ _13240_/A vssd1 vssd1 vccd1 vccd1 _19416_/A sky130_fd_sc_hd__buf_4
X_25226_ _25678_/CLK hold697/X vssd1 vssd1 vccd1 vccd1 hold695/A sky130_fd_sc_hd__dfxtp_1
X_22438_ _22438_/A _22438_/B vssd1 vssd1 vccd1 vccd1 _22438_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_150_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13171_ _26293_/Q _19257_/A vssd1 vssd1 vccd1 vccd1 _14542_/A sky130_fd_sc_hd__xor2_1
X_25157_ _26248_/CLK hold836/X vssd1 vssd1 vccd1 vccd1 hold835/A sky130_fd_sc_hd__dfxtp_1
X_22369_ _22369_/A _25887_/Q vssd1 vssd1 vccd1 vccd1 _22369_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24108_ hold2351/X hold2034/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24109_/A sky130_fd_sc_hd__mux2_1
X_25088_ _26301_/CLK _25088_/D vssd1 vssd1 vccd1 vccd1 _25088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16930_ _16930_/A _16930_/B vssd1 vssd1 vccd1 vccd1 _16930_/Y sky130_fd_sc_hd__nand2_1
X_24039_ _24039_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24040_/A sky130_fd_sc_hd__and2_1
X_16861_ _16862_/B _16862_/A vssd1 vssd1 vccd1 vccd1 _16861_/X sky130_fd_sc_hd__or2_1
X_18600_ _18600_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18600_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_189_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15812_ _23188_/B _15812_/B vssd1 vssd1 vccd1 vccd1 _15813_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_176_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19580_ _19578_/X _19579_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19580_/Y sky130_fd_sc_hd__a21oi_1
X_16792_ _16789_/Y _16790_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16792_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18531_ _20139_/C _22181_/A vssd1 vssd1 vccd1 vccd1 _20131_/A sky130_fd_sc_hd__nand2_2
X_15743_ _15743_/A vssd1 vssd1 vccd1 vccd1 _15745_/A sky130_fd_sc_hd__inv_2
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12955_ _12930_/X _12953_/X _12917_/X _12954_/X vssd1 vssd1 vccd1 vccd1 _12955_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18462_ _20011_/B _19588_/A vssd1 vssd1 vccd1 vccd1 _18463_/B sky130_fd_sc_hd__nand2_1
X_15674_ _15674_/A _15674_/B vssd1 vssd1 vccd1 vccd1 _15675_/A sky130_fd_sc_hd__nor2_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _26240_/Q _25609_/Q vssd1 vssd1 vccd1 vccd1 _14373_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_59_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17413_ _17413_/A _17413_/B vssd1 vssd1 vccd1 vccd1 _17413_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_96_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14625_ _14623_/Y hold471/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold472/A sky130_fd_sc_hd__a21oi_1
X_18393_ _18535_/A _18393_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _18393_/X sky130_fd_sc_hd__and3_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17344_ _17342_/X _17241_/X _17343_/X vssd1 vssd1 vccd1 vccd1 _17345_/A sky130_fd_sc_hd__a21o_1
X_14556_ _14554_/Y hold375/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold376/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13507_ _26219_/Q _13426_/X _13468_/X _13506_/Y vssd1 vssd1 vccd1 vccd1 _13508_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17275_ _20965_/B _25864_/Q _20991_/B vssd1 vssd1 vccd1 vccd1 _17276_/B sky130_fd_sc_hd__mux2_2
X_14487_ _14485_/Y hold312/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold313/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19014_ _19014_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _19014_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16226_ _16228_/B vssd1 vssd1 vccd1 vccd1 _16245_/B sky130_fd_sc_hd__inv_2
X_13438_ _26336_/Q _25705_/Q vssd1 vssd1 vccd1 vccd1 _14675_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_3_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16157_ _16161_/B _16157_/B vssd1 vssd1 vccd1 vccd1 _16158_/A sky130_fd_sc_hd__and2_1
XFILLER_0_140_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13369_ _18968_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13369_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15108_ _15108_/A _15110_/B vssd1 vssd1 vccd1 vccd1 _15269_/B sky130_fd_sc_hd__and2_1
X_16088_ _16088_/A _16088_/B vssd1 vssd1 vccd1 vccd1 _16097_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_80_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15039_ _15270_/A _15051_/A vssd1 vssd1 vccd1 vccd1 _15039_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19916_ _19909_/X _19915_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19916_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2707 _26256_/Q vssd1 vssd1 vccd1 vccd1 hold2707/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2718 _26283_/Q vssd1 vssd1 vccd1 vccd1 hold2718/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2729 _26233_/Q vssd1 vssd1 vccd1 vccd1 hold2729/X sky130_fd_sc_hd__dlygate4sd3_1
X_19847_ _19862_/B _19928_/B vssd1 vssd1 vccd1 vccd1 _19849_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19778_ _19779_/B _19779_/A vssd1 vssd1 vccd1 vccd1 _19778_/X sky130_fd_sc_hd__or2_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18729_ _18792_/A _18733_/B vssd1 vssd1 vccd1 vccd1 _18731_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21740_ _21740_/A _21740_/B vssd1 vssd1 vccd1 vccd1 _21740_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21671_ _22058_/A _21671_/B vssd1 vssd1 vccd1 vccd1 _21671_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23410_ hold26/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23410_/X sky130_fd_sc_hd__or2b_1
X_20622_ _20660_/A _20622_/B vssd1 vssd1 vccd1 vccd1 _20622_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24390_ _24390_/A vssd1 vssd1 vccd1 vccd1 _26194_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23341_ _23342_/B _23342_/A vssd1 vssd1 vccd1 vccd1 _23343_/A sky130_fd_sc_hd__or2_1
XFILLER_0_144_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20553_ _20553_/A _20553_/B vssd1 vssd1 vccd1 vccd1 _20555_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26060_ _26060_/CLK _26060_/D vssd1 vssd1 vccd1 vccd1 _26060_/Q sky130_fd_sc_hd__dfxtp_1
X_23272_ hold829/X _23273_/A vssd1 vssd1 vccd1 vccd1 _23272_/X sky130_fd_sc_hd__or2_1
X_20484_ _20487_/A _20487_/C vssd1 vssd1 vccd1 vccd1 _20486_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_132_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25011_ _26096_/CLK _25011_/D vssd1 vssd1 vccd1 vccd1 _25011_/Q sky130_fd_sc_hd__dfxtp_1
X_22223_ _22224_/B _22224_/A vssd1 vssd1 vccd1 vccd1 _22225_/A sky130_fd_sc_hd__or2_2
XFILLER_0_104_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22154_ _22154_/A _22838_/B vssd1 vssd1 vccd1 vccd1 _22155_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_113_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21105_ _25869_/Q _21105_/B _21105_/C vssd1 vssd1 vccd1 vccd1 _21109_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_22_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22085_ _22083_/X _22084_/Y _21789_/X vssd1 vssd1 vccd1 vccd1 _22085_/Y sky130_fd_sc_hd__a21oi_2
Xclkbuf_4_1__f_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_clk/A
+ sky130_fd_sc_hd__clkbuf_16
X_25913_ _25913_/CLK _25913_/D vssd1 vssd1 vccd1 vccd1 _25913_/Q sky130_fd_sc_hd__dfxtp_1
X_21036_ _21036_/A _21036_/B _21036_/C vssd1 vssd1 vccd1 vccd1 _21037_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_22_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25844_ _25859_/CLK _25844_/D vssd1 vssd1 vccd1 vccd1 _25844_/Q sky130_fd_sc_hd__dfxtp_4
X_22987_ _22978_/Y _22986_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22987_/X sky130_fd_sc_hd__a21o_1
X_25775_ _26251_/CLK _25775_/D vssd1 vssd1 vccd1 vccd1 _25775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12740_ _16711_/A _16773_/A vssd1 vssd1 vccd1 vccd1 _14064_/A sky130_fd_sc_hd__nor2_8
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21938_ _25799_/Q _21938_/B vssd1 vssd1 vccd1 vccd1 _21938_/Y sky130_fd_sc_hd__nor2_1
X_24726_ _24726_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24727_/A sky130_fd_sc_hd__and2_1
XFILLER_0_96_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12671_ _12662_/C _12671_/B _12671_/C vssd1 vssd1 vccd1 vccd1 _12681_/B sky130_fd_sc_hd__nand3b_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24657_ _24657_/A vssd1 vssd1 vccd1 vccd1 _26281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21869_ _25797_/Q _21869_/B vssd1 vssd1 vccd1 vccd1 _21869_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14590_/A vssd1 vssd1 vccd1 vccd1 _14465_/A sky130_fd_sc_hd__clkbuf_8
X_23608_ _23608_/A _23629_/B vssd1 vssd1 vccd1 vccd1 _23609_/A sky130_fd_sc_hd__and2_1
XFILLER_0_139_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15390_ _15378_/A _15374_/B _15372_/A vssd1 vssd1 vccd1 vccd1 _15392_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24588_ _24588_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24589_/A sky130_fd_sc_hd__and2_1
XFILLER_0_181_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14341_ _14344_/A hold116/X vssd1 vssd1 vccd1 vccd1 hold117/A sky130_fd_sc_hd__nand2_1
X_26327_ _26330_/CLK _26327_/D vssd1 vssd1 vccd1 vccd1 _26327_/Q sky130_fd_sc_hd__dfxtp_2
X_23539_ _24942_/S hold293/A _23538_/X vssd1 vssd1 vccd1 vccd1 _23539_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17060_ _17630_/A _17060_/B vssd1 vssd1 vccd1 vccd1 _17060_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_107_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14272_ _14277_/B _14277_/C _23629_/B _14271_/Y vssd1 vssd1 vccd1 vccd1 _25258_/D
+ sky130_fd_sc_hd__o211a_1
X_26258_ _26264_/CLK _26258_/D vssd1 vssd1 vccd1 vccd1 _26258_/Q sky130_fd_sc_hd__dfxtp_4
X_16011_ _16011_/A _16676_/A _22144_/B vssd1 vssd1 vccd1 vccd1 _16028_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25209_ _26292_/CLK hold854/X vssd1 vssd1 vccd1 vccd1 hold853/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13223_ _13220_/X _14566_/A _13067_/X _19373_/A vssd1 vssd1 vccd1 vccd1 _13223_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26189_ _26190_/CLK _26189_/D vssd1 vssd1 vccd1 vccd1 _26189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13154_ _13049_/X _14533_/A _13067_/X _19216_/A vssd1 vssd1 vccd1 vccd1 _13154_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _19039_/A _17962_/B vssd1 vssd1 vccd1 vccd1 _17962_/X sky130_fd_sc_hd__xor2_1
X_13085_ _26149_/Q _13065_/X _13084_/X vssd1 vssd1 vccd1 vccd1 _13085_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_97_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19701_ _19701_/A _20322_/B vssd1 vssd1 vccd1 vccd1 _19701_/Y sky130_fd_sc_hd__nor2_1
X_16913_ _16913_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16913_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_100_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17893_ _17893_/A _25786_/Q _17893_/C vssd1 vssd1 vccd1 vccd1 _20474_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_109_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19632_ _20131_/A _19630_/Y _20135_/C vssd1 vssd1 vccd1 vccd1 _19720_/B sky130_fd_sc_hd__o21a_2
X_16844_ _16842_/Y _15458_/A _16843_/Y vssd1 vssd1 vccd1 vccd1 _16844_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19563_ _19579_/B _19649_/B vssd1 vssd1 vccd1 vccd1 _19565_/A sky130_fd_sc_hd__xnor2_1
X_16775_ _25871_/Q _13468_/X _16774_/Y vssd1 vssd1 vccd1 vccd1 _16775_/Y sky130_fd_sc_hd__a21oi_1
X_13987_ _14000_/A hold656/X vssd1 vssd1 vccd1 vccd1 hold657/A sky130_fd_sc_hd__nand2_1
X_18514_ _18514_/A _18514_/B vssd1 vssd1 vccd1 vccd1 _18514_/X sky130_fd_sc_hd__xor2_1
X_15726_ _15795_/A _16625_/B vssd1 vssd1 vccd1 vccd1 _15729_/A sky130_fd_sc_hd__nor2_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _26121_/Q _12907_/X _12937_/X vssd1 vssd1 vccd1 vccd1 _12938_/X sky130_fd_sc_hd__a21o_1
X_19494_ _21789_/A vssd1 vssd1 vccd1 vccd1 _19494_/X sky130_fd_sc_hd__buf_6
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18445_ _18445_/A _18449_/B vssd1 vssd1 vccd1 vccd1 _18447_/A sky130_fd_sc_hd__nand2_1
X_15657_ _15657_/A _15657_/B vssd1 vssd1 vccd1 vccd1 _15658_/A sky130_fd_sc_hd__nor2_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ hold983/X _12974_/B vssd1 vssd1 vccd1 vccd1 _12869_/X sky130_fd_sc_hd__or2_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14608_ _14608_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14608_/Y sky130_fd_sc_hd__nand2_1
X_18376_ _18641_/A _19275_/A vssd1 vssd1 vccd1 vccd1 _18376_/Y sky130_fd_sc_hd__nand2_1
X_15588_ _15588_/A vssd1 vssd1 vccd1 vccd1 _16890_/A sky130_fd_sc_hd__inv_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17327_ _25612_/Q vssd1 vssd1 vccd1 vccd1 _21075_/B sky130_fd_sc_hd__inv_2
X_14539_ _14539_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14539_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17258_ _17258_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17258_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_183_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16209_ _16214_/B _16210_/A vssd1 vssd1 vccd1 vccd1 _16209_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17189_ _17189_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17189_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2504 _26058_/Q vssd1 vssd1 vccd1 vccd1 hold2504/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2515 _25683_/Q vssd1 vssd1 vccd1 vccd1 _13303_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2526 _15180_/X vssd1 vssd1 vccd1 vccd1 _15182_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2537 _12674_/B vssd1 vssd1 vccd1 vccd1 _12667_/C sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1803 hold2759/X vssd1 vssd1 vccd1 vccd1 _17685_/C sky130_fd_sc_hd__buf_1
Xhold2548 _25688_/Q vssd1 vssd1 vccd1 vccd1 _13335_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2559 _26230_/Q vssd1 vssd1 vccd1 vccd1 hold2559/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1814 _17540_/Y vssd1 vssd1 vccd1 vccd1 _25629_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1825 _25856_/Q vssd1 vssd1 vccd1 vccd1 _22320_/B sky130_fd_sc_hd__dlygate4sd3_1
X_22910_ _22910_/A _23027_/B vssd1 vssd1 vccd1 vccd1 _22910_/Y sky130_fd_sc_hd__nand2_1
Xhold1836 _21932_/Y vssd1 vssd1 vccd1 vccd1 _25843_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23890_ _23890_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23891_/A sky130_fd_sc_hd__and2_1
Xhold1847 _25914_/Q vssd1 vssd1 vccd1 vccd1 _23581_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1858 _25857_/Q vssd1 vssd1 vccd1 vccd1 _22341_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1869 _17561_/Y vssd1 vssd1 vccd1 vccd1 _25632_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22841_ _22841_/A _23152_/B vssd1 vssd1 vccd1 vccd1 _22842_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25560_ _26065_/CLK _25560_/D vssd1 vssd1 vccd1 vccd1 _25560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22772_ _22937_/A _22772_/B vssd1 vssd1 vccd1 vccd1 _22772_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_149_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24511_ _24511_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24512_/A sky130_fd_sc_hd__and2_1
XFILLER_0_17_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21723_ _14267_/A _24871_/B _21203_/A vssd1 vssd1 vccd1 vccd1 _22421_/A sky130_fd_sc_hd__a21o_4
XFILLER_0_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25491_ _25491_/CLK hold706/X vssd1 vssd1 vccd1 vccd1 hold704/A sky130_fd_sc_hd__dfxtp_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24442_ _24442_/A vssd1 vssd1 vccd1 vccd1 _26211_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21654_ _21654_/A _22902_/B vssd1 vssd1 vccd1 vccd1 _21654_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20605_ _20605_/A _20605_/B _20605_/C vssd1 vssd1 vccd1 vccd1 _20606_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_164_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24373_ _24373_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24374_/A sky130_fd_sc_hd__and2_1
X_21585_ _21584_/Y _21203_/X _20986_/X _20957_/A vssd1 vssd1 vccd1 vccd1 _21585_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_35_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26112_ _26112_/CLK _26112_/D vssd1 vssd1 vccd1 vccd1 _26112_/Q sky130_fd_sc_hd__dfxtp_1
X_23324_ _23324_/A _23324_/B vssd1 vssd1 vccd1 vccd1 _23330_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20536_ _20536_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20541_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26043_ _26073_/CLK _26043_/D vssd1 vssd1 vccd1 vccd1 _26043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23255_ _23255_/A vssd1 vssd1 vccd1 vccd1 _23256_/B sky130_fd_sc_hd__inv_2
XFILLER_0_162_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20467_ _20467_/A _22131_/B vssd1 vssd1 vccd1 vccd1 _20468_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_162_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22206_ _22206_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _22206_/X sky130_fd_sc_hd__and2_1
XFILLER_0_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23186_ _23186_/A _23186_/B vssd1 vssd1 vccd1 vccd1 _23187_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20398_ _20398_/A _20398_/B vssd1 vssd1 vccd1 vccd1 _21222_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_63_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22137_ _22137_/A _22137_/B vssd1 vssd1 vccd1 vccd1 _23090_/A sky130_fd_sc_hd__nand2_8
X_22068_ _19574_/A _22067_/A _22067_/Y vssd1 vssd1 vccd1 vccd1 _22070_/A sky130_fd_sc_hd__o21ai_2
X_21019_ _21235_/A _21019_/B vssd1 vssd1 vccd1 vccd1 _21019_/Y sky130_fd_sc_hd__nand2_1
X_13910_ _13941_/A _13910_/B vssd1 vssd1 vccd1 vccd1 _13910_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14890_ _14890_/A _14899_/B vssd1 vssd1 vccd1 vccd1 _14890_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_173_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25827_ _25827_/CLK _25827_/D vssd1 vssd1 vccd1 vccd1 _25827_/Q sky130_fd_sc_hd__dfxtp_4
X_13841_ _26272_/Q _13801_/X _13793_/X _13840_/Y vssd1 vssd1 vccd1 vccd1 _13842_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16560_ _16561_/A _16691_/B hold910/X vssd1 vssd1 vccd1 vccd1 _16562_/A sky130_fd_sc_hd__a21oi_1
X_13772_ _13823_/A _13772_/B vssd1 vssd1 vccd1 vccd1 _13772_/Y sky130_fd_sc_hd__nand2_1
X_25758_ _25773_/CLK _25758_/D vssd1 vssd1 vccd1 vccd1 _25758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15511_ _15621_/A _16464_/B vssd1 vssd1 vccd1 vccd1 _15514_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_167_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24709_ _24709_/A vssd1 vssd1 vccd1 vccd1 _26298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12723_ _12529_/Y _17009_/B _12721_/Y _20023_/B vssd1 vssd1 vccd1 vccd1 _12723_/X
+ sky130_fd_sc_hd__a31o_1
X_16491_ _16491_/A _16491_/B vssd1 vssd1 vccd1 vccd1 _16491_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25689_ _25689_/CLK _25689_/D vssd1 vssd1 vccd1 vccd1 _25689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18230_ _18228_/X _17528_/X _18229_/X vssd1 vssd1 vccd1 vccd1 _18231_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_183_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15442_ _15442_/A _15442_/B vssd1 vssd1 vccd1 vccd1 _15466_/B sky130_fd_sc_hd__nor2_1
X_12654_ _12654_/A _12654_/B _12654_/C vssd1 vssd1 vccd1 vccd1 _12656_/A sky130_fd_sc_hd__and3_1
XFILLER_0_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18161_ _18161_/A _20309_/A vssd1 vssd1 vccd1 vccd1 _19074_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_81_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15373_ _16810_/A _15373_/B vssd1 vssd1 vccd1 vccd1 _15374_/B sky130_fd_sc_hd__nand2_1
X_12585_ _12585_/A vssd1 vssd1 vccd1 vccd1 _23923_/B sky130_fd_sc_hd__inv_2
XFILLER_0_65_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17112_ _17272_/A _17112_/B vssd1 vssd1 vccd1 vccd1 _17112_/Y sky130_fd_sc_hd__nand2_1
X_14324_ _14322_/Y hold282/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold283/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18092_ _20883_/B _19359_/A vssd1 vssd1 vccd1 vccd1 _18093_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14255_ _25836_/Q vssd1 vssd1 vccd1 vccd1 _18936_/B sky130_fd_sc_hd__inv_2
X_17043_ _17423_/A _17505_/A vssd1 vssd1 vccd1 vccd1 _17044_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13206_ _13109_/X _13204_/X _13192_/X _13205_/X vssd1 vssd1 vccd1 vccd1 _13206_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14186_ _14264_/A _14186_/B vssd1 vssd1 vccd1 vccd1 _14186_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_110_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _26159_/Q _13065_/X _13136_/X vssd1 vssd1 vccd1 vccd1 _13137_/X sky130_fd_sc_hd__a21o_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18994_ _19186_/A _19744_/A vssd1 vssd1 vccd1 vccd1 _18994_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _17945_/A _17945_/B _17945_/C vssd1 vssd1 vccd1 vccd1 _22162_/A sky130_fd_sc_hd__nand3_2
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _13049_/X _14482_/A _13067_/X _25643_/Q vssd1 vssd1 vccd1 vccd1 _13068_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17876_ _17877_/B _17877_/A vssd1 vssd1 vccd1 vccd1 _17878_/A sky130_fd_sc_hd__or2_1
X_19615_ _19612_/Y _19615_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19615_/X sky130_fd_sc_hd__and3b_1
X_16827_ _16858_/A _16827_/B vssd1 vssd1 vccd1 vccd1 _16827_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_177_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19546_ _19546_/A _21238_/B vssd1 vssd1 vccd1 vccd1 _19546_/Y sky130_fd_sc_hd__nor2_1
X_16758_ _16756_/Y _16757_/Y _16594_/X vssd1 vssd1 vccd1 vccd1 _16758_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_177_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15709_ _15709_/A vssd1 vssd1 vccd1 vccd1 _16617_/A sky130_fd_sc_hd__inv_2
X_19477_ _19478_/B _19478_/A vssd1 vssd1 vccd1 vccd1 _19477_/X sky130_fd_sc_hd__or2_1
X_16689_ _16695_/A _16695_/B vssd1 vssd1 vccd1 vccd1 _16694_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18428_ _18792_/A _25747_/Q vssd1 vssd1 vccd1 vccd1 _18430_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_158_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18359_ _21947_/B _25616_/Q vssd1 vssd1 vccd1 vccd1 _18361_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21370_ _21370_/A _21418_/A vssd1 vssd1 vccd1 vccd1 _21371_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20321_ _20321_/A _22327_/B vssd1 vssd1 vccd1 vccd1 _20322_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_142_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold900 hold900/A vssd1 vssd1 vccd1 vccd1 hold900/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 hold911/A vssd1 vssd1 vccd1 vccd1 hold911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 hold922/A vssd1 vssd1 vccd1 vccd1 hold922/X sky130_fd_sc_hd__dlygate4sd3_1
X_23040_ _23186_/A _23040_/B vssd1 vssd1 vccd1 vccd1 _23041_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_101_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold933 hold933/A vssd1 vssd1 vccd1 vccd1 hold933/X sky130_fd_sc_hd__dlygate4sd3_1
X_20252_ _20252_/A vssd1 vssd1 vccd1 vccd1 _20254_/B sky130_fd_sc_hd__inv_2
Xhold944 hold944/A vssd1 vssd1 vccd1 vccd1 hold944/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 hold955/A vssd1 vssd1 vccd1 vccd1 hold955/X sky130_fd_sc_hd__buf_1
XFILLER_0_12_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold966 hold966/A vssd1 vssd1 vccd1 vccd1 hold966/X sky130_fd_sc_hd__buf_1
Xhold977 hold977/A vssd1 vssd1 vccd1 vccd1 hold977/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold988 hold988/A vssd1 vssd1 vccd1 vccd1 hold988/X sky130_fd_sc_hd__dlygate4sd3_1
X_20183_ _21433_/A _21062_/B vssd1 vssd1 vccd1 vccd1 _20187_/A sky130_fd_sc_hd__nand2_1
Xhold999 hold999/A vssd1 vssd1 vccd1 vccd1 hold999/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2301 _15431_/Y vssd1 vssd1 vccd1 vccd1 _25453_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2312 _26142_/Q vssd1 vssd1 vccd1 vccd1 hold2312/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2323 _26114_/Q vssd1 vssd1 vccd1 vccd1 hold2323/X sky130_fd_sc_hd__dlygate4sd3_1
X_24991_ _25491_/CLK _24991_/D vssd1 vssd1 vccd1 vccd1 _24991_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2334 _26180_/Q vssd1 vssd1 vccd1 vccd1 hold2334/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1600 _25899_/Q vssd1 vssd1 vccd1 vccd1 _23165_/B sky130_fd_sc_hd__clkbuf_2
Xhold2345 _25667_/Q vssd1 vssd1 vccd1 vccd1 _13201_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1611 _21558_/Y vssd1 vssd1 vccd1 vccd1 _25827_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2356 _25690_/Q vssd1 vssd1 vccd1 vccd1 _13347_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23942_ _23942_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23943_/A sky130_fd_sc_hd__and2_1
Xhold2367 _24826_/X vssd1 vssd1 vccd1 vccd1 _24827_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1622 _25651_/Q vssd1 vssd1 vccd1 vccd1 _19176_/A sky130_fd_sc_hd__buf_2
Xhold2378 _25673_/Q vssd1 vssd1 vccd1 vccd1 _13240_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1633 _17657_/Y vssd1 vssd1 vccd1 vccd1 _25645_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2389 _26079_/Q vssd1 vssd1 vccd1 vccd1 hold2389/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1644 _25642_/Q vssd1 vssd1 vccd1 vccd1 _17635_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1655 _25877_/Q vssd1 vssd1 vccd1 vccd1 _22805_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23873_ _23873_/A vssd1 vssd1 vccd1 vccd1 _26028_/D sky130_fd_sc_hd__clkbuf_1
Xhold1666 _19892_/Y vssd1 vssd1 vccd1 vccd1 _25764_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1677 _22938_/Y vssd1 vssd1 vccd1 vccd1 _25885_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1688 _25599_/Q vssd1 vssd1 vccd1 vccd1 _17259_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1699 _17377_/Y vssd1 vssd1 vccd1 vccd1 _25609_/D sky130_fd_sc_hd__dlygate4sd3_1
X_22824_ _22824_/A _23136_/B vssd1 vssd1 vccd1 vccd1 _22825_/B sky130_fd_sc_hd__nand2_1
X_25612_ _26117_/CLK _25612_/D vssd1 vssd1 vccd1 vccd1 _25612_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_184_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25543_ _26047_/CLK _25543_/D vssd1 vssd1 vccd1 vccd1 _25543_/Q sky130_fd_sc_hd__dfxtp_1
X_22755_ _22746_/Y _22754_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22755_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_165_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21706_ _21708_/A _21709_/B vssd1 vssd1 vccd1 vccd1 _21707_/B sky130_fd_sc_hd__nand2_1
X_25474_ _25535_/CLK hold903/X vssd1 vssd1 vccd1 vccd1 hold902/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22686_ _16776_/B _22421_/X _22679_/X _22681_/Y _22685_/X vssd1 vssd1 vccd1 vccd1
+ _22687_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_82_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24425_ _24425_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24426_/A sky130_fd_sc_hd__and2_1
XFILLER_0_137_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21637_ _21637_/A _21637_/B vssd1 vssd1 vccd1 vccd1 _21638_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_180_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24356_ hold2491/X hold2265/X _24356_/S vssd1 vssd1 vccd1 vccd1 _24357_/A sky130_fd_sc_hd__mux2_1
X_21568_ _26331_/Q hold473/X vssd1 vssd1 vccd1 vccd1 _21568_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_105_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23307_ _23307_/A _23307_/B vssd1 vssd1 vccd1 vccd1 _23310_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20519_ _20522_/A _20522_/C vssd1 vssd1 vccd1 vccd1 _20520_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_105_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24287_ hold1909/X _26161_/Q _24356_/S vssd1 vssd1 vccd1 vccd1 _24287_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_160_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21499_ _21499_/A _21547_/A vssd1 vssd1 vccd1 vccd1 _21500_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14040_ _25801_/Q vssd1 vssd1 vccd1 vccd1 _18224_/B sky130_fd_sc_hd__inv_2
X_23238_ _23238_/A _24949_/S vssd1 vssd1 vccd1 vccd1 _23238_/Y sky130_fd_sc_hd__nand2_1
X_26026_ _26042_/CLK _26026_/D vssd1 vssd1 vccd1 vccd1 _26026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23169_ _23169_/A _23169_/B vssd1 vssd1 vccd1 vccd1 _23170_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_101_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15991_ _16212_/A hold771/X vssd1 vssd1 vccd1 vccd1 hold772/A sky130_fd_sc_hd__nand2_1
X_17730_ _17734_/A _17794_/A vssd1 vssd1 vccd1 vccd1 _17733_/A sky130_fd_sc_hd__nand2_1
X_14942_ _14942_/A _14947_/B vssd1 vssd1 vccd1 vccd1 _14942_/Y sky130_fd_sc_hd__nand2_1
X_17661_ _25838_/Q vssd1 vssd1 vccd1 vccd1 _20025_/A sky130_fd_sc_hd__inv_2
X_14873_ _14900_/A _14873_/B vssd1 vssd1 vccd1 vccd1 _14873_/Y sky130_fd_sc_hd__nand2_1
X_19400_ _19399_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19401_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16612_ _16610_/B _16610_/A _16611_/Y vssd1 vssd1 vccd1 vccd1 _16612_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_159_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13824_ hold804/X _13823_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold805/A sky130_fd_sc_hd__a21oi_1
X_17592_ _17590_/Y _17591_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _25636_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19331_ _19331_/A _20818_/B vssd1 vssd1 vccd1 vccd1 _19331_/Y sky130_fd_sc_hd__nor2_1
X_16543_ _16543_/A _16543_/B vssd1 vssd1 vccd1 vccd1 _16598_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13755_ _25756_/Q vssd1 vssd1 vccd1 vccd1 _18612_/B sky130_fd_sc_hd__inv_2
XFILLER_0_168_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12706_ hold837/X _12702_/B _12705_/X vssd1 vssd1 vccd1 vccd1 hold838/A sky130_fd_sc_hd__o21a_1
XFILLER_0_155_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19262_ _26223_/Q hold509/X vssd1 vssd1 vccd1 vccd1 _19262_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16474_ _16472_/X _16473_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 hold971/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13686_ hold615/X _13685_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold616/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18213_ _18211_/Y _18212_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25655_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15425_ _16831_/A _15425_/B vssd1 vssd1 vccd1 vccd1 _15426_/B sky130_fd_sc_hd__and2_1
XFILLER_0_156_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12637_ _12637_/A vssd1 vssd1 vccd1 vccd1 _24980_/D sky130_fd_sc_hd__clkbuf_1
X_19193_ _19192_/Y _21228_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19195_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18144_ _18535_/A _18144_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _18144_/X sky130_fd_sc_hd__and3_1
X_15356_ _16803_/A _15356_/B vssd1 vssd1 vccd1 vccd1 _15357_/B sky130_fd_sc_hd__and2_1
X_12568_ _23598_/A _12570_/A vssd1 vssd1 vccd1 vccd1 _12575_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_53_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14307_ _14307_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14307_/Y sky130_fd_sc_hd__nand2_1
X_18075_ _18075_/A _20252_/A vssd1 vssd1 vccd1 vccd1 _20247_/A sky130_fd_sc_hd__nand2_2
X_15287_ _15287_/A vssd1 vssd1 vccd1 vccd1 _16294_/A sky130_fd_sc_hd__inv_2
X_12499_ _24997_/Q vssd1 vssd1 vccd1 vccd1 _21203_/A sky130_fd_sc_hd__buf_8
XFILLER_0_123_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold207 hold207/A vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 hold218/A vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold229 hold229/A vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
X_17026_ _19630_/A _17026_/B vssd1 vssd1 vccd1 vccd1 _17498_/A sky130_fd_sc_hd__xor2_4
X_14238_ _18874_/B _14262_/B vssd1 vssd1 vccd1 vccd1 _14238_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_123_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14169_ _14236_/A hold440/X vssd1 vssd1 vccd1 vccd1 hold441/A sky130_fd_sc_hd__nand2_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ _18975_/X _18879_/X _18976_/X vssd1 vssd1 vccd1 vccd1 _18978_/A sky130_fd_sc_hd__a21o_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17928_ _17928_/A _17928_/B vssd1 vssd1 vccd1 vccd1 _17931_/A sky130_fd_sc_hd__nand2_1
X_17859_ _17859_/A _17859_/B _17859_/C vssd1 vssd1 vccd1 vccd1 _17860_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_117_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20870_ _21677_/A _21451_/B vssd1 vssd1 vccd1 vccd1 _20871_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_117_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19529_ _26242_/Q hold416/X vssd1 vssd1 vccd1 vccd1 _19529_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22540_ _18816_/A _25830_/Q _22538_/Y _22539_/Y vssd1 vssd1 vccd1 vccd1 _22541_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22471_ _23023_/A _22874_/B vssd1 vssd1 vccd1 vccd1 _22473_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24210_ hold2280/X hold2001/X _24279_/S vssd1 vssd1 vccd1 vccd1 _24211_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_106_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21422_ _26322_/Q _21228_/X hold825/X vssd1 vssd1 vccd1 vccd1 _21425_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25190_ _26273_/CLK hold782/X vssd1 vssd1 vccd1 vccd1 hold780/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24141_ _24141_/A vssd1 vssd1 vccd1 vccd1 _26113_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21353_ _21707_/C _21402_/A vssd1 vssd1 vccd1 vccd1 _21354_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_31_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20304_ _21042_/A _20304_/B _20303_/X vssd1 vssd1 vccd1 vccd1 _20305_/B sky130_fd_sc_hd__or3b_1
X_24072_ _24072_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24073_/A sky130_fd_sc_hd__and2_1
Xhold730 hold730/A vssd1 vssd1 vccd1 vccd1 hold730/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21284_ _21283_/Y _21203_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21284_/X
+ sky130_fd_sc_hd__a211o_1
Xhold741 hold741/A vssd1 vssd1 vccd1 vccd1 hold741/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold752 hold752/A vssd1 vssd1 vccd1 vccd1 hold752/X sky130_fd_sc_hd__dlygate4sd3_1
X_23023_ _23023_/A _23023_/B vssd1 vssd1 vccd1 vccd1 _23025_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold763 hold763/A vssd1 vssd1 vccd1 vccd1 hold763/X sky130_fd_sc_hd__dlygate4sd3_1
X_20235_ _20235_/A _22267_/B vssd1 vssd1 vccd1 vccd1 _20236_/A sky130_fd_sc_hd__nand2_1
Xhold774 hold774/A vssd1 vssd1 vccd1 vccd1 hold774/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 hold785/A vssd1 vssd1 vccd1 vccd1 hold785/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold796 hold796/A vssd1 vssd1 vccd1 vccd1 hold796/X sky130_fd_sc_hd__buf_1
X_20166_ _25881_/Q vssd1 vssd1 vccd1 vccd1 _20167_/B sky130_fd_sc_hd__inv_2
Xhold2120 _26015_/Q vssd1 vssd1 vccd1 vccd1 hold2120/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2131 _23871_/X vssd1 vssd1 vccd1 vccd1 _23872_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2142 _25986_/Q vssd1 vssd1 vccd1 vccd1 _14743_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2153 _26148_/Q vssd1 vssd1 vccd1 vccd1 hold2153/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24974_ _25420_/CLK _24974_/D vssd1 vssd1 vccd1 vccd1 _24974_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2164 _26091_/Q vssd1 vssd1 vccd1 vccd1 hold2164/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20097_ _21709_/A vssd1 vssd1 vccd1 vccd1 _21708_/A sky130_fd_sc_hd__inv_2
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2175 _26168_/Q vssd1 vssd1 vccd1 vccd1 hold2175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1430 _20907_/Y vssd1 vssd1 vccd1 vccd1 _25797_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2186 _25968_/Q vssd1 vssd1 vccd1 vccd1 hold2186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 _25806_/Q vssd1 vssd1 vccd1 vccd1 _21154_/B sky130_fd_sc_hd__buf_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2197 _15010_/Y vssd1 vssd1 vccd1 vccd1 hold2197/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23925_ _23924_/Y _23599_/A _24969_/Q _23924_/C vssd1 vssd1 vccd1 vccd1 _23925_/X
+ sky130_fd_sc_hd__o2bb2a_1
Xhold1452 _13038_/X vssd1 vssd1 vccd1 vccd1 _25057_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1463 _25731_/Q vssd1 vssd1 vccd1 vccd1 _19424_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1474 _13238_/X vssd1 vssd1 vccd1 vccd1 _25092_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1485 _25897_/Q vssd1 vssd1 vccd1 vccd1 _23133_/B sky130_fd_sc_hd__buf_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1496 _13017_/X vssd1 vssd1 vccd1 vccd1 _25053_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23856_ hold2039/X hold1907/X _23907_/S vssd1 vssd1 vccd1 vccd1 _23857_/A sky130_fd_sc_hd__mux2_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22807_ _23119_/B _22807_/B vssd1 vssd1 vccd1 vccd1 _22809_/A sky130_fd_sc_hd__nand2_1
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23787_ _23787_/A vssd1 vssd1 vccd1 vccd1 _26000_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20999_ _21002_/A _21002_/C vssd1 vssd1 vccd1 vccd1 _21001_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25526_ _25533_/CLK hold865/X vssd1 vssd1 vccd1 vccd1 hold864/A sky130_fd_sc_hd__dfxtp_1
X_13540_ _13583_/A _13540_/B vssd1 vssd1 vccd1 vccd1 _13540_/Y sky130_fd_sc_hd__nand2_1
X_22738_ _22738_/A _22900_/B vssd1 vssd1 vccd1 vccd1 _22738_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13471_ _26213_/Q _13426_/X _13468_/X _13470_/Y vssd1 vssd1 vccd1 vccd1 _13472_/B
+ sky130_fd_sc_hd__a22o_1
X_25457_ _26064_/CLK _25457_/D vssd1 vssd1 vccd1 vccd1 _25457_/Q sky130_fd_sc_hd__dfxtp_1
X_22669_ _22670_/B _22670_/A vssd1 vssd1 vccd1 vccd1 _22671_/A sky130_fd_sc_hd__or2_1
XFILLER_0_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15210_ _15210_/A vssd1 vssd1 vccd1 vccd1 _16235_/A sky130_fd_sc_hd__inv_2
X_24408_ _24408_/A vssd1 vssd1 vccd1 vccd1 _26200_/D sky130_fd_sc_hd__clkbuf_1
X_16190_ _16216_/A _16215_/A vssd1 vssd1 vccd1 vccd1 _16190_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_164_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25388_ _26339_/CLK hold277/X vssd1 vssd1 vccd1 vccd1 hold275/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15141_ _15141_/A vssd1 vssd1 vccd1 vccd1 _16179_/A sky130_fd_sc_hd__inv_2
XFILLER_0_51_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24339_ _24339_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24340_/A sky130_fd_sc_hd__and2_1
XFILLER_0_105_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15072_ _15085_/A _15073_/A vssd1 vssd1 vccd1 vccd1 _15072_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14023_ _26301_/Q _13988_/X _13981_/X _14022_/Y vssd1 vssd1 vccd1 vccd1 _14024_/B
+ sky130_fd_sc_hd__a22o_1
X_18900_ _19026_/A _18900_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18900_/X sky130_fd_sc_hd__and3_1
X_26009_ _26009_/CLK _26009_/D vssd1 vssd1 vccd1 vccd1 _26009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19880_ _26267_/Q hold944/X vssd1 vssd1 vccd1 vccd1 _19880_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_120_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18831_ _18831_/A _25831_/Q _18831_/C vssd1 vssd1 vccd1 vccd1 _20720_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_175_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18762_ _18986_/A _19546_/A vssd1 vssd1 vccd1 vccd1 _18762_/Y sky130_fd_sc_hd__nand2_1
X_15974_ _15961_/B _16000_/A _15960_/B vssd1 vssd1 vccd1 vccd1 _15975_/A sky130_fd_sc_hd__o21ai_1
X_17713_ _17719_/A _17719_/B vssd1 vssd1 vccd1 vccd1 _17722_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_175_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14925_ _14925_/A _14925_/B vssd1 vssd1 vccd1 vccd1 _14927_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18693_ _18793_/A _18693_/B _18894_/C vssd1 vssd1 vccd1 vccd1 _18694_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
X_17644_ _17644_/A _17644_/B vssd1 vssd1 vccd1 vccd1 _17645_/B sky130_fd_sc_hd__xnor2_1
X_14856_ _14864_/A _14856_/B vssd1 vssd1 vccd1 vccd1 _14856_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13807_ _13880_/A hold944/X vssd1 vssd1 vccd1 vccd1 _13807_/Y sky130_fd_sc_hd__nand2_1
X_17575_ _17605_/A _17575_/B vssd1 vssd1 vccd1 vccd1 _17575_/Y sky130_fd_sc_hd__nand2_1
X_14787_ _14785_/Y _14786_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14787_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19314_ _26227_/Q hold446/X vssd1 vssd1 vccd1 vccd1 _19314_/Y sky130_fd_sc_hd__nand2_1
X_16526_ _16599_/A _16543_/B _16525_/Y vssd1 vssd1 vccd1 vccd1 _16528_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_133_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13738_ _18550_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13738_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19245_ _20585_/A _22219_/B _25597_/Q vssd1 vssd1 vccd1 vccd1 _20590_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16457_ _16455_/X _16456_/Y _16231_/A vssd1 vssd1 vccd1 vccd1 _16457_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_128_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13669_ _25742_/Q vssd1 vssd1 vccd1 vccd1 _18327_/B sky130_fd_sc_hd__inv_2
XFILLER_0_171_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15408_ _15408_/A _15408_/B vssd1 vssd1 vccd1 vccd1 _15411_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19176_ _19176_/A _19176_/B vssd1 vssd1 vccd1 vccd1 _19176_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_182_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16388_ _16390_/B _16390_/A vssd1 vssd1 vccd1 vccd1 _16389_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18127_ _18127_/A _20284_/A vssd1 vssd1 vccd1 vccd1 _19017_/A sky130_fd_sc_hd__xor2_4
X_15339_ hold975/X vssd1 vssd1 vccd1 vccd1 _15341_/A sky130_fd_sc_hd__inv_2
XFILLER_0_182_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18058_ _18535_/A _18058_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _18058_/X sky130_fd_sc_hd__and3_1
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17009_ _17009_/A _17009_/B vssd1 vssd1 vccd1 vccd1 _23199_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20020_ _21676_/A _21370_/A vssd1 vssd1 vccd1 vccd1 _20028_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21971_ _21971_/A _25864_/Q vssd1 vssd1 vccd1 vccd1 _21971_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_174_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23710_ _23710_/A vssd1 vssd1 vccd1 vccd1 _25975_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20922_ _21708_/A _21480_/C vssd1 vssd1 vccd1 vccd1 _20924_/A sky130_fd_sc_hd__nand2_1
X_24690_ _24690_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24691_/A sky130_fd_sc_hd__and2_1
XFILLER_0_174_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23641_ hold2188/X hold2118/X _23677_/S vssd1 vssd1 vccd1 vccd1 _23642_/A sky130_fd_sc_hd__mux2_1
X_20853_ _21235_/A _20853_/B vssd1 vssd1 vccd1 vccd1 _20853_/Y sky130_fd_sc_hd__nand2_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23572_ hold275/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23572_/X sky130_fd_sc_hd__or2b_1
X_20784_ _20784_/A _21769_/B _20784_/C vssd1 vssd1 vccd1 vccd1 _20787_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22523_ _22523_/A _22523_/B vssd1 vssd1 vccd1 vccd1 _22524_/B sky130_fd_sc_hd__nand2_1
X_25311_ _26139_/CLK hold274/X vssd1 vssd1 vccd1 vccd1 hold272/A sky130_fd_sc_hd__dfxtp_1
X_26291_ _26292_/CLK _26291_/D vssd1 vssd1 vccd1 vccd1 _26291_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_9_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22454_ _23191_/C vssd1 vssd1 vccd1 vccd1 _22454_/X sky130_fd_sc_hd__buf_6
X_25242_ _25709_/CLK hold442/X vssd1 vssd1 vccd1 vccd1 hold440/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21405_ _21405_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21410_/A sky130_fd_sc_hd__nand2_1
X_25173_ _25174_/CLK hold367/X vssd1 vssd1 vccd1 vccd1 hold365/A sky130_fd_sc_hd__dfxtp_1
X_22385_ _22383_/Y _22384_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _22385_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24124_ _24124_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24125_/A sky130_fd_sc_hd__and2_1
XFILLER_0_60_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21336_ _21694_/B _21385_/A vssd1 vssd1 vccd1 vccd1 _21338_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_130_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24055_ _24055_/A vssd1 vssd1 vccd1 vccd1 _26085_/D sky130_fd_sc_hd__clkbuf_1
Xhold560 hold560/A vssd1 vssd1 vccd1 vccd1 hold560/X sky130_fd_sc_hd__dlygate4sd3_1
X_21267_ _21267_/A _25875_/Q vssd1 vssd1 vccd1 vccd1 _21271_/B sky130_fd_sc_hd__nand2_1
Xhold571 hold571/A vssd1 vssd1 vccd1 vccd1 hold571/X sky130_fd_sc_hd__dlygate4sd3_1
X_23006_ _23004_/X _23005_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _23006_/Y sky130_fd_sc_hd__a21oi_1
Xhold582 hold582/A vssd1 vssd1 vccd1 vccd1 hold582/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold593 hold593/A vssd1 vssd1 vccd1 vccd1 hold593/X sky130_fd_sc_hd__dlygate4sd3_1
X_20218_ _20218_/A _20218_/B vssd1 vssd1 vccd1 vccd1 _21086_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_99_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21198_ _21198_/A _21198_/B _21198_/C vssd1 vssd1 vccd1 vccd1 _21199_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_60_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20149_ _20151_/A _20151_/B vssd1 vssd1 vccd1 vccd1 _20150_/A sky130_fd_sc_hd__nand2_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24957_ _24955_/X _24956_/X _24957_/S vssd1 vssd1 vccd1 vccd1 _24958_/A sky130_fd_sc_hd__mux2_1
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _26256_/Q _25625_/Q vssd1 vssd1 vccd1 vccd1 _14425_/A sky130_fd_sc_hd__xor2_1
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1260 _25892_/Q vssd1 vssd1 vccd1 vccd1 _23053_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ _25839_/Q _13466_/A _14709_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14711_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1271 _12945_/X vssd1 vssd1 vccd1 vccd1 _25039_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1282 _25561_/Q vssd1 vssd1 vccd1 vccd1 _16851_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_23908_ _24560_/A vssd1 vssd1 vccd1 vccd1 _24002_/B sky130_fd_sc_hd__buf_8
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15690_ _16930_/A _15690_/B vssd1 vssd1 vccd1 vccd1 _15691_/B sky130_fd_sc_hd__nand2_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1293 _12834_/X vssd1 vssd1 vccd1 vccd1 _25018_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24888_ _16081_/B _16095_/B _24942_/S vssd1 vssd1 vccd1 vccd1 _24889_/A sky130_fd_sc_hd__mux2_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _14641_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14641_/Y sky130_fd_sc_hd__nand2_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23839_ _23839_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23840_/A sky130_fd_sc_hd__and2_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17360_ _19504_/A _17360_/B vssd1 vssd1 vccd1 vccd1 _17601_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_170_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14572_ _14572_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14572_/Y sky130_fd_sc_hd__nand2_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16311_ _16490_/A _16334_/A _16310_/X vssd1 vssd1 vccd1 vccd1 _16313_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_137_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25509_ _26052_/CLK _25509_/D vssd1 vssd1 vccd1 vccd1 _25509_/Q sky130_fd_sc_hd__dfxtp_1
X_13523_ hold891/A vssd1 vssd1 vccd1 vccd1 _18186_/B sky130_fd_sc_hd__inv_2
XFILLER_0_165_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17291_ _25643_/Q vssd1 vssd1 vccd1 vccd1 _20000_/B sky130_fd_sc_hd__inv_2
XFILLER_0_138_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19030_ _19028_/Y _19029_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25701_/D sky130_fd_sc_hd__a21oi_1
X_16242_ _16473_/A hold972/X vssd1 vssd1 vccd1 vccd1 _16242_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_125_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13454_ _13220_/A _14684_/A _13242_/A _25708_/Q vssd1 vssd1 vccd1 vccd1 _13454_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16173_ _16182_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16173_/Y sky130_fd_sc_hd__nand2_1
X_13385_ _13220_/X _14648_/A _13242_/X _19744_/A vssd1 vssd1 vccd1 vccd1 _13385_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15124_ _15124_/A _15124_/B vssd1 vssd1 vccd1 vccd1 _15162_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15055_ _15055_/A _15067_/A vssd1 vssd1 vccd1 vccd1 _15055_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19932_ _19930_/Y _19931_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _19932_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14006_ hold555/X _14005_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold556/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19863_ _19861_/X _19862_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19863_/Y sky130_fd_sc_hd__a21oi_1
X_18814_ _18814_/A _18814_/B _18814_/C vssd1 vssd1 vccd1 vccd1 _22541_/A sky130_fd_sc_hd__nand3_2
X_19794_ _19792_/X _19793_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19794_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18745_ _22463_/B _25635_/Q vssd1 vssd1 vccd1 vccd1 _18747_/A sky130_fd_sc_hd__nand2_1
X_15957_ _15955_/X _15956_/Y _15805_/X vssd1 vssd1 vccd1 vccd1 hold881/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_163_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14908_ _14909_/B _14909_/A vssd1 vssd1 vccd1 vccd1 _14910_/A sky130_fd_sc_hd__or2_1
XFILLER_0_76_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18676_ _18676_/A _20400_/A vssd1 vssd1 vccd1 vccd1 _18981_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_37_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15888_ hold653/X vssd1 vssd1 vccd1 vccd1 _15891_/B sky130_fd_sc_hd__inv_2
XFILLER_0_114_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17627_ _18252_/A _17627_/B vssd1 vssd1 vccd1 vccd1 _17627_/Y sky130_fd_sc_hd__nand2_1
X_14839_ _14839_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14839_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17558_ _17556_/X _17528_/X _17557_/X vssd1 vssd1 vccd1 vccd1 _17559_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_175_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16509_ _16676_/A _15568_/A _16508_/Y vssd1 vssd1 vccd1 vccd1 _16511_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_46_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17489_ _17605_/A _17489_/B vssd1 vssd1 vccd1 vccd1 _17489_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19228_ _19452_/A hold937/X vssd1 vssd1 vccd1 vccd1 hold938/A sky130_fd_sc_hd__nand2_1
XFILLER_0_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19159_ _19159_/A _21889_/A vssd1 vssd1 vccd1 vccd1 _20174_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22170_ _22147_/X _22169_/Y _21791_/X vssd1 vssd1 vccd1 vccd1 _22170_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_124_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21121_ _26308_/Q hold620/X vssd1 vssd1 vccd1 vccd1 _21121_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_140_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21052_ _21054_/B _21054_/C vssd1 vssd1 vccd1 vccd1 _21053_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20003_ _20003_/A _22670_/B vssd1 vssd1 vccd1 vccd1 _20007_/B sky130_fd_sc_hd__nand2_1
X_25860_ _25860_/CLK _25860_/D vssd1 vssd1 vccd1 vccd1 _25860_/Q sky130_fd_sc_hd__dfxtp_4
X_24811_ hold2693/X hold2684/X _24817_/S vssd1 vssd1 vccd1 vccd1 _24812_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25791_ _25791_/CLK _25791_/D vssd1 vssd1 vccd1 vccd1 _25791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24742_ _24742_/A vssd1 vssd1 vccd1 vccd1 _26309_/D sky130_fd_sc_hd__clkbuf_1
X_21954_ _23151_/A _22703_/A vssd1 vssd1 vccd1 vccd1 _21962_/A sky130_fd_sc_hd__nand2_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20905_ _20905_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _20905_/Y sky130_fd_sc_hd__nand2_1
X_21885_ _23119_/A _22651_/A vssd1 vssd1 vccd1 vccd1 _21893_/A sky130_fd_sc_hd__nand2_1
X_24673_ _24673_/A vssd1 vssd1 vccd1 vccd1 _26286_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23624_ _23624_/A vssd1 vssd1 vccd1 vccd1 _25947_/D sky130_fd_sc_hd__clkbuf_1
X_20836_ _20835_/B _20836_/B _20836_/C vssd1 vssd1 vccd1 vccd1 _20837_/B sky130_fd_sc_hd__nand3b_4
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20767_ _20767_/A _21351_/C _20767_/C vssd1 vssd1 vccd1 vccd1 _20768_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23555_ _23543_/X _23554_/X _24949_/S vssd1 vssd1 vccd1 vccd1 _23555_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22506_ _22506_/A _23001_/B _22506_/C vssd1 vssd1 vccd1 vccd1 _22506_/X sky130_fd_sc_hd__and3_1
XFILLER_0_92_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23486_ _24940_/S hold296/A _23485_/X vssd1 vssd1 vccd1 vccd1 _23486_/Y sky130_fd_sc_hd__o21ai_1
X_26274_ _26279_/CLK _26274_/D vssd1 vssd1 vccd1 vccd1 _26274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20698_ _22586_/A vssd1 vssd1 vccd1 vccd1 _21235_/A sky130_fd_sc_hd__buf_6
XFILLER_0_135_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22437_ _18736_/A _25826_/Q _22435_/Y _22436_/Y vssd1 vssd1 vccd1 vccd1 _22438_/B
+ sky130_fd_sc_hd__a31o_1
X_25225_ _25678_/CLK hold622/X vssd1 vssd1 vccd1 vccd1 hold620/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13170_ _13170_/A vssd1 vssd1 vccd1 vccd1 _19257_/A sky130_fd_sc_hd__buf_4
X_22368_ _22368_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _22368_/X sky130_fd_sc_hd__and2_1
XFILLER_0_27_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25156_ _25738_/CLK hold842/X vssd1 vssd1 vccd1 vccd1 hold841/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24107_ _24107_/A vssd1 vssd1 vccd1 vccd1 _26102_/D sky130_fd_sc_hd__clkbuf_1
X_21319_ _21319_/A _21319_/B _21319_/C vssd1 vssd1 vccd1 vccd1 _21323_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25087_ _26299_/CLK _25087_/D vssd1 vssd1 vccd1 vccd1 _25087_/Q sky130_fd_sc_hd__dfxtp_1
X_22299_ _22299_/A _22299_/B vssd1 vssd1 vccd1 vccd1 _22299_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_103_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24038_ hold2286/X _26081_/Q _24047_/S vssd1 vssd1 vccd1 vccd1 _24038_/X sky130_fd_sc_hd__mux2_1
Xhold390 hold390/A vssd1 vssd1 vccd1 vccd1 hold390/X sky130_fd_sc_hd__dlygate4sd3_1
X_16860_ _16935_/A _16865_/B vssd1 vssd1 vccd1 vccd1 _16862_/B sky130_fd_sc_hd__nand2_1
X_15811_ _23191_/B _15811_/B vssd1 vssd1 vccd1 vccd1 _23188_/B sky130_fd_sc_hd__xor2_1
X_16791_ _17568_/A vssd1 vssd1 vccd1 vccd1 _16791_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_189_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25989_ _25991_/CLK _25989_/D vssd1 vssd1 vccd1 vccd1 _25989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18530_ _18530_/A _18530_/B _18530_/C vssd1 vssd1 vccd1 vccd1 _22181_/A sky130_fd_sc_hd__nand3_2
X_15742_ _15743_/A _15744_/A vssd1 vssd1 vccd1 vccd1 _15746_/A sky130_fd_sc_hd__nor2_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _17479_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12954_/X sky130_fd_sc_hd__or2_1
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1090 _19611_/Y vssd1 vssd1 vccd1 vccd1 _25744_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _22095_/B _25621_/Q vssd1 vssd1 vccd1 vccd1 _18463_/A sky130_fd_sc_hd__nand2_1
X_15673_ _16923_/A _15673_/B vssd1 vssd1 vccd1 vccd1 _15674_/B sky130_fd_sc_hd__and2_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _12840_/X _12883_/X _12827_/X _12884_/X vssd1 vssd1 vccd1 vccd1 _12885_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_193_clk _26093_/CLK vssd1 vssd1 vccd1 vccd1 _25619_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17412_ _17586_/A _17637_/B vssd1 vssd1 vccd1 vccd1 _17413_/B sky130_fd_sc_hd__xnor2_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _14645_/A hold470/X vssd1 vssd1 vccd1 vccd1 hold471/A sky130_fd_sc_hd__nand2_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18392_ _18392_/A _18392_/B vssd1 vssd1 vccd1 vccd1 _18392_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _17393_/A _17343_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17343_/X sky130_fd_sc_hd__and3_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14555_ _14585_/A hold374/X vssd1 vssd1 vccd1 vccd1 hold375/A sky130_fd_sc_hd__nand2_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13506_ _18070_/B _13518_/B vssd1 vssd1 vccd1 vccd1 _13506_/Y sky130_fd_sc_hd__nor2_1
X_17274_ _25608_/Q vssd1 vssd1 vccd1 vccd1 _20965_/B sky130_fd_sc_hd__inv_2
XFILLER_0_183_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14486_ _14525_/A hold311/X vssd1 vssd1 vccd1 vccd1 hold312/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19013_ _19011_/X _18879_/X _19012_/X vssd1 vssd1 vccd1 vccd1 _19014_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_183_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16225_ _16238_/B _16225_/B vssd1 vssd1 vccd1 vccd1 _16228_/B sky130_fd_sc_hd__and2_1
XFILLER_0_180_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13437_ _13522_/A _13435_/X _23629_/B _13436_/X vssd1 vssd1 vccd1 vccd1 _13437_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16156_ _16156_/A _16156_/B vssd1 vssd1 vccd1 vccd1 _16161_/B sky130_fd_sc_hd__nor2_1
X_13368_ _26196_/Q _13239_/X _13367_/X vssd1 vssd1 vccd1 vccd1 _13368_/X sky130_fd_sc_hd__a21o_1
X_15107_ _15107_/A _15085_/Y vssd1 vssd1 vccd1 vccd1 _15110_/B sky130_fd_sc_hd__nor2b_1
XFILLER_0_122_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16087_ _16088_/B _16088_/A vssd1 vssd1 vccd1 vccd1 _16089_/A sky130_fd_sc_hd__or2_1
X_13299_ _24745_/A vssd1 vssd1 vccd1 vccd1 _24560_/A sky130_fd_sc_hd__buf_12
X_15038_ _15051_/A _15270_/A vssd1 vssd1 vccd1 vccd1 _15038_/X sky130_fd_sc_hd__or2_1
X_19915_ _19913_/X _19914_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19915_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2708 _26255_/Q vssd1 vssd1 vccd1 vccd1 hold2708/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2719 _26265_/Q vssd1 vssd1 vccd1 vccd1 hold2719/X sky130_fd_sc_hd__dlygate4sd3_1
X_19846_ _20711_/A _19844_/Y _20716_/C vssd1 vssd1 vccd1 vccd1 _19928_/B sky130_fd_sc_hd__o21a_2
X_16989_ _25623_/Q vssd1 vssd1 vccd1 vccd1 _20099_/B sky130_fd_sc_hd__inv_2
X_19777_ _19793_/B _19862_/B vssd1 vssd1 vccd1 vccd1 _19779_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18728_ _25890_/Q _22435_/A vssd1 vssd1 vccd1 vccd1 _18736_/A sky130_fd_sc_hd__or2_2
XFILLER_0_189_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18659_ _18657_/X _18269_/X _18658_/X vssd1 vssd1 vccd1 vccd1 _18660_/A sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_184_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _25738_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21670_ _21670_/A _22902_/B vssd1 vssd1 vccd1 vccd1 _21670_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20621_ _20621_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _20621_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23340_ _23340_/A vssd1 vssd1 vccd1 vccd1 _25930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20552_ _20554_/B _20554_/C vssd1 vssd1 vccd1 vccd1 _20553_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23271_ _23271_/A vssd1 vssd1 vccd1 vccd1 _25916_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20483_ _20483_/A _22413_/B _20483_/C vssd1 vssd1 vccd1 vccd1 _20487_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_144_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22222_ _19244_/A _22221_/A _22221_/Y vssd1 vssd1 vccd1 vccd1 _22224_/A sky130_fd_sc_hd__o21ai_1
X_25010_ _26221_/CLK hold3/X vssd1 vssd1 vccd1 vccd1 _25010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22153_ _22838_/B _22154_/A vssd1 vssd1 vccd1 vccd1 _22155_/A sky130_fd_sc_hd__or2_1
XFILLER_0_112_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21104_ _21104_/A _25869_/Q vssd1 vssd1 vccd1 vccd1 _21109_/A sky130_fd_sc_hd__nand2_1
X_22084_ _22084_/A _23058_/A _22084_/C vssd1 vssd1 vccd1 vccd1 _22084_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25912_ _25913_/CLK _25912_/D vssd1 vssd1 vccd1 vccd1 _25912_/Q sky130_fd_sc_hd__dfxtp_4
X_21035_ _21548_/B _21497_/C vssd1 vssd1 vccd1 vccd1 _21036_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25843_ _26208_/CLK _25843_/D vssd1 vssd1 vccd1 vccd1 _25843_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_22_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25774_ _26251_/CLK _25774_/D vssd1 vssd1 vccd1 vccd1 _25774_/Q sky130_fd_sc_hd__dfxtp_1
X_22986_ _22986_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _22986_/Y sky130_fd_sc_hd__nand2_1
X_24725_ hold2103/X _26304_/Q _24740_/S vssd1 vssd1 vccd1 vccd1 _24725_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_175_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _26236_/CLK sky130_fd_sc_hd__clkbuf_16
X_21937_ _21937_/A _25863_/Q vssd1 vssd1 vccd1 vccd1 _21937_/Y sky130_fd_sc_hd__nand2_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12674_/B _12674_/A vssd1 vssd1 vccd1 vccd1 _12670_/Y sky130_fd_sc_hd__nand2_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24656_ _24656_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24657_/A sky130_fd_sc_hd__and2_1
XFILLER_0_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21868_ _21868_/A _25861_/Q vssd1 vssd1 vccd1 vccd1 _21868_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_167_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23607_ hold2283/X hold2258/X _23677_/S vssd1 vssd1 vccd1 vccd1 _23608_/A sky130_fd_sc_hd__mux2_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20819_ _20822_/A _20822_/C vssd1 vssd1 vccd1 vccd1 _20820_/A sky130_fd_sc_hd__nand2_1
X_21799_ _21799_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _21799_/X sky130_fd_sc_hd__and2_1
X_24587_ hold2575/X _26259_/Q _24587_/S vssd1 vssd1 vccd1 vccd1 _24587_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_182_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26326_ _26330_/CLK _26326_/D vssd1 vssd1 vccd1 vccd1 _26326_/Q sky130_fd_sc_hd__dfxtp_2
X_14340_ _14340_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14340_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_80_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23538_ hold23/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23538_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_93_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14271_ _14270_/Y _14277_/C _14277_/B vssd1 vssd1 vccd1 vccd1 _14271_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26257_ _26264_/CLK _26257_/D vssd1 vssd1 vccd1 vccd1 _26257_/Q sky130_fd_sc_hd__dfxtp_4
X_23469_ _23463_/X _23468_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _23469_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_123_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16010_ _16018_/B vssd1 vssd1 vccd1 vccd1 _16011_/A sky130_fd_sc_hd__inv_2
XFILLER_0_122_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25208_ _25793_/CLK hold779/X vssd1 vssd1 vccd1 vccd1 hold777/A sky130_fd_sc_hd__dfxtp_1
X_13222_ _26301_/Q _19373_/A vssd1 vssd1 vccd1 vccd1 _14566_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_104_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26188_ _26190_/CLK _26188_/D vssd1 vssd1 vccd1 vccd1 _26188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13153_ _26290_/Q _19216_/A vssd1 vssd1 vccd1 vccd1 _14533_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_0_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25139_ _25785_/CLK hold535/X vssd1 vssd1 vccd1 vccd1 hold533/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17961_ _19059_/A _18434_/A vssd1 vssd1 vccd1 vccd1 _17962_/B sky130_fd_sc_hd__xnor2_4
X_13084_ _13049_/X _14491_/A _13067_/X _21749_/A vssd1 vssd1 vccd1 vccd1 _13084_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16912_ _16910_/X _16711_/X _16911_/Y _25891_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16913_/A sky130_fd_sc_hd__a32o_1
X_19700_ _19697_/Y _19700_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19700_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_109_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17892_ _18612_/A _25722_/Q _18955_/C vssd1 vssd1 vccd1 vccd1 _17893_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_40_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16843_ _16424_/B _16842_/Y _15621_/A vssd1 vssd1 vccd1 vccd1 _16843_/Y sky130_fd_sc_hd__a21oi_1
X_19631_ _20131_/A _22179_/B _25624_/Q vssd1 vssd1 vccd1 vccd1 _20135_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_189_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19562_ _21264_/A _19560_/Y _21268_/C vssd1 vssd1 vccd1 vccd1 _19649_/B sky130_fd_sc_hd__o21a_2
X_16774_ _16976_/B _16774_/B vssd1 vssd1 vccd1 vccd1 _16774_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_88_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13986_ hold719/X _13985_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold720/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_177_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18513_ _18718_/A _18858_/A vssd1 vssd1 vccd1 vccd1 _18514_/B sky130_fd_sc_hd__xnor2_1
X_15725_ _23108_/B _15812_/B vssd1 vssd1 vccd1 vccd1 _16625_/B sky130_fd_sc_hd__nand2_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12937_ _12891_/X _14400_/A _12909_/X _25618_/Q vssd1 vssd1 vccd1 vccd1 _12937_/X
+ sky130_fd_sc_hd__a22o_1
X_19493_ _19493_/A _19493_/B vssd1 vssd1 vccd1 vccd1 _19493_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_87_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_166_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _26289_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18444_ _25876_/Q _22064_/A vssd1 vssd1 vccd1 vccd1 _18452_/A sky130_fd_sc_hd__or2_2
X_15656_ _15656_/A _15656_/B vssd1 vssd1 vccd1 vccd1 _15657_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _26108_/Q _12748_/X _12867_/X vssd1 vssd1 vccd1 vccd1 _12868_/X sky130_fd_sc_hd__a21o_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _14605_/Y hold294/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold295/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18375_ _18375_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18375_/Y sky130_fd_sc_hd__nand2_1
X_15587_ hold908/X vssd1 vssd1 vccd1 vccd1 _15589_/A sky130_fd_sc_hd__inv_2
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _12726_/B _14319_/A _12752_/X _25592_/Q vssd1 vssd1 vccd1 vccd1 _12799_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17326_ _17324_/Y _17325_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _17326_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_141_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14538_ _14536_/Y hold270/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold271/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17257_ _17255_/X _17241_/X _17256_/X vssd1 vssd1 vccd1 vccd1 _17258_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_126_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14469_ _14469_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14469_/Y sky130_fd_sc_hd__nand2_1
X_16208_ _16208_/A _16208_/B vssd1 vssd1 vccd1 vccd1 _16210_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_183_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17188_ _17186_/X _23187_/B _17187_/X vssd1 vssd1 vccd1 vccd1 _17189_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16139_ _16139_/A _16139_/B vssd1 vssd1 vccd1 vccd1 _16140_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2505 _23971_/X vssd1 vssd1 vccd1 vccd1 _23972_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2516 _24980_/Q vssd1 vssd1 vccd1 vccd1 _12632_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2527 _15182_/Y vssd1 vssd1 vccd1 vccd1 hold2527/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2538 _12667_/X vssd1 vssd1 vccd1 vccd1 _12668_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1804 _25591_/Q vssd1 vssd1 vccd1 vccd1 _17151_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2549 _24989_/Q vssd1 vssd1 vccd1 vccd1 _12686_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1815 _25842_/Q vssd1 vssd1 vccd1 vccd1 _21896_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1826 _22321_/Y vssd1 vssd1 vccd1 vccd1 _25856_/D sky130_fd_sc_hd__dlygate4sd3_1
X_19829_ _19826_/Y _19829_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19829_/X sky130_fd_sc_hd__and3b_1
Xhold1837 _25848_/Q vssd1 vssd1 vccd1 vccd1 _22088_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1848 _23581_/Y vssd1 vssd1 vccd1 vccd1 hold1848/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1859 _22342_/Y vssd1 vssd1 vccd1 vccd1 _25857_/D sky130_fd_sc_hd__dlygate4sd3_1
X_22840_ _23151_/B _22840_/B vssd1 vssd1 vccd1 vccd1 _22842_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22771_ _22762_/Y _22770_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22771_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_17_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_157_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _25797_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_189_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24510_ hold2729/X hold2683/X _24510_/S vssd1 vssd1 vccd1 vccd1 _24511_/A sky130_fd_sc_hd__mux2_1
X_21722_ _21722_/A _22145_/B vssd1 vssd1 vccd1 vccd1 _21722_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_38_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25490_ _25933_/CLK hold664/X vssd1 vssd1 vccd1 vccd1 hold662/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24441_ _24441_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24442_/A sky130_fd_sc_hd__and2_1
X_21653_ _21653_/A _21653_/B vssd1 vssd1 vccd1 vccd1 _21654_/A sky130_fd_sc_hd__nand2_1
X_20604_ _20604_/A _20604_/B vssd1 vssd1 vccd1 vccd1 _20606_/A sky130_fd_sc_hd__nand2_1
X_21584_ _26332_/Q hold751/X vssd1 vssd1 vccd1 vccd1 _21584_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24372_ hold2409/X hold2325/X _24433_/S vssd1 vssd1 vccd1 vccd1 _24373_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_90_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26111_ _26112_/CLK _26111_/D vssd1 vssd1 vccd1 vccd1 _26111_/Q sky130_fd_sc_hd__dfxtp_1
X_23323_ _23324_/B _23324_/A vssd1 vssd1 vccd1 vccd1 _23323_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20535_ _20535_/A _20535_/B vssd1 vssd1 vccd1 vccd1 _20536_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26042_ _26042_/CLK _26042_/D vssd1 vssd1 vccd1 vccd1 _26042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23254_ _23254_/A _25912_/Q vssd1 vssd1 vccd1 vccd1 _23255_/A sky130_fd_sc_hd__nand2_1
X_20466_ _20463_/Y _20464_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _20466_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_162_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22205_ _22203_/X _15839_/B _22204_/Y hold955/X _21725_/X vssd1 vssd1 vccd1 vccd1
+ _22206_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_132_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23185_ _23185_/A _23185_/B vssd1 vssd1 vccd1 vccd1 _23186_/B sky130_fd_sc_hd__nand2_1
X_20397_ _20396_/B _20397_/B _20397_/C vssd1 vssd1 vccd1 vccd1 _20398_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_24_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22136_ _22136_/A _22136_/B vssd1 vssd1 vccd1 vccd1 _22137_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_100_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22067_ _22067_/A _22067_/B vssd1 vssd1 vccd1 vccd1 _22067_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21018_ _21018_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _21018_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25826_ _25865_/CLK _25826_/D vssd1 vssd1 vccd1 vccd1 _25826_/Q sky130_fd_sc_hd__dfxtp_2
X_13840_ _18873_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13840_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_96_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_148_clk clkbuf_4_11__f_clk/X vssd1 vssd1 vccd1 vccd1 _26184_/CLK sky130_fd_sc_hd__clkbuf_16
X_13771_ _26261_/Q _13612_/X _13605_/X _13770_/Y vssd1 vssd1 vccd1 vccd1 _13772_/B
+ sky130_fd_sc_hd__a22o_1
X_25757_ _25773_/CLK _25757_/D vssd1 vssd1 vccd1 vccd1 _25757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22969_ _22969_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _22969_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15510_ _22911_/B _16369_/B vssd1 vssd1 vccd1 vccd1 _16464_/B sky130_fd_sc_hd__nand2_1
X_24708_ _24708_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24709_/A sky130_fd_sc_hd__and2_1
XFILLER_0_85_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12722_ _25582_/Q vssd1 vssd1 vccd1 vccd1 _20023_/B sky130_fd_sc_hd__inv_2
XFILLER_0_97_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16490_ _16490_/A _16490_/B vssd1 vssd1 vccd1 vccd1 _16495_/A sky130_fd_sc_hd__nand2_1
X_25688_ _26317_/CLK _25688_/D vssd1 vssd1 vccd1 vccd1 _25688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15441_ _15441_/A _15441_/B vssd1 vssd1 vccd1 vccd1 _15442_/B sky130_fd_sc_hd__nor2_1
X_12653_ _12653_/A vssd1 vssd1 vccd1 vccd1 _24982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24639_ hold2663/X hold2632/X _24664_/S vssd1 vssd1 vccd1 vccd1 _24640_/A sky130_fd_sc_hd__mux2_1
X_18160_ _18160_/A _20317_/A vssd1 vssd1 vccd1 vccd1 _20309_/A sky130_fd_sc_hd__nand2_4
X_15372_ _15372_/A vssd1 vssd1 vccd1 vccd1 _15374_/A sky130_fd_sc_hd__inv_2
XFILLER_0_68_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12584_ _12584_/A vssd1 vssd1 vccd1 vccd1 _24969_/D sky130_fd_sc_hd__inv_2
XFILLER_0_81_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17111_ _17111_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17111_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14323_ _14344_/A hold281/X vssd1 vssd1 vccd1 vccd1 hold282/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26309_ _26313_/CLK _26309_/D vssd1 vssd1 vccd1 vccd1 _26309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18091_ _21869_/B _25605_/Q vssd1 vssd1 vccd1 vccd1 _18093_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_180_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17042_ _19644_/A _17042_/B vssd1 vssd1 vccd1 vccd1 _17505_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_162_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14254_ _14260_/A hold431/X vssd1 vssd1 vccd1 vccd1 hold432/A sky130_fd_sc_hd__nand2_1
XFILLER_0_52_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13205_ _18455_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13205_/X sky130_fd_sc_hd__or2_1
X_14185_ _26327_/Q _13518_/B _14170_/X _14184_/Y vssd1 vssd1 vccd1 vccd1 _14186_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13136_ _13049_/X _14521_/A _13067_/X _25656_/Q vssd1 vssd1 vccd1 vccd1 _13136_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ _19199_/A vssd1 vssd1 vccd1 vccd1 _19186_/A sky130_fd_sc_hd__buf_8
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17944_ _18529_/A _17944_/B _18083_/C vssd1 vssd1 vccd1 vccd1 _17945_/C sky130_fd_sc_hd__nand3_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _13242_/A vssd1 vssd1 vccd1 vccd1 _13067_/X sky130_fd_sc_hd__buf_12
XFILLER_0_40_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17875_ _17875_/A _17875_/B vssd1 vssd1 vccd1 vccd1 _17877_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_174_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19614_ _19613_/Y _19272_/X _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19615_/B
+ sky130_fd_sc_hd__a211o_1
X_16826_ _16826_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16826_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16757_ _16858_/A _16757_/B vssd1 vssd1 vccd1 vccd1 _16757_/Y sky130_fd_sc_hd__nand2_1
X_19545_ _19542_/Y _19545_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19545_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_177_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13969_ _25790_/Q vssd1 vssd1 vccd1 vccd1 _18087_/B sky130_fd_sc_hd__inv_2
XFILLER_0_49_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_139_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _25808_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15708_ _23092_/B _15776_/B vssd1 vssd1 vccd1 vccd1 _15709_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16688_ _16686_/Y hold609/X _16594_/X vssd1 vssd1 vccd1 vccd1 hold610/A sky130_fd_sc_hd__a21oi_1
X_19476_ _19493_/B _19565_/B vssd1 vssd1 vccd1 vccd1 _19478_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15639_ _15640_/B _16911_/A vssd1 vssd1 vccd1 vccd1 _15641_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_75_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18427_ _18427_/A _25811_/Q _18427_/C vssd1 vssd1 vccd1 vccd1 _21270_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_189_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18358_ _19518_/A vssd1 vssd1 vccd1 vccd1 _21947_/B sky130_fd_sc_hd__inv_2
XFILLER_0_17_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17309_ _17393_/A _17309_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17309_/X sky130_fd_sc_hd__and3_1
XFILLER_0_173_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18289_ _21080_/B _21812_/A vssd1 vssd1 vccd1 vccd1 _21074_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20320_ _21169_/C vssd1 vssd1 vccd1 vccd1 _21172_/B sky130_fd_sc_hd__inv_2
XFILLER_0_4_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold901 hold901/A vssd1 vssd1 vccd1 vccd1 hold901/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 hold912/A vssd1 vssd1 vccd1 vccd1 hold912/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 hold923/A vssd1 vssd1 vccd1 vccd1 hold923/X sky130_fd_sc_hd__dlygate4sd3_1
X_20251_ _20251_/A _20251_/B _20251_/C vssd1 vssd1 vccd1 vccd1 _20254_/C sky130_fd_sc_hd__nand3_1
Xhold934 hold934/A vssd1 vssd1 vccd1 vccd1 hold934/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 hold945/A vssd1 vssd1 vccd1 vccd1 hold945/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold956 hold956/A vssd1 vssd1 vccd1 vccd1 hold956/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 hold967/A vssd1 vssd1 vccd1 vccd1 hold967/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold978 hold978/A vssd1 vssd1 vccd1 vccd1 hold978/X sky130_fd_sc_hd__dlygate4sd3_1
X_20182_ _21059_/C vssd1 vssd1 vccd1 vccd1 _21062_/B sky130_fd_sc_hd__inv_2
Xhold989 hold989/A vssd1 vssd1 vccd1 vccd1 hold989/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2302 _26122_/Q vssd1 vssd1 vccd1 vccd1 hold2302/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24990_ _24990_/CLK _24990_/D vssd1 vssd1 vccd1 vccd1 _24990_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2313 _24231_/X vssd1 vssd1 vccd1 vccd1 _24232_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2324 _26119_/Q vssd1 vssd1 vccd1 vccd1 hold2324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2335 _26145_/Q vssd1 vssd1 vccd1 vccd1 hold2335/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2346 _25994_/Q vssd1 vssd1 vccd1 vccd1 hold2346/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1601 _23166_/Y vssd1 vssd1 vccd1 vccd1 _25899_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23941_ hold2471/X hold2469/X _24001_/S vssd1 vssd1 vccd1 vccd1 _23942_/A sky130_fd_sc_hd__mux2_1
Xhold2357 _26057_/Q vssd1 vssd1 vccd1 vccd1 hold2357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1612 _25832_/Q vssd1 vssd1 vccd1 vccd1 _21639_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1623 _25649_/Q vssd1 vssd1 vccd1 vccd1 _17966_/B sky130_fd_sc_hd__clkbuf_2
Xhold2368 _26052_/Q vssd1 vssd1 vccd1 vccd1 hold2368/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2379 _25664_/Q vssd1 vssd1 vccd1 vccd1 _13182_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1634 _25644_/Q vssd1 vssd1 vccd1 vccd1 _17649_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1645 _25614_/Q vssd1 vssd1 vccd1 vccd1 _17427_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1656 _22806_/Y vssd1 vssd1 vccd1 vccd1 _25877_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23872_ _23872_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23873_/A sky130_fd_sc_hd__and2_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1667 _25807_/Q vssd1 vssd1 vccd1 vccd1 _21181_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1678 _25608_/Q vssd1 vssd1 vccd1 vccd1 _17366_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1689 _17260_/Y vssd1 vssd1 vccd1 vccd1 _25599_/D sky130_fd_sc_hd__dlygate4sd3_1
X_25611_ _26117_/CLK _25611_/D vssd1 vssd1 vccd1 vccd1 _25611_/Q sky130_fd_sc_hd__dfxtp_4
X_22823_ _23135_/B _22823_/B vssd1 vssd1 vccd1 vccd1 _22825_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25542_ _26047_/CLK _25542_/D vssd1 vssd1 vccd1 vccd1 _25542_/Q sky130_fd_sc_hd__dfxtp_1
X_22754_ _22754_/A _22900_/B vssd1 vssd1 vccd1 vccd1 _22754_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_177_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21705_ _21708_/B _21709_/A vssd1 vssd1 vccd1 vccd1 _21707_/A sky130_fd_sc_hd__nand2_1
X_25473_ _26064_/CLK _25473_/D vssd1 vssd1 vccd1 vccd1 _25473_/Q sky130_fd_sc_hd__dfxtp_1
X_22685_ _22685_/A _23001_/B _22685_/C vssd1 vssd1 vccd1 vccd1 _22685_/X sky130_fd_sc_hd__and3_1
XFILLER_0_137_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24424_ hold2214/X _26206_/Q _24433_/S vssd1 vssd1 vccd1 vccd1 _24424_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_165_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21636_ _21636_/A _21636_/B _21635_/X vssd1 vssd1 vccd1 vccd1 _21637_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24355_ _24355_/A vssd1 vssd1 vccd1 vccd1 _26183_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21567_ _26331_/Q _19130_/X hold473/X vssd1 vssd1 vccd1 vccd1 _21570_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23306_ _23306_/A hold985/X _25922_/Q vssd1 vssd1 vccd1 vccd1 _23307_/B sky130_fd_sc_hd__and3_1
XFILLER_0_50_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20518_ _20518_/A _20518_/B vssd1 vssd1 vccd1 vccd1 _20522_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24286_ _24286_/A vssd1 vssd1 vccd1 vccd1 _26160_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21498_ _21498_/A _21546_/A vssd1 vssd1 vccd1 vccd1 _21500_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_127_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26025_ _26042_/CLK _26025_/D vssd1 vssd1 vccd1 vccd1 _26025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23237_ _24949_/S _23238_/A vssd1 vssd1 vccd1 vccd1 _23237_/X sky130_fd_sc_hd__or2_1
X_20449_ _21252_/B _21547_/A vssd1 vssd1 vccd1 vccd1 _20452_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_120_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23168_ _23168_/A _23168_/B vssd1 vssd1 vccd1 vccd1 _23169_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22119_ _22119_/A _25878_/Q vssd1 vssd1 vccd1 vccd1 _22119_/Y sky130_fd_sc_hd__nand2_1
X_15990_ _15988_/X _15989_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _15990_/X sky130_fd_sc_hd__a21o_1
X_23099_ _23099_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _23099_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_98_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14941_ _14947_/B _14942_/A vssd1 vssd1 vccd1 vccd1 _14941_/X sky130_fd_sc_hd__or2_1
X_17660_ _19089_/B _25582_/Q vssd1 vssd1 vccd1 vccd1 _17662_/B sky130_fd_sc_hd__nand2_1
X_14872_ _14872_/A _14899_/B vssd1 vssd1 vccd1 vccd1 _14872_/Y sky130_fd_sc_hd__nand2_1
X_16611_ _16620_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16611_/Y sky130_fd_sc_hd__nand2_1
X_25809_ _25812_/CLK _25809_/D vssd1 vssd1 vccd1 vccd1 _25809_/Q sky130_fd_sc_hd__dfxtp_2
X_13823_ _13823_/A _13823_/B vssd1 vssd1 vccd1 vccd1 _13823_/Y sky130_fd_sc_hd__nand2_1
X_17591_ _17605_/A _17591_/B vssd1 vssd1 vccd1 vccd1 _17591_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16542_ _16542_/A vssd1 vssd1 vccd1 vccd1 _16543_/A sky130_fd_sc_hd__inv_2
X_19330_ _19327_/Y _19330_/B _19980_/B vssd1 vssd1 vccd1 vccd1 _19330_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13754_ _13760_/A hold500/X vssd1 vssd1 vccd1 vccd1 hold501/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12705_ _12707_/B _23377_/B vssd1 vssd1 vccd1 vccd1 _12705_/X sky130_fd_sc_hd__and2_1
X_19261_ _19261_/A _19261_/B vssd1 vssd1 vccd1 vccd1 _19261_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16473_ _16473_/A hold970/X vssd1 vssd1 vccd1 vccd1 _16473_/Y sky130_fd_sc_hd__nand2_1
X_13685_ _13703_/A _13685_/B vssd1 vssd1 vccd1 vccd1 _13685_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_155_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18212_ _18252_/A _18212_/B vssd1 vssd1 vccd1 vccd1 _18212_/Y sky130_fd_sc_hd__nand2_1
X_15424_ _15425_/B _16831_/A vssd1 vssd1 vccd1 vccd1 _15426_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_66_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12636_ _12636_/A _24836_/B _12636_/C vssd1 vssd1 vccd1 vccd1 _12636_/X sky130_fd_sc_hd__and3_1
X_19192_ _26218_/Q hold530/X vssd1 vssd1 vccd1 vccd1 _19192_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_182_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18143_ _19067_/A _18143_/B vssd1 vssd1 vccd1 vccd1 _18143_/X sky130_fd_sc_hd__xor2_2
X_15355_ _15356_/B _16803_/A vssd1 vssd1 vccd1 vccd1 _15357_/A sky130_fd_sc_hd__nor2_1
X_12567_ _12567_/A vssd1 vssd1 vccd1 vccd1 _23598_/A sky130_fd_sc_hd__inv_2
XFILLER_0_136_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14306_ _14304_/Y hold12/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_170_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18074_ _18074_/A _25780_/Q _18074_/C vssd1 vssd1 vccd1 vccd1 _20252_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_81_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15286_ _22679_/B _15812_/B vssd1 vssd1 vccd1 vccd1 _15287_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_145_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12498_ _14270_/B _24836_/B _23001_/B _12726_/B _12497_/Y vssd1 vssd1 vccd1 vccd1
+ _12498_/X sky130_fd_sc_hd__a32o_1
Xhold208 hold208/A vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 hold219/A vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__dlygate4sd3_1
X_17025_ _20132_/B _25880_/Q _25816_/Q vssd1 vssd1 vccd1 vccd1 _17026_/B sky130_fd_sc_hd__mux2_2
X_14237_ _25833_/Q vssd1 vssd1 vccd1 vccd1 _18874_/B sky130_fd_sc_hd__inv_2
XFILLER_0_145_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14168_ _14163_/Y _14167_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold840/A sky130_fd_sc_hd__a21oi_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _13109_/X _13117_/X _13096_/X _13118_/X vssd1 vssd1 vccd1 vccd1 _13119_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18976_ _19026_/A _18976_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18976_/X sky130_fd_sc_hd__and3_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ hold540/X _14098_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold541/A sky130_fd_sc_hd__a21oi_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _17927_/A _17927_/B vssd1 vssd1 vccd1 vccd1 _17928_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_56_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17858_ _18612_/A _17858_/B _18083_/C vssd1 vssd1 vccd1 vccd1 _17859_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_79_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16809_ _16810_/B _16810_/A vssd1 vssd1 vccd1 vccd1 _16809_/X sky130_fd_sc_hd__or2_1
XFILLER_0_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17789_ _18122_/C _17789_/B vssd1 vssd1 vccd1 vccd1 _18100_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_178_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19528_ _26242_/Q _19483_/X hold416/X vssd1 vssd1 vccd1 vccd1 _19528_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19459_ _21074_/A _21810_/B _25612_/Q vssd1 vssd1 vccd1 vccd1 _21078_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_147_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22470_ _23024_/B vssd1 vssd1 vccd1 vccd1 _23023_/A sky130_fd_sc_hd__inv_2
XFILLER_0_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21421_ _21421_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21426_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24140_ _24140_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24141_/A sky130_fd_sc_hd__and2_1
XFILLER_0_32_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21352_ _21710_/B _21401_/A vssd1 vssd1 vccd1 vccd1 _21354_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20303_ _20302_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20303_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_102_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24071_ hold992/X hold2164/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24072_/A sky130_fd_sc_hd__mux2_1
X_21283_ _26314_/Q hold794/X vssd1 vssd1 vccd1 vccd1 _21283_/Y sky130_fd_sc_hd__nand2_1
Xhold720 hold720/A vssd1 vssd1 vccd1 vccd1 hold720/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 hold731/A vssd1 vssd1 vccd1 vccd1 hold731/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold742 hold742/A vssd1 vssd1 vccd1 vccd1 hold742/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23022_ _23020_/X _23021_/Y _22856_/X vssd1 vssd1 vccd1 vccd1 _25890_/D sky130_fd_sc_hd__a21oi_1
Xhold753 hold753/A vssd1 vssd1 vccd1 vccd1 hold753/X sky130_fd_sc_hd__dlygate4sd3_1
X_20234_ _20232_/Y _20233_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _20234_/Y sky130_fd_sc_hd__a21oi_1
Xhold764 hold764/A vssd1 vssd1 vccd1 vccd1 hold764/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold775 hold775/A vssd1 vssd1 vccd1 vccd1 hold775/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 hold786/A vssd1 vssd1 vccd1 vccd1 hold786/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 hold797/A vssd1 vssd1 vccd1 vccd1 hold797/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20165_ _20165_/A _25881_/Q vssd1 vssd1 vccd1 vccd1 _20171_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_110_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2110 _26132_/Q vssd1 vssd1 vccd1 vccd1 hold2110/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2121 _23835_/X vssd1 vssd1 vccd1 vccd1 _23836_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2132 _25001_/Q vssd1 vssd1 vccd1 vccd1 _12522_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24973_ _25425_/CLK _24973_/D vssd1 vssd1 vccd1 vccd1 _24973_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2143 _23745_/X vssd1 vssd1 vccd1 vccd1 _23746_/A sky130_fd_sc_hd__dlygate4sd3_1
X_20096_ _20096_/A _20096_/B vssd1 vssd1 vccd1 vccd1 _21709_/A sky130_fd_sc_hd__nand2_4
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2154 _24249_/X vssd1 vssd1 vccd1 vccd1 _24250_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2165 _26013_/Q vssd1 vssd1 vccd1 vccd1 hold2165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1420 _13346_/X vssd1 vssd1 vccd1 vccd1 _25109_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2176 _24311_/X vssd1 vssd1 vccd1 vccd1 _24312_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1431 _25747_/Q vssd1 vssd1 vccd1 vccd1 _19652_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23924_ _23924_/A _24968_/Q _23924_/C vssd1 vssd1 vccd1 vccd1 _23924_/Y sky130_fd_sc_hd__nor3_1
Xhold1442 _21155_/Y vssd1 vssd1 vccd1 vccd1 _25806_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2187 _26165_/Q vssd1 vssd1 vccd1 vccd1 hold2187/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2198 _15011_/Y vssd1 vssd1 vccd1 vccd1 _25425_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1453 _25765_/Q vssd1 vssd1 vccd1 vccd1 _19904_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1464 _19425_/Y vssd1 vssd1 vccd1 vccd1 _25731_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1475 _25799_/Q vssd1 vssd1 vccd1 vccd1 _20962_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1486 _23134_/Y vssd1 vssd1 vccd1 vccd1 _25897_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23855_ _23855_/A vssd1 vssd1 vccd1 vccd1 _26022_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1497 _25818_/Q vssd1 vssd1 vccd1 vccd1 _21412_/B sky130_fd_sc_hd__buf_1
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22806_ _22804_/X _22805_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22806_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23786_ _23786_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23787_/A sky130_fd_sc_hd__and2_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20998_ _20998_/A _22011_/B _20998_/C vssd1 vssd1 vccd1 vccd1 _21002_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_184_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25525_ _26012_/CLK hold941/X vssd1 vssd1 vccd1 vccd1 hold940/A sky130_fd_sc_hd__dfxtp_1
X_22737_ _16790_/B _22421_/X _22731_/X _22732_/Y _22736_/X vssd1 vssd1 vccd1 vccd1
+ _22738_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_165_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25456_ _26064_/CLK hold917/X vssd1 vssd1 vccd1 vccd1 hold916/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13470_ _13470_/A _13518_/B vssd1 vssd1 vccd1 vccd1 _13470_/Y sky130_fd_sc_hd__nor2_1
X_22668_ _25707_/Q _22667_/A _22667_/Y vssd1 vssd1 vccd1 vccd1 _22670_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_164_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24407_ _24407_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24408_/A sky130_fd_sc_hd__and2_1
XFILLER_0_35_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21619_ _21618_/Y _21203_/X _20986_/A _20957_/A vssd1 vssd1 vccd1 vccd1 _21619_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_180_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25387_ _26339_/CLK hold319/X vssd1 vssd1 vccd1 vccd1 hold317/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22599_ _22957_/B _23104_/B vssd1 vssd1 vccd1 vccd1 _22600_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15140_ _22476_/B _16369_/B vssd1 vssd1 vccd1 vccd1 _15141_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24338_ hold2404/X _26178_/Q _24356_/S vssd1 vssd1 vccd1 vccd1 _24338_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_105_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15071_ _15270_/A _15108_/A _15110_/A vssd1 vssd1 vccd1 vccd1 _15073_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_132_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24269_ _24269_/A vssd1 vssd1 vccd1 vccd1 _26155_/D sky130_fd_sc_hd__clkbuf_1
X_26008_ _26009_/CLK _26008_/D vssd1 vssd1 vccd1 vccd1 _26008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14022_ _18139_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14022_/Y sky130_fd_sc_hd__nor2_1
X_18830_ _18952_/A _25767_/Q _18891_/C vssd1 vssd1 vccd1 vccd1 _18831_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_101_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15973_ _15999_/A vssd1 vssd1 vccd1 vccd1 _15978_/B sky130_fd_sc_hd__inv_2
X_18761_ _18761_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18761_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_175_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14924_ _14924_/A _14923_/Y vssd1 vssd1 vccd1 vccd1 _14927_/B sky130_fd_sc_hd__or2b_1
X_17712_ _17721_/A _25904_/Q vssd1 vssd1 vccd1 vccd1 _17719_/A sky130_fd_sc_hd__nand2_1
X_18692_ _18792_/A _25760_/Q vssd1 vssd1 vccd1 vccd1 _18694_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_175_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14855_ _25855_/Q _14170_/A _15042_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14856_/B
+ sky130_fd_sc_hd__a22o_1
X_17643_ _17641_/Y _17642_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _17643_/Y sky130_fd_sc_hd__a21oi_1
X_13806_ hold618/X _13805_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold619/A sky130_fd_sc_hd__a21oi_1
X_17574_ _17574_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17574_/Y sky130_fd_sc_hd__nand2_1
X_14786_ _14900_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14786_/Y sky130_fd_sc_hd__nand2_1
X_16525_ _16512_/A _16500_/A _16511_/B vssd1 vssd1 vccd1 vccd1 _16525_/Y sky130_fd_sc_hd__a21oi_1
X_19313_ _26227_/Q _12537_/B hold446/X vssd1 vssd1 vccd1 vccd1 _19313_/Y sky130_fd_sc_hd__a21oi_1
X_13737_ _25753_/Q vssd1 vssd1 vccd1 vccd1 _18550_/B sky130_fd_sc_hd__inv_2
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_70_clk _25472_/CLK vssd1 vssd1 vccd1 vccd1 _26066_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16456_ _16456_/A _16456_/B vssd1 vssd1 vccd1 vccd1 _16456_/Y sky130_fd_sc_hd__nand2_1
X_19244_ _19244_/A _20586_/B vssd1 vssd1 vccd1 vccd1 _19244_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_45_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13668_ _13760_/A hold791/X vssd1 vssd1 vccd1 vccd1 hold792/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15407_ _15408_/B _15407_/B vssd1 vssd1 vccd1 vccd1 _15822_/B sky130_fd_sc_hd__and2_1
XFILLER_0_54_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12619_ _12624_/A _24836_/B _12619_/C vssd1 vssd1 vccd1 vccd1 _12620_/A sky130_fd_sc_hd__and3_1
XFILLER_0_26_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19175_ _19175_/A _19980_/B _19175_/C vssd1 vssd1 vccd1 vccd1 _19175_/X sky130_fd_sc_hd__and3_1
XFILLER_0_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16387_ _16387_/A _16401_/C vssd1 vssd1 vccd1 vccd1 _16390_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13599_ _25731_/Q vssd1 vssd1 vccd1 vccd1 _18002_/B sky130_fd_sc_hd__inv_2
XFILLER_0_171_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18126_ _18126_/A _20290_/B vssd1 vssd1 vccd1 vccd1 _20284_/A sky130_fd_sc_hd__nand2_4
X_15338_ hold975/X _15340_/A vssd1 vssd1 vccd1 vccd1 _15342_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_83_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18057_ _19053_/A _18057_/B vssd1 vssd1 vccd1 vccd1 _18057_/X sky130_fd_sc_hd__xor2_1
X_15269_ _15272_/B _15269_/B _15271_/B vssd1 vssd1 vccd1 vccd1 _15270_/B sky130_fd_sc_hd__and3_1
XFILLER_0_124_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17008_ _17008_/A _17008_/B vssd1 vssd1 vccd1 vccd1 _17009_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18959_ _19031_/A _19080_/B vssd1 vssd1 vccd1 vccd1 _18960_/B sky130_fd_sc_hd__xnor2_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21970_ _21970_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _21970_/X sky130_fd_sc_hd__and2_1
XFILLER_0_179_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20921_ _20921_/A _20921_/B _21435_/B vssd1 vssd1 vccd1 vccd1 _20925_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23640_ _23640_/A vssd1 vssd1 vccd1 vccd1 _25952_/D sky130_fd_sc_hd__clkbuf_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20852_ _20852_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _20852_/Y sky130_fd_sc_hd__nand2_1
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23571_ _23568_/Y _23570_/Y _24957_/S vssd1 vssd1 vccd1 vccd1 _23571_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20783_ _25858_/Q vssd1 vssd1 vccd1 vccd1 _21769_/B sky130_fd_sc_hd__inv_2
XFILLER_0_14_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_61_clk _25472_/CLK vssd1 vssd1 vccd1 vccd1 _25537_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25310_ _26139_/CLK hold19/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22522_ _22907_/B _23056_/B vssd1 vssd1 vccd1 vccd1 _22523_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_119_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26290_ _26292_/CLK _26290_/D vssd1 vssd1 vccd1 vccd1 _26290_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_119_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25241_ _25817_/CLK hold840/X vssd1 vssd1 vccd1 vccd1 hold839/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22453_ _22453_/A _22453_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22456_/A sky130_fd_sc_hd__or3_1
XFILLER_0_134_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21404_ _21404_/A _21404_/B vssd1 vssd1 vccd1 vccd1 _21405_/A sky130_fd_sc_hd__nand2_1
X_25172_ _25779_/CLK hold382/X vssd1 vssd1 vccd1 vccd1 hold380/A sky130_fd_sc_hd__dfxtp_1
X_22384_ _22561_/A _22384_/B vssd1 vssd1 vccd1 vccd1 _22384_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_60_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24123_ hold2145/X _26108_/Q _24126_/S vssd1 vssd1 vccd1 vccd1 _24123_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21335_ _21335_/A _21335_/B _21335_/C vssd1 vssd1 vccd1 vccd1 _21339_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_20_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24054_ _24054_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24055_/A sky130_fd_sc_hd__and2_1
Xhold550 hold550/A vssd1 vssd1 vccd1 vccd1 hold550/X sky130_fd_sc_hd__dlygate4sd3_1
X_21266_ _21268_/B _21268_/C vssd1 vssd1 vccd1 vccd1 _21267_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_130_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold561 hold561/A vssd1 vssd1 vccd1 vccd1 hold561/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 hold572/A vssd1 vssd1 vccd1 vccd1 hold572/X sky130_fd_sc_hd__dlygate4sd3_1
X_23005_ _23197_/A _23005_/B vssd1 vssd1 vccd1 vccd1 _23005_/Y sky130_fd_sc_hd__nand2_1
Xhold583 hold583/A vssd1 vssd1 vccd1 vccd1 hold583/X sky130_fd_sc_hd__dlygate4sd3_1
X_20217_ _20216_/B _20217_/B _20217_/C vssd1 vssd1 vccd1 vccd1 _20218_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_99_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold594 hold594/A vssd1 vssd1 vccd1 vccd1 hold594/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21197_ _21643_/C _21594_/C vssd1 vssd1 vccd1 vccd1 _21198_/C sky130_fd_sc_hd__nand2_1
X_20148_ _20148_/A _21036_/B _20148_/C vssd1 vssd1 vccd1 vccd1 _20151_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_99_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24956_ _16678_/B _16692_/A _24956_/S vssd1 vssd1 vccd1 vccd1 _24956_/X sky130_fd_sc_hd__mux2_1
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ _12930_/X _12968_/X _12917_/X _12969_/X vssd1 vssd1 vccd1 vccd1 _12970_/X
+ sky130_fd_sc_hd__o211a_1
X_20079_ _26278_/Q _20078_/X hold602/X vssd1 vssd1 vccd1 vccd1 _20082_/B sky130_fd_sc_hd__a21oi_1
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1250 _25100_/Q vssd1 vssd1 vccd1 vccd1 _18719_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1261 _16920_/Y vssd1 vssd1 vccd1 vccd1 _25571_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23907_ hold2003/X hold1912/X _23907_/S vssd1 vssd1 vccd1 vccd1 _23909_/A sky130_fd_sc_hd__mux2_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1272 _25112_/Q vssd1 vssd1 vccd1 vccd1 _18961_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24887_ _24887_/A _24946_/A vssd1 vssd1 vccd1 vccd1 _24887_/Y sky130_fd_sc_hd__nand2_1
Xhold1283 _16852_/Y vssd1 vssd1 vccd1 vccd1 _25561_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1294 _25563_/Q vssd1 vssd1 vccd1 vccd1 _16865_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _14638_/Y hold33/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_185_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23838_ hold2238/X hold2119/X _23907_/S vssd1 vssd1 vccd1 vccd1 _23839_/A sky130_fd_sc_hd__mux2_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _14569_/Y hold120/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold121/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23769_ _23769_/A vssd1 vssd1 vccd1 vccd1 _25994_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _26012_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_184_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16310_ _16296_/A _16284_/A _16295_/B vssd1 vssd1 vccd1 vccd1 _16310_/X sky130_fd_sc_hd__a21o_1
X_25508_ _25510_/CLK hold703/X vssd1 vssd1 vccd1 vccd1 hold701/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13522_ _13522_/A hold533/X vssd1 vssd1 vccd1 vccd1 hold534/A sky130_fd_sc_hd__nand2_1
X_17290_ _19416_/A _17290_/B vssd1 vssd1 vccd1 vccd1 _17556_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_94_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16241_ _16239_/X _16240_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _16241_/X sky130_fd_sc_hd__a21o_1
X_25439_ _26002_/CLK _25439_/D vssd1 vssd1 vccd1 vccd1 _25439_/Q sky130_fd_sc_hd__dfxtp_1
X_13453_ _26339_/Q _25708_/Q vssd1 vssd1 vccd1 vccd1 _14684_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_152_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16172_ _16216_/A _16172_/B vssd1 vssd1 vccd1 vccd1 _16182_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_153_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13384_ _26327_/Q _19744_/A vssd1 vssd1 vccd1 vccd1 _14648_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15123_ _15123_/A _16712_/A vssd1 vssd1 vccd1 vccd1 _15124_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_106_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15054_ _15067_/A _15055_/A vssd1 vssd1 vccd1 vccd1 _15054_/X sky130_fd_sc_hd__or2_1
X_19931_ _19975_/A _19931_/B vssd1 vssd1 vccd1 vccd1 _19931_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_120_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14005_ _14061_/A _14005_/B vssd1 vssd1 vccd1 vccd1 _14005_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_103_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19862_ _19862_/A _19862_/B vssd1 vssd1 vccd1 vccd1 _19862_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18813_ _18955_/A _18813_/B _18894_/C vssd1 vssd1 vccd1 vccd1 _18814_/C sky130_fd_sc_hd__nand3_1
X_19793_ _19793_/A _19793_/B vssd1 vssd1 vccd1 vccd1 _19793_/Y sky130_fd_sc_hd__nand2_1
X_18744_ _19788_/A vssd1 vssd1 vccd1 vccd1 _22463_/B sky130_fd_sc_hd__inv_2
X_15956_ _15956_/A hold880/X vssd1 vssd1 vccd1 vccd1 _15956_/Y sky130_fd_sc_hd__nand2_1
X_14907_ _14916_/B _14907_/B vssd1 vssd1 vccd1 vccd1 _14907_/Y sky130_fd_sc_hd__xnor2_1
X_15887_ _15885_/X hold462/X _15805_/X vssd1 vssd1 vccd1 vccd1 hold463/A sky130_fd_sc_hd__a21oi_1
X_18675_ _20409_/B _22372_/A vssd1 vssd1 vccd1 vccd1 _20400_/A sky130_fd_sc_hd__nand2_2
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17626_ _17626_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _17626_/Y sky130_fd_sc_hd__nand2_1
X_14838_ _25853_/Q _13466_/A _14837_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14839_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14769_ _14767_/Y _14768_/Y _14741_/X vssd1 vssd1 vccd1 vccd1 _14769_/Y sky130_fd_sc_hd__a21oi_1
X_17557_ _17624_/A _17557_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17557_/X sky130_fd_sc_hd__and3_1
XFILLER_0_74_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_43_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _26079_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16508_ hold940/X vssd1 vssd1 vccd1 vccd1 _16508_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_73_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17488_ _17488_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17488_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19227_ _19227_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _19227_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_183_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16439_ _16441_/B _16439_/B vssd1 vssd1 vccd1 vccd1 _16439_/X sky130_fd_sc_hd__or2_1
XFILLER_0_143_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19158_ _25650_/Q _20174_/B vssd1 vssd1 vccd1 vccd1 _19158_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_171_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18109_ _18109_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _18109_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19089_ _19089_/A _19089_/B vssd1 vssd1 vccd1 vccd1 _20023_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21120_ _26308_/Q _20731_/X hold620/X vssd1 vssd1 vccd1 vccd1 _21123_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_160_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21051_ _25867_/Q _21051_/B _21051_/C vssd1 vssd1 vccd1 vccd1 _21054_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_100_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20002_ _23165_/B vssd1 vssd1 vccd1 vccd1 _22670_/B sky130_fd_sc_hd__inv_2
X_24810_ _24810_/A vssd1 vssd1 vccd1 vccd1 _26331_/D sky130_fd_sc_hd__clkbuf_1
X_25790_ _25793_/CLK _25790_/D vssd1 vssd1 vccd1 vccd1 _25790_/Q sky130_fd_sc_hd__dfxtp_2
X_24741_ _24741_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24742_/A sky130_fd_sc_hd__and2_1
X_21953_ _21953_/A _21953_/B vssd1 vssd1 vccd1 vccd1 _22703_/A sky130_fd_sc_hd__nand2_2
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20904_ _20904_/A _20904_/B vssd1 vssd1 vccd1 vccd1 _20905_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24672_ _24672_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24673_/A sky130_fd_sc_hd__and2_1
X_21884_ _21884_/A _21884_/B vssd1 vssd1 vccd1 vccd1 _22651_/A sky130_fd_sc_hd__nand2_2
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23623_ _23623_/A _23629_/B vssd1 vssd1 vccd1 vccd1 _23624_/A sky130_fd_sc_hd__and2_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20835_ _20835_/A _20835_/B vssd1 vssd1 vccd1 vccd1 _20837_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_178_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_clk _25184_/CLK vssd1 vssd1 vccd1 vccd1 _25765_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23554_ _23548_/X _23553_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _23554_/X sky130_fd_sc_hd__mux2_1
X_20766_ _21403_/B _21677_/B vssd1 vssd1 vccd1 vccd1 _20767_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22505_ _22504_/A _22454_/X _22504_/B vssd1 vssd1 vccd1 vccd1 _22506_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26273_ _26273_/CLK _26273_/D vssd1 vssd1 vccd1 vccd1 _26273_/Q sky130_fd_sc_hd__dfxtp_1
X_23485_ hold110/A _24860_/S vssd1 vssd1 vccd1 vccd1 _23485_/X sky130_fd_sc_hd__or2b_1
X_20697_ _20697_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _20697_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25224_ _25678_/CLK hold797/X vssd1 vssd1 vccd1 vccd1 hold796/A sky130_fd_sc_hd__dfxtp_1
X_22436_ _25826_/Q _22436_/B vssd1 vssd1 vccd1 vccd1 _22436_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25155_ _25738_/CLK hold496/X vssd1 vssd1 vccd1 vccd1 hold494/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22367_ _22365_/X _15839_/B _22366_/Y _14891_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _22368_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_102_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24106_ _24106_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24107_/A sky130_fd_sc_hd__and2_1
X_21318_ _21369_/A _21675_/C vssd1 vssd1 vccd1 vccd1 _21319_/B sky130_fd_sc_hd__nand2_1
X_25086_ _26299_/CLK _25086_/D vssd1 vssd1 vccd1 vccd1 _25086_/Q sky130_fd_sc_hd__dfxtp_1
X_22298_ _18615_/A _25820_/Q _22296_/Y _22297_/Y vssd1 vssd1 vccd1 vccd1 _22299_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_102_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24037_ _24037_/A vssd1 vssd1 vccd1 vccd1 _26080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21249_ _21249_/A _21249_/B _21249_/C vssd1 vssd1 vccd1 vccd1 _21253_/A sky130_fd_sc_hd__nand3_1
Xhold380 hold380/A vssd1 vssd1 vccd1 vccd1 hold380/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 hold391/A vssd1 vssd1 vccd1 vccd1 hold391/X sky130_fd_sc_hd__dlygate4sd3_1
X_15810_ _15810_/A _15810_/B vssd1 vssd1 vccd1 vccd1 _15811_/B sky130_fd_sc_hd__nand2_2
X_16790_ _16858_/A _16790_/B vssd1 vssd1 vccd1 vccd1 _16790_/Y sky130_fd_sc_hd__nand2_1
X_25988_ _25991_/CLK _25988_/D vssd1 vssd1 vccd1 vccd1 _25988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15741_ _15795_/A _16638_/B vssd1 vssd1 vccd1 vccd1 _15744_/A sky130_fd_sc_hd__nor2_1
X_24939_ _24867_/S _24932_/Y _24934_/Y _24938_/X vssd1 vssd1 vccd1 vccd1 _24939_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ _26124_/Q _12907_/X _12952_/X vssd1 vssd1 vccd1 vccd1 _12953_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_88_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1080 _12950_/X vssd1 vssd1 vccd1 vccd1 _25040_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1091 _25070_/Q vssd1 vssd1 vccd1 vccd1 _18008_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15672_ _15673_/B _16923_/A vssd1 vssd1 vccd1 vccd1 _15674_/A sky130_fd_sc_hd__nor2_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18460_ _19588_/A vssd1 vssd1 vccd1 vccd1 _22095_/B sky130_fd_sc_hd__inv_2
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _17363_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12884_/X sky130_fd_sc_hd__or2_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _19574_/A _17411_/B vssd1 vssd1 vccd1 vccd1 _17637_/B sky130_fd_sc_hd__xor2_4
X_14623_ _14623_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14623_/Y sky130_fd_sc_hd__nand2_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18391_ _18596_/A _18738_/A vssd1 vssd1 vccd1 vccd1 _18392_/B sky130_fd_sc_hd__xnor2_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _25779_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17342_ _17616_/A _17342_/B vssd1 vssd1 vccd1 vccd1 _17342_/X sky130_fd_sc_hd__xor2_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14554_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14554_/Y sky130_fd_sc_hd__nand2_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13505_ _25716_/Q vssd1 vssd1 vccd1 vccd1 _18070_/B sky130_fd_sc_hd__inv_2
X_17273_ _17271_/Y _17272_/Y _17204_/X vssd1 vssd1 vccd1 vccd1 _17273_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14485_ _14485_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14485_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16224_ _16224_/A _16224_/B vssd1 vssd1 vccd1 vccd1 _16225_/B sky130_fd_sc_hd__nand2_1
X_19012_ _19026_/A hold995/X _22786_/A vssd1 vssd1 vccd1 vccd1 _19012_/X sky130_fd_sc_hd__and3_1
XFILLER_0_10_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13436_ _19047_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13436_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16155_ _16153_/X _16154_/Y _16076_/X vssd1 vssd1 vccd1 vccd1 hold862/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13367_ _13220_/X _14638_/A _13242_/X _19701_/A vssd1 vssd1 vccd1 vccd1 _13367_/X
+ sky130_fd_sc_hd__a22o_1
X_15106_ _15106_/A _15106_/B vssd1 vssd1 vccd1 vccd1 _15107_/A sky130_fd_sc_hd__or2_1
X_16086_ _16160_/A _16104_/A _16107_/A vssd1 vssd1 vccd1 vccd1 _16088_/A sky130_fd_sc_hd__a21o_1
X_13298_ _26185_/Q _13239_/X _13297_/X vssd1 vssd1 vccd1 vccd1 _13298_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_122_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15037_ _15037_/A _15037_/B vssd1 vssd1 vccd1 vccd1 _15270_/A sky130_fd_sc_hd__nand2_4
X_19914_ _19914_/A _19914_/B vssd1 vssd1 vccd1 vccd1 _19914_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_20_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2709 _24575_/X vssd1 vssd1 vccd1 vccd1 _24576_/A sky130_fd_sc_hd__dlygate4sd3_1
X_19845_ _20711_/A _22564_/B _25639_/Q vssd1 vssd1 vccd1 vccd1 _20716_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_120_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19776_ _20517_/A _19774_/Y _20522_/C vssd1 vssd1 vccd1 vccd1 _19862_/B sky130_fd_sc_hd__o21a_2
X_16988_ _18147_/B _16988_/B vssd1 vssd1 vccd1 vccd1 _17402_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18727_ _18727_/A _18727_/B vssd1 vssd1 vccd1 vccd1 _22435_/A sky130_fd_sc_hd__nand2_1
X_15939_ _15937_/X hold444/X _15805_/X vssd1 vssd1 vccd1 vccd1 hold445/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18658_ _19026_/A _18658_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18658_/X sky130_fd_sc_hd__and3_1
XFILLER_0_94_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17609_ _17624_/A _17609_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _17609_/X sky130_fd_sc_hd__and3_1
XFILLER_0_148_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18589_ _18589_/A _25819_/Q _18589_/C vssd1 vssd1 vccd1 vccd1 _20244_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_clk _25184_/CLK vssd1 vssd1 vccd1 vccd1 _25711_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20620_ _20620_/A _20620_/B vssd1 vssd1 vccd1 vccd1 _20621_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20551_ _20551_/A _22195_/B _20551_/C vssd1 vssd1 vccd1 vccd1 _20554_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_74_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23270_ _23270_/A _23377_/B _23270_/C vssd1 vssd1 vccd1 vccd1 _23271_/A sky130_fd_sc_hd__and3_1
XFILLER_0_144_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20482_ _23005_/B vssd1 vssd1 vccd1 vccd1 _22413_/B sky130_fd_sc_hd__inv_2
XFILLER_0_14_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22221_ _22221_/A _22221_/B vssd1 vssd1 vccd1 vccd1 _22221_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22152_ _19616_/A _22151_/A _22151_/Y vssd1 vssd1 vccd1 vccd1 _22154_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_140_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21103_ _21105_/B _21105_/C vssd1 vssd1 vccd1 vccd1 _21104_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22083_ _22084_/A _22084_/C _23058_/A vssd1 vssd1 vccd1 vccd1 _22083_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_121_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25911_ _25913_/CLK _25911_/D vssd1 vssd1 vccd1 vccd1 _25911_/Q sky130_fd_sc_hd__dfxtp_1
X_21034_ _21545_/C _21500_/B vssd1 vssd1 vccd1 vccd1 _21036_/A sky130_fd_sc_hd__nand2_1
X_25842_ _26339_/CLK _25842_/D vssd1 vssd1 vccd1 vccd1 _25842_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_96_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25773_ _25773_/CLK _25773_/D vssd1 vssd1 vccd1 vccd1 _25773_/Q sky130_fd_sc_hd__dfxtp_1
X_22985_ _16893_/B _22421_/X _22979_/X _22980_/Y _22984_/X vssd1 vssd1 vccd1 vccd1
+ _22986_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_69_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24724_ _24724_/A vssd1 vssd1 vccd1 vccd1 _26303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21936_ _21936_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _21936_/X sky130_fd_sc_hd__and2_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24655_ hold2620/X _26281_/Q _24664_/S vssd1 vssd1 vccd1 vccd1 _24655_/X sky130_fd_sc_hd__mux2_1
X_21867_ _21867_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _21867_/X sky130_fd_sc_hd__and2_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23606_ _23606_/A vssd1 vssd1 vccd1 vccd1 _25941_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20818_ _20818_/A _20818_/B vssd1 vssd1 vccd1 vccd1 _20822_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24586_ _24586_/A vssd1 vssd1 vccd1 vccd1 _26258_/D sky130_fd_sc_hd__clkbuf_1
X_21798_ _21796_/X _14270_/A _21797_/Y _14721_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _21799_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_93_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26325_ _26325_/CLK _26325_/D vssd1 vssd1 vccd1 vccd1 _26325_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23537_ _23534_/Y _23536_/Y _24957_/S vssd1 vssd1 vccd1 vccd1 _23537_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_181_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20749_ _20749_/A _20749_/B vssd1 vssd1 vccd1 vccd1 _21403_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14270_ _14270_/A _14270_/B vssd1 vssd1 vccd1 vccd1 _14270_/Y sky130_fd_sc_hd__nor2_1
X_26256_ _26267_/CLK _26256_/D vssd1 vssd1 vccd1 vccd1 _26256_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_92_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23468_ _23465_/Y _23467_/Y _24957_/S vssd1 vssd1 vccd1 vccd1 _23468_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25207_ _26289_/CLK hold730/X vssd1 vssd1 vccd1 vccd1 hold728/A sky130_fd_sc_hd__dfxtp_1
X_13221_ _13221_/A vssd1 vssd1 vccd1 vccd1 _19373_/A sky130_fd_sc_hd__buf_4
X_22419_ _23120_/A _22419_/B vssd1 vssd1 vccd1 vccd1 _22420_/A sky130_fd_sc_hd__xor2_1
X_26187_ _26190_/CLK _26187_/D vssd1 vssd1 vccd1 vccd1 _26187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23399_ _24940_/S hold188/A _23398_/X vssd1 vssd1 vccd1 vccd1 _23399_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25138_ _26239_/CLK hold844/X vssd1 vssd1 vccd1 vccd1 hold843/A sky130_fd_sc_hd__dfxtp_1
X_13152_ _13152_/A vssd1 vssd1 vccd1 vccd1 _19216_/A sky130_fd_sc_hd__buf_4
XFILLER_0_104_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17960_ _17960_/A _20779_/A vssd1 vssd1 vccd1 vccd1 _18434_/A sky130_fd_sc_hd__xor2_4
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25069_ _26152_/CLK _25069_/D vssd1 vssd1 vccd1 vccd1 _25069_/Q sky130_fd_sc_hd__dfxtp_1
X_13083_ _26277_/Q _21749_/A vssd1 vssd1 vccd1 vccd1 _14491_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_103_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16911_ _16911_/A _16911_/B vssd1 vssd1 vccd1 vccd1 _16911_/Y sky130_fd_sc_hd__nand2_1
X_17891_ _18529_/C vssd1 vssd1 vccd1 vccd1 _18955_/C sky130_fd_sc_hd__buf_8
XFILLER_0_109_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19630_ _19630_/A _20132_/B vssd1 vssd1 vccd1 vccd1 _19630_/Y sky130_fd_sc_hd__nor2_1
X_16842_ _16980_/A _16842_/B vssd1 vssd1 vccd1 vccd1 _16842_/Y sky130_fd_sc_hd__nand2_1
X_19561_ _21264_/A _22040_/B _25619_/Q vssd1 vssd1 vccd1 vccd1 _21268_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_189_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16773_ _16773_/A vssd1 vssd1 vccd1 vccd1 _16977_/A sky130_fd_sc_hd__clkbuf_8
X_13985_ _14061_/A _13985_/B vssd1 vssd1 vccd1 vccd1 _13985_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18512_ _18512_/A _20098_/A vssd1 vssd1 vccd1 vccd1 _18858_/A sky130_fd_sc_hd__xor2_4
X_15724_ _23111_/B _15724_/B vssd1 vssd1 vccd1 vccd1 _23108_/B sky130_fd_sc_hd__xor2_1
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12936_ _26249_/Q _25618_/Q vssd1 vssd1 vccd1 vccd1 _14400_/A sky130_fd_sc_hd__xor2_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19492_ _19493_/B _19493_/A vssd1 vssd1 vccd1 vccd1 _19492_/X sky130_fd_sc_hd__or2_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18443_ _18443_/A _18443_/B vssd1 vssd1 vccd1 vccd1 _22064_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_185_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15655_ _15655_/A vssd1 vssd1 vccd1 vccd1 _15656_/B sky130_fd_sc_hd__inv_2
X_12867_ _12726_/B _14361_/A _12752_/X _25605_/Q vssd1 vssd1 vccd1 vccd1 _12867_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14606_ _14645_/A hold293/X vssd1 vssd1 vccd1 vccd1 hold294/A sky130_fd_sc_hd__nand2_1
X_15586_ hold908/X _15588_/A vssd1 vssd1 vccd1 vccd1 _15590_/A sky130_fd_sc_hd__nor2_1
X_18374_ _18372_/X _18269_/X _18373_/X vssd1 vssd1 vccd1 vccd1 _18375_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12798_ _26223_/Q _25592_/Q vssd1 vssd1 vccd1 vccd1 _14319_/A sky130_fd_sc_hd__xor2_2
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _17467_/A _17325_/B vssd1 vssd1 vccd1 vccd1 _17325_/Y sky130_fd_sc_hd__nand2_1
X_14537_ _14585_/A hold269/X vssd1 vssd1 vccd1 vccd1 hold270/A sky130_fd_sc_hd__nand2_1
XFILLER_0_154_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17256_ _17393_/A _17256_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17256_/X sky130_fd_sc_hd__and3_1
X_14468_ _14588_/A vssd1 vssd1 vccd1 vccd1 _14524_/B sky130_fd_sc_hd__buf_8
XFILLER_0_71_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16207_ _16207_/A vssd1 vssd1 vccd1 vccd1 _16214_/B sky130_fd_sc_hd__inv_2
X_13419_ _14125_/A vssd1 vssd1 vccd1 vccd1 _13522_/A sky130_fd_sc_hd__buf_8
X_17187_ _17393_/A _17187_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17187_/X sky130_fd_sc_hd__and3_1
XFILLER_0_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14399_ _14397_/Y hold285/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold286/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_141_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16138_ _16139_/B _16139_/A vssd1 vssd1 vccd1 vccd1 _16150_/B sky130_fd_sc_hd__or2_1
XFILLER_0_51_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16069_ _16069_/A _16069_/B vssd1 vssd1 vccd1 vccd1 _16070_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _25636_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2506 _25697_/Q vssd1 vssd1 vccd1 vccd1 _13389_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2517 _12635_/Y vssd1 vssd1 vccd1 vccd1 _12636_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold2528 _15183_/Y vssd1 vssd1 vccd1 vccd1 _25439_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2539 _24991_/Q vssd1 vssd1 vccd1 vccd1 _12694_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1805 _25636_/Q vssd1 vssd1 vccd1 vccd1 _17591_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1816 _21898_/Y vssd1 vssd1 vccd1 vccd1 _25842_/D sky130_fd_sc_hd__dlygate4sd3_1
X_19828_ _19827_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19829_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1827 _25850_/Q vssd1 vssd1 vccd1 vccd1 _22142_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1838 _22089_/Y vssd1 vssd1 vccd1 vccd1 _25848_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1849 _23595_/X vssd1 vssd1 vccd1 vccd1 _25940_/D sky130_fd_sc_hd__dlygate4sd3_1
X_19759_ _20478_/A _22408_/B _25633_/Q vssd1 vssd1 vccd1 vccd1 _20483_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_79_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22770_ _22770_/A _22900_/B vssd1 vssd1 vccd1 vccd1 _22770_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21721_ _22893_/A _21721_/B vssd1 vssd1 vccd1 vccd1 _21721_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24440_ hold1938/X _26211_/Q _24510_/S vssd1 vssd1 vccd1 vccd1 _24440_/X sky130_fd_sc_hd__mux2_1
X_21652_ _21716_/A _21652_/B _21651_/X vssd1 vssd1 vccd1 vccd1 _21653_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20603_ _20605_/B vssd1 vssd1 vccd1 vccd1 _20604_/B sky130_fd_sc_hd__inv_2
XFILLER_0_117_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24371_ _24371_/A vssd1 vssd1 vccd1 vccd1 _26188_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21583_ _26332_/Q _19130_/X hold751/X vssd1 vssd1 vccd1 vccd1 _21586_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26110_ _26112_/CLK _26110_/D vssd1 vssd1 vccd1 vccd1 _26110_/Q sky130_fd_sc_hd__dfxtp_1
X_23322_ _23322_/A vssd1 vssd1 vccd1 vccd1 _25926_/D sky130_fd_sc_hd__clkbuf_1
X_20534_ _20534_/A _21225_/B _20534_/C vssd1 vssd1 vccd1 vccd1 _20535_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26041_ _26041_/CLK _26041_/D vssd1 vssd1 vccd1 vccd1 _26041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23253_ _24959_/C _24867_/S _23253_/C vssd1 vssd1 vccd1 vccd1 _23256_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_104_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20465_ _21099_/A vssd1 vssd1 vccd1 vccd1 _20465_/X sky130_fd_sc_hd__buf_6
XFILLER_0_43_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22204_ _22204_/A _22387_/B vssd1 vssd1 vccd1 vccd1 _22204_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_162_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23184_ _23184_/A _23184_/B vssd1 vssd1 vccd1 vccd1 _23185_/B sky130_fd_sc_hd__nand2_1
X_20396_ _20396_/A _20396_/B vssd1 vssd1 vccd1 vccd1 _20398_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22135_ _22136_/B _22136_/A vssd1 vssd1 vccd1 vccd1 _22137_/A sky130_fd_sc_hd__or2_2
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22066_ _18452_/A _25812_/Q _22064_/Y _22065_/Y vssd1 vssd1 vccd1 vccd1 _22067_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21017_ _21017_/A _21017_/B vssd1 vssd1 vccd1 vccd1 _21018_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25825_ _25827_/CLK _25825_/D vssd1 vssd1 vccd1 vccd1 _25825_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_173_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13770_ _18652_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13770_/Y sky130_fd_sc_hd__nor2_1
X_25756_ _25756_/CLK _25756_/D vssd1 vssd1 vccd1 vccd1 _25756_/Q sky130_fd_sc_hd__dfxtp_1
X_22968_ _16886_/B _22421_/X _22962_/X _22963_/Y _22967_/X vssd1 vssd1 vccd1 vccd1
+ _22969_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_139_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12721_ _19483_/A vssd1 vssd1 vccd1 vccd1 _12721_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_179_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21919_ _21919_/A _21919_/B vssd1 vssd1 vccd1 vccd1 _22676_/A sky130_fd_sc_hd__nand2_2
X_24707_ hold2580/X _26298_/Q _24740_/S vssd1 vssd1 vccd1 vccd1 _24707_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25687_ _25687_/CLK _25687_/D vssd1 vssd1 vccd1 vccd1 _25687_/Q sky130_fd_sc_hd__dfxtp_1
X_22899_ _16858_/B _22421_/X _22893_/X _22894_/Y _22898_/X vssd1 vssd1 vccd1 vccd1
+ _22900_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15440_ _15440_/A vssd1 vssd1 vccd1 vccd1 _15441_/B sky130_fd_sc_hd__inv_2
X_12652_ _12652_/A _24836_/B _12661_/B vssd1 vssd1 vccd1 vccd1 _12652_/X sky130_fd_sc_hd__and3_1
X_24638_ _24638_/A vssd1 vssd1 vccd1 vccd1 _26275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15371_ _15373_/B _16810_/A vssd1 vssd1 vccd1 vccd1 _15372_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_154_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12583_ _12587_/A _14910_/B _12583_/C vssd1 vssd1 vccd1 vccd1 _12583_/Y sky130_fd_sc_hd__nand3_1
X_24569_ hold2664/X _26253_/Q _24587_/S vssd1 vssd1 vccd1 vccd1 _24569_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17110_ _17108_/X _23187_/B _17109_/X vssd1 vssd1 vccd1 vccd1 _17111_/A sky130_fd_sc_hd__a21o_1
X_14322_ _14322_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14322_/Y sky130_fd_sc_hd__nand2_1
X_18090_ _19359_/A vssd1 vssd1 vccd1 vccd1 _21869_/B sky130_fd_sc_hd__inv_2
X_26308_ _26308_/CLK _26308_/D vssd1 vssd1 vccd1 vccd1 _26308_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17041_ _20163_/B _25881_/Q _25817_/Q vssd1 vssd1 vccd1 vccd1 _17042_/B sky130_fd_sc_hd__mux2_2
X_26239_ _26239_/CLK _26239_/D vssd1 vssd1 vccd1 vccd1 _26239_/Q sky130_fd_sc_hd__dfxtp_2
X_14253_ hold651/X _14252_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold652/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13204_ _26170_/Q _13065_/X _13203_/X vssd1 vssd1 vccd1 vccd1 _13204_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14184_ _18694_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14184_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13135_ _26287_/Q _25656_/Q vssd1 vssd1 vccd1 vccd1 _14521_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18992_ _18992_/A _19126_/B vssd1 vssd1 vccd1 vccd1 _18992_/Y sky130_fd_sc_hd__nand2_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ _18528_/A _25723_/Q vssd1 vssd1 vccd1 vccd1 _17945_/A sky130_fd_sc_hd__nand2_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _26274_/Q _25643_/Q vssd1 vssd1 vccd1 vccd1 _14482_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_178_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17874_ _17874_/A _17874_/B vssd1 vssd1 vccd1 vccd1 _17875_/A sky130_fd_sc_hd__or2_1
X_19613_ _26248_/Q hold401/X vssd1 vssd1 vccd1 vccd1 _19613_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16825_ _16823_/X _16711_/X _16824_/Y _25878_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16826_/A sky130_fd_sc_hd__a32o_1
X_19544_ _19543_/Y _19272_/X _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19545_/B
+ sky130_fd_sc_hd__a211o_1
X_16756_ _16756_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16756_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13968_ _14000_/A hold638/X vssd1 vssd1 vccd1 vccd1 hold639/A sky130_fd_sc_hd__nand2_1
X_15707_ _23095_/B _15707_/B vssd1 vssd1 vccd1 vccd1 _23092_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12919_ _12840_/X _12916_/X _12917_/X _12918_/X vssd1 vssd1 vccd1 vccd1 _12919_/X
+ sky130_fd_sc_hd__o211a_1
X_19475_ _21101_/A _19473_/Y _21105_/C vssd1 vssd1 vccd1 vccd1 _19565_/B sky130_fd_sc_hd__o21a_1
X_16687_ _16698_/A hold608/X vssd1 vssd1 vccd1 vccd1 hold609/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13899_ hold558/X _13898_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold559/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18426_ _18446_/A _25747_/Q _21716_/A vssd1 vssd1 vccd1 vccd1 _18427_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_174_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15638_ _16561_/A _16711_/A vssd1 vssd1 vccd1 vccd1 _16911_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18357_ _18355_/Y _18356_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25662_/D sky130_fd_sc_hd__a21oi_1
X_15569_ _16510_/A _16711_/A vssd1 vssd1 vccd1 vccd1 _16883_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17308_ _17513_/A _17308_/B vssd1 vssd1 vccd1 vccd1 _17308_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_72_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18288_ _18288_/A _18288_/B _18288_/C vssd1 vssd1 vccd1 vccd1 _21812_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_126_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17239_ _17478_/A _17239_/B vssd1 vssd1 vccd1 vccd1 _17239_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_47_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold902 hold902/A vssd1 vssd1 vccd1 vccd1 hold902/X sky130_fd_sc_hd__buf_1
Xhold913 hold913/A vssd1 vssd1 vccd1 vccd1 hold913/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20250_ _20250_/A _25844_/Q vssd1 vssd1 vccd1 vccd1 _20254_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold924 hold924/A vssd1 vssd1 vccd1 vccd1 hold924/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 hold935/A vssd1 vssd1 vccd1 vccd1 hold935/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 hold946/A vssd1 vssd1 vccd1 vccd1 hold946/X sky130_fd_sc_hd__buf_1
XFILLER_0_101_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold957 hold957/A vssd1 vssd1 vccd1 vccd1 hold957/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 hold968/A vssd1 vssd1 vccd1 vccd1 hold968/X sky130_fd_sc_hd__dlygate4sd3_1
X_20181_ _20181_/A _20181_/B vssd1 vssd1 vccd1 vccd1 _21059_/C sky130_fd_sc_hd__nand2_4
Xhold979 hold979/A vssd1 vssd1 vccd1 vccd1 hold979/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2303 _24169_/X vssd1 vssd1 vccd1 vccd1 _24170_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2314 _26012_/Q vssd1 vssd1 vccd1 vccd1 hold2314/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2325 _26189_/Q vssd1 vssd1 vccd1 vccd1 hold2325/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23940_ _23940_/A vssd1 vssd1 vccd1 vccd1 _26048_/D sky130_fd_sc_hd__clkbuf_1
Xhold2336 _26113_/Q vssd1 vssd1 vccd1 vccd1 hold2336/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2347 _25426_/Q vssd1 vssd1 vccd1 vccd1 _15013_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1602 _25610_/Q vssd1 vssd1 vccd1 vccd1 _17386_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2358 _23968_/X vssd1 vssd1 vccd1 vccd1 _23969_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1613 _21640_/Y vssd1 vssd1 vccd1 vccd1 _25832_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2369 _24976_/Q vssd1 vssd1 vccd1 vccd1 _12613_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1624 _25783_/Q vssd1 vssd1 vccd1 vccd1 _20387_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1635 _25836_/Q vssd1 vssd1 vccd1 vccd1 _21703_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1646 _17429_/Y vssd1 vssd1 vccd1 vccd1 _25614_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23871_ _26027_/Q hold2130/X _23907_/S vssd1 vssd1 vccd1 vccd1 _23871_/X sky130_fd_sc_hd__mux2_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1657 _25606_/Q vssd1 vssd1 vccd1 vccd1 _17346_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1668 _21182_/Y vssd1 vssd1 vccd1 vccd1 _25807_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1679 _25879_/Q vssd1 vssd1 vccd1 vccd1 _22838_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_25610_ _26116_/CLK _25610_/D vssd1 vssd1 vccd1 vccd1 _25610_/Q sky130_fd_sc_hd__dfxtp_2
X_22822_ _22820_/X _22821_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22822_/Y sky130_fd_sc_hd__a21oi_1
X_25541_ _26047_/CLK _25541_/D vssd1 vssd1 vccd1 vccd1 _25541_/Q sky130_fd_sc_hd__dfxtp_1
X_22753_ _16799_/B _22421_/X _22747_/X _22748_/Y _22752_/X vssd1 vssd1 vccd1 vccd1
+ _22754_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_17_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21704_ _21702_/Y _21703_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21704_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25472_ _25472_/CLK _25472_/D vssd1 vssd1 vccd1 vccd1 _25472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22684_ _22683_/A _22454_/X _22683_/B vssd1 vssd1 vccd1 vccd1 _22685_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_137_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24423_ _24423_/A vssd1 vssd1 vccd1 vccd1 _26205_/D sky130_fd_sc_hd__clkbuf_1
X_21635_ _21634_/Y _21203_/X _20986_/A _20957_/A vssd1 vssd1 vccd1 vccd1 _21635_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_164_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24354_ _24354_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24355_/A sky130_fd_sc_hd__and2_1
XFILLER_0_118_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21566_ _21566_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21571_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23305_ _23305_/A vssd1 vssd1 vccd1 vccd1 _23310_/B sky130_fd_sc_hd__inv_2
XFILLER_0_145_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20517_ _20517_/A _22436_/B vssd1 vssd1 vccd1 vccd1 _20518_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24285_ _24285_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24286_/A sky130_fd_sc_hd__and2_1
XFILLER_0_133_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21497_ _21497_/A _21497_/B _21497_/C vssd1 vssd1 vccd1 vccd1 _21501_/A sky130_fd_sc_hd__nand3_1
X_26024_ _26042_/CLK _26024_/D vssd1 vssd1 vccd1 vccd1 _26024_/Q sky130_fd_sc_hd__dfxtp_1
X_23236_ _23236_/A vssd1 vssd1 vccd1 vccd1 _24949_/S sky130_fd_sc_hd__buf_12
XFILLER_0_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20448_ _20448_/A _20448_/B vssd1 vssd1 vccd1 vccd1 _21547_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_132_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23167_ _23167_/A _23167_/B vssd1 vssd1 vccd1 vccd1 _23169_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20379_ _20379_/A _20379_/B vssd1 vssd1 vccd1 vccd1 _20380_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22118_ _22118_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _22118_/X sky130_fd_sc_hd__and2_1
XFILLER_0_24_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23098_ _16940_/B _22421_/A _23092_/X _23093_/Y _23097_/X vssd1 vssd1 vccd1 vccd1
+ _23099_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_101_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14940_ _14948_/A _14932_/A _14932_/B vssd1 vssd1 vccd1 vccd1 _14942_/A sky130_fd_sc_hd__a21bo_1
X_22049_ _22550_/A _22758_/B vssd1 vssd1 vccd1 vccd1 _22055_/C sky130_fd_sc_hd__nand2_1
X_14871_ _25857_/Q _13466_/A _14870_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14872_/A
+ sky130_fd_sc_hd__a22o_1
X_16610_ _16610_/A _16610_/B vssd1 vssd1 vccd1 vccd1 _16620_/A sky130_fd_sc_hd__or2_1
XFILLER_0_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25808_ _25808_/CLK _25808_/D vssd1 vssd1 vccd1 vccd1 _25808_/Q sky130_fd_sc_hd__dfxtp_2
X_13822_ _26269_/Q _13801_/X _13793_/X _13821_/Y vssd1 vssd1 vccd1 vccd1 _13823_/B
+ sky130_fd_sc_hd__a22o_1
X_17590_ _17590_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _17590_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16541_ _16541_/A _16541_/B vssd1 vssd1 vccd1 vccd1 _16542_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_173_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13753_ hold525/X _13752_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold526/A sky130_fd_sc_hd__a21oi_1
X_25739_ _25808_/CLK _25739_/D vssd1 vssd1 vccd1 vccd1 _25739_/Q sky130_fd_sc_hd__dfxtp_1
X_12704_ _12704_/A hold997/X hold837/X vssd1 vssd1 vccd1 vccd1 _12707_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_85_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19260_ _19280_/B _19350_/B vssd1 vssd1 vccd1 vccd1 _19261_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16472_ _16468_/B _16468_/A _16486_/B _16471_/Y vssd1 vssd1 vccd1 vccd1 _16472_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13684_ _26247_/Q _13612_/X _13605_/X _13683_/Y vssd1 vssd1 vccd1 vccd1 _13685_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18211_ _18211_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18211_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_54_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15423_ _16401_/A _15778_/B vssd1 vssd1 vccd1 vccd1 _16831_/A sky130_fd_sc_hd__nand2_1
X_12635_ _12635_/A _12635_/B vssd1 vssd1 vccd1 vccd1 _12635_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19191_ _19989_/A _19191_/B vssd1 vssd1 vccd1 vccd1 _19191_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15354_ _16346_/A _16711_/A vssd1 vssd1 vccd1 vccd1 _16803_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18142_ _18372_/A _18514_/A vssd1 vssd1 vccd1 vccd1 _18143_/B sky130_fd_sc_hd__xnor2_1
X_12566_ _12566_/A vssd1 vssd1 vccd1 vccd1 _24966_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14305_ _14344_/A hold11/X vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15285_ _22683_/B _15285_/B vssd1 vssd1 vccd1 vccd1 _22679_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_123_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18073_ _18073_/A _18073_/B vssd1 vssd1 vccd1 vccd1 _18075_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12497_ _14345_/A _23199_/C vssd1 vssd1 vccd1 vccd1 _12497_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14236_ _14236_/A hold632/X vssd1 vssd1 vccd1 vccd1 hold633/A sky130_fd_sc_hd__nand2_1
Xhold209 hold209/A vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
X_17024_ _25624_/Q vssd1 vssd1 vccd1 vccd1 _20132_/B sky130_fd_sc_hd__inv_2
XFILLER_0_106_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14167_ _14180_/A _14167_/B vssd1 vssd1 vccd1 vccd1 _14167_/Y sky130_fd_sc_hd__nand2_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _18107_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13118_/X sky130_fd_sc_hd__or2_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _14180_/A _14098_/B vssd1 vssd1 vccd1 vccd1 _14098_/Y sky130_fd_sc_hd__nand2_1
X_18975_ _19025_/A _18975_/B vssd1 vssd1 vccd1 vccd1 _18975_/X sky130_fd_sc_hd__xor2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ _17927_/B _17927_/A vssd1 vssd1 vccd1 vccd1 _17928_/A sky130_fd_sc_hd__or2_1
X_13049_ _13220_/A vssd1 vssd1 vccd1 vccd1 _13049_/X sky130_fd_sc_hd__buf_12
XFILLER_0_147_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17857_ _18611_/A _25721_/Q vssd1 vssd1 vccd1 vccd1 _17859_/A sky130_fd_sc_hd__nand2_1
X_16808_ _16935_/A _16813_/B vssd1 vssd1 vccd1 vccd1 _16810_/B sky130_fd_sc_hd__nand2_1
X_17788_ _18153_/C vssd1 vssd1 vccd1 vccd1 _17789_/B sky130_fd_sc_hd__inv_2
XFILLER_0_89_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19527_ _19525_/Y _19526_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19527_/Y sky130_fd_sc_hd__a21oi_1
X_16739_ _16740_/B _16740_/A vssd1 vssd1 vccd1 vccd1 _16739_/X sky130_fd_sc_hd__or2_1
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19458_ _19458_/A _21075_/B vssd1 vssd1 vccd1 vccd1 _19458_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_158_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18409_ _18409_/A _18409_/B _18409_/C vssd1 vssd1 vccd1 vccd1 _22017_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_9_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19389_ _20935_/A _21938_/B _25607_/Q vssd1 vssd1 vccd1 vccd1 _20940_/C sky130_fd_sc_hd__nand3_1
X_21420_ _21420_/A _21420_/B vssd1 vssd1 vccd1 vccd1 _21421_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21351_ _21351_/A _21351_/B _21351_/C vssd1 vssd1 vccd1 vccd1 _21355_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20302_ _26284_/Q hold736/X vssd1 vssd1 vccd1 vccd1 _20302_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24070_ _24070_/A vssd1 vssd1 vccd1 vccd1 _26090_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold710 hold710/A vssd1 vssd1 vccd1 vccd1 hold710/X sky130_fd_sc_hd__dlygate4sd3_1
X_21282_ _26314_/Q _21228_/X hold794/X vssd1 vssd1 vccd1 vccd1 _21285_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_188_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold721 hold721/A vssd1 vssd1 vccd1 vccd1 hold721/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold732 hold732/A vssd1 vssd1 vccd1 vccd1 hold732/X sky130_fd_sc_hd__dlygate4sd3_1
X_23021_ _23197_/A _23021_/B vssd1 vssd1 vccd1 vccd1 _23021_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_13_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold743 hold743/A vssd1 vssd1 vccd1 vccd1 hold743/X sky130_fd_sc_hd__dlygate4sd3_1
X_20233_ _20660_/A _20233_/B vssd1 vssd1 vccd1 vccd1 _20233_/Y sky130_fd_sc_hd__nand2_1
Xhold754 hold754/A vssd1 vssd1 vccd1 vccd1 hold754/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold765 hold765/A vssd1 vssd1 vccd1 vccd1 hold765/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold776 hold776/A vssd1 vssd1 vccd1 vccd1 hold776/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 hold787/A vssd1 vssd1 vccd1 vccd1 hold787/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold798 hold798/A vssd1 vssd1 vccd1 vccd1 hold798/X sky130_fd_sc_hd__dlygate4sd3_1
X_20164_ _20167_/A _20167_/C vssd1 vssd1 vccd1 vccd1 _20165_/A sky130_fd_sc_hd__nand2_1
Xhold2100 _23367_/X vssd1 vssd1 vccd1 vccd1 _23368_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2111 _25970_/Q vssd1 vssd1 vccd1 vccd1 hold2111/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2122 _25991_/Q vssd1 vssd1 vccd1 vccd1 _14788_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2133 _25956_/Q vssd1 vssd1 vccd1 vccd1 hold2133/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24972_ _24983_/CLK _24972_/D vssd1 vssd1 vccd1 vccd1 _24972_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2144 _25662_/Q vssd1 vssd1 vccd1 vccd1 _13170_/A sky130_fd_sc_hd__dlygate4sd3_1
X_20095_ _20094_/B _20095_/B _20095_/C vssd1 vssd1 vccd1 vccd1 _20096_/B sky130_fd_sc_hd__nand3b_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1410 _16784_/Y vssd1 vssd1 vccd1 vccd1 _25551_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2155 _25988_/Q vssd1 vssd1 vccd1 vccd1 _14761_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1421 _25019_/Q vssd1 vssd1 vccd1 vccd1 _17256_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2166 _26161_/Q vssd1 vssd1 vccd1 vccd1 hold2166/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2177 _26031_/Q vssd1 vssd1 vccd1 vccd1 hold2177/X sky130_fd_sc_hd__dlygate4sd3_1
X_23923_ _23923_/A _23923_/B vssd1 vssd1 vccd1 vccd1 _23924_/C sky130_fd_sc_hd__nand2_1
Xhold1432 _19654_/Y vssd1 vssd1 vccd1 vccd1 _25747_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2188 _25952_/Q vssd1 vssd1 vccd1 vccd1 hold2188/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1443 _25570_/Q vssd1 vssd1 vccd1 vccd1 _16914_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2199 _25995_/Q vssd1 vssd1 vccd1 vccd1 _14824_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1454 _19905_/Y vssd1 vssd1 vccd1 vccd1 _25765_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1465 _25051_/Q vssd1 vssd1 vccd1 vccd1 _17550_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23854_ _23854_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23855_/A sky130_fd_sc_hd__and2_1
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1476 _20963_/Y vssd1 vssd1 vccd1 vccd1 _25799_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1487 _25097_/Q vssd1 vssd1 vccd1 vccd1 _18658_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1498 _21413_/Y vssd1 vssd1 vccd1 vccd1 _25818_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22805_ _22937_/A _22805_/B vssd1 vssd1 vccd1 vccd1 _22805_/Y sky130_fd_sc_hd__nand2_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23785_ _14859_/B _26000_/Q _23831_/S vssd1 vssd1 vccd1 vccd1 _23785_/X sky130_fd_sc_hd__mux2_1
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20997_ _22536_/B vssd1 vssd1 vccd1 vccd1 _22011_/B sky130_fd_sc_hd__inv_2
XFILLER_0_79_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25524_ _25533_/CLK hold747/X vssd1 vssd1 vccd1 vccd1 hold745/A sky130_fd_sc_hd__dfxtp_1
X_22736_ _22736_/A _23001_/B _22736_/C vssd1 vssd1 vccd1 vccd1 _22736_/X sky130_fd_sc_hd__and3_1
X_25455_ _25535_/CLK _25455_/D vssd1 vssd1 vccd1 vccd1 _25455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22667_ _22667_/A _22667_/B vssd1 vssd1 vccd1 vccd1 _22667_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24406_ hold2353/X hold2321/X _24433_/S vssd1 vssd1 vccd1 vccd1 _24407_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_180_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21618_ _26334_/Q hold566/X vssd1 vssd1 vccd1 vccd1 _21618_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_118_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25386_ _26336_/CLK hold148/X vssd1 vssd1 vccd1 vccd1 hold146/A sky130_fd_sc_hd__dfxtp_1
X_22598_ _23103_/B _22958_/B vssd1 vssd1 vccd1 vccd1 _22600_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_7__f_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _25472_/CLK sky130_fd_sc_hd__clkbuf_16
X_24337_ _24337_/A vssd1 vssd1 vccd1 vccd1 _26177_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21549_ _21549_/A _21549_/B vssd1 vssd1 vccd1 vccd1 _21550_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_161_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15070_ _15050_/B _15067_/B _15067_/X _15052_/X _15059_/B vssd1 vssd1 vccd1 vccd1
+ _15110_/A sky130_fd_sc_hd__o221ai_4
XFILLER_0_161_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24268_ _24268_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24269_/A sky130_fd_sc_hd__and2_1
XFILLER_0_132_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26007_ _26009_/CLK _26007_/D vssd1 vssd1 vccd1 vccd1 _26007_/Q sky130_fd_sc_hd__dfxtp_1
X_14021_ _25798_/Q vssd1 vssd1 vccd1 vccd1 _18139_/B sky130_fd_sc_hd__inv_2
X_23219_ _23278_/B _24956_/S vssd1 vssd1 vccd1 vccd1 _23227_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24199_ _24199_/A vssd1 vssd1 vccd1 vccd1 _26132_/D sky130_fd_sc_hd__clkbuf_1
X_18760_ _18758_/X _18269_/X _18759_/X vssd1 vssd1 vccd1 vccd1 _18761_/A sky130_fd_sc_hd__a21o_1
X_15972_ _15987_/B _15972_/B vssd1 vssd1 vccd1 vccd1 _15999_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_175_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17711_ _17711_/A _23201_/B vssd1 vssd1 vccd1 vccd1 _17721_/A sky130_fd_sc_hd__nand2_1
X_14923_ _14923_/A _14923_/B vssd1 vssd1 vccd1 vccd1 _14923_/Y sky130_fd_sc_hd__nand2_1
X_18691_ _18691_/A _25824_/Q _18691_/C vssd1 vssd1 vccd1 vccd1 _20447_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_211_clk _26093_/CLK vssd1 vssd1 vccd1 vccd1 _26089_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
X_17642_ _18252_/A _17642_/B vssd1 vssd1 vccd1 vccd1 _17642_/Y sky130_fd_sc_hd__nand2_1
X_14854_ _14854_/A vssd1 vssd1 vccd1 vccd1 _15042_/A sky130_fd_sc_hd__inv_2
XFILLER_0_37_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13805_ _13823_/A _13805_/B vssd1 vssd1 vccd1 vccd1 _13805_/Y sky130_fd_sc_hd__nand2_1
X_17573_ _17571_/X _17528_/X _17572_/X vssd1 vssd1 vccd1 vccd1 _17574_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_98_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14785_ _14785_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14785_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_98_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19312_ _19310_/Y _19311_/Y _19086_/X vssd1 vssd1 vccd1 vccd1 _19312_/Y sky130_fd_sc_hd__a21oi_1
X_16524_ _16524_/A _16524_/B vssd1 vssd1 vccd1 vccd1 _16543_/B sky130_fd_sc_hd__nor2_1
X_13736_ _13760_/A hold365/X vssd1 vssd1 vccd1 vccd1 hold366/A sky130_fd_sc_hd__nand2_1
XFILLER_0_129_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19243_ _19241_/Y hold923/X _19086_/X vssd1 vssd1 vccd1 vccd1 hold924/A sky130_fd_sc_hd__a21oi_1
X_16455_ _16456_/B _16456_/A vssd1 vssd1 vccd1 vccd1 _16455_/X sky130_fd_sc_hd__or2_1
X_13667_ hold675/X _13666_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold676/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15406_ _15406_/A _15406_/B _15406_/C vssd1 vssd1 vccd1 vccd1 _15408_/B sky130_fd_sc_hd__and3_1
XFILLER_0_155_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12618_ _12618_/A _12618_/B vssd1 vssd1 vccd1 vccd1 _12619_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19174_ _26217_/Q _19134_/X hold766/X vssd1 vssd1 vccd1 vccd1 _19175_/C sky130_fd_sc_hd__a21o_1
X_16386_ hold518/X vssd1 vssd1 vccd1 vccd1 _16390_/B sky130_fd_sc_hd__inv_2
X_13598_ _13642_/A hold563/X vssd1 vssd1 vccd1 vccd1 hold564/A sky130_fd_sc_hd__nand2_1
XFILLER_0_54_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18125_ _18125_/A _18125_/B _25781_/Q vssd1 vssd1 vccd1 vccd1 _20290_/B sky130_fd_sc_hd__nand3_2
X_15337_ _15621_/A _16329_/B vssd1 vssd1 vccd1 vccd1 _15340_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12549_ _17707_/B _12546_/X _17742_/A vssd1 vssd1 vccd1 vccd1 _12549_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_124_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18056_ _19073_/A _18474_/A vssd1 vssd1 vccd1 vccd1 _18057_/B sky130_fd_sc_hd__xnor2_4
XANTENNA_1 _21007_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15268_ _15268_/A _15268_/B _15268_/C vssd1 vssd1 vccd1 vccd1 _15272_/B sky130_fd_sc_hd__and3_1
XFILLER_0_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17007_ _16993_/X _23187_/B _17006_/X vssd1 vssd1 vccd1 vccd1 _17012_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_50_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14219_ _25830_/Q vssd1 vssd1 vccd1 vccd1 _18814_/B sky130_fd_sc_hd__inv_2
XFILLER_0_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15199_ _15199_/A _15199_/B vssd1 vssd1 vccd1 vccd1 _15268_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_111_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18958_ _18958_/A _20087_/A vssd1 vssd1 vccd1 vccd1 _19080_/B sky130_fd_sc_hd__xor2_4
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17909_ _17909_/A _17909_/B _17909_/C vssd1 vssd1 vccd1 vccd1 _21731_/A sky130_fd_sc_hd__nand3_2
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18889_ _25898_/Q _22639_/A vssd1 vssd1 vccd1 vccd1 _18897_/A sky130_fd_sc_hd__or2_2
XFILLER_0_154_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_202_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _26231_/CLK sky130_fd_sc_hd__clkbuf_16
X_20920_ _21708_/A _21483_/B vssd1 vssd1 vccd1 vccd1 _20921_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20851_ _20851_/A _20851_/B vssd1 vssd1 vccd1 vccd1 _20852_/A sky130_fd_sc_hd__nand2_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23570_ _24922_/S hold347/A _23569_/X vssd1 vssd1 vccd1 vccd1 _23570_/Y sky130_fd_sc_hd__o21ai_1
X_20782_ _20782_/A _25858_/Q vssd1 vssd1 vccd1 vccd1 _20787_/B sky130_fd_sc_hd__nand2_1
X_22521_ _22906_/B _23055_/B vssd1 vssd1 vccd1 vccd1 _22523_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25240_ _25817_/CLK hold649/X vssd1 vssd1 vccd1 vccd1 hold647/A sky130_fd_sc_hd__dfxtp_1
X_22452_ _23191_/C vssd1 vssd1 vccd1 vccd1 _22999_/C sky130_fd_sc_hd__buf_8
XFILLER_0_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21403_ _21403_/A _21403_/B _21403_/C vssd1 vssd1 vccd1 vccd1 _21404_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_162_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25171_ _25752_/CLK hold517/X vssd1 vssd1 vccd1 vccd1 hold515/A sky130_fd_sc_hd__dfxtp_1
X_22383_ _22368_/X _22382_/Y _17229_/B vssd1 vssd1 vccd1 vccd1 _22383_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24122_ _24122_/A vssd1 vssd1 vccd1 vccd1 _26107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21334_ _21385_/A _21691_/C vssd1 vssd1 vccd1 vccd1 _21335_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_170_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24053_ input5/X hold2277/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24054_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21265_ _21265_/A _21265_/B vssd1 vssd1 vccd1 vccd1 _21268_/B sky130_fd_sc_hd__nand2_1
Xhold540 hold540/A vssd1 vssd1 vccd1 vccd1 hold540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 hold551/A vssd1 vssd1 vccd1 vccd1 hold551/X sky130_fd_sc_hd__dlygate4sd3_1
X_23004_ _22995_/Y _23003_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _23004_/X sky130_fd_sc_hd__a21o_1
Xhold562 hold562/A vssd1 vssd1 vccd1 vccd1 hold562/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20216_ _20216_/A _20216_/B vssd1 vssd1 vccd1 vccd1 _20218_/A sky130_fd_sc_hd__nand2_1
Xhold573 hold573/A vssd1 vssd1 vccd1 vccd1 hold573/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold584 hold584/A vssd1 vssd1 vccd1 vccd1 hold584/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 hold595/A vssd1 vssd1 vccd1 vccd1 hold595/X sky130_fd_sc_hd__dlygate4sd3_1
X_21196_ _21646_/B _21597_/B vssd1 vssd1 vccd1 vccd1 _21198_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_15__f_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_99_clk/A
+ sky130_fd_sc_hd__clkbuf_16
X_20147_ _21033_/C vssd1 vssd1 vccd1 vccd1 _21036_/B sky130_fd_sc_hd__inv_2
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24955_ _16655_/A _16667_/B _24956_/S vssd1 vssd1 vccd1 vccd1 _24955_/X sky130_fd_sc_hd__mux2_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20078_ _21228_/A vssd1 vssd1 vccd1 vccd1 _20078_/X sky130_fd_sc_hd__buf_8
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1240 _25761_/Q vssd1 vssd1 vccd1 vccd1 _19852_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1251 _13288_/X vssd1 vssd1 vccd1 vccd1 _25100_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23906_ _23906_/A vssd1 vssd1 vccd1 vccd1 _26039_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1262 _25757_/Q vssd1 vssd1 vccd1 vccd1 _19796_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1273 _13364_/X vssd1 vssd1 vccd1 vccd1 _25112_/D sky130_fd_sc_hd__dlygate4sd3_1
X_24886_ _16049_/B _16069_/B _24922_/S vssd1 vssd1 vccd1 vccd1 _24887_/A sky130_fd_sc_hd__mux2_1
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1284 _25724_/Q vssd1 vssd1 vccd1 vccd1 _19325_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1295 _16866_/Y vssd1 vssd1 vccd1 vccd1 _25563_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23837_ _23837_/A vssd1 vssd1 vccd1 vccd1 _26016_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14570_ _14585_/A hold119/X vssd1 vssd1 vccd1 vccd1 hold120/A sky130_fd_sc_hd__nand2_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23768_ _23768_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23769_/A sky130_fd_sc_hd__and2_1
XFILLER_0_67_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25507_ _25510_/CLK _25507_/D vssd1 vssd1 vccd1 vccd1 hold999/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13521_ _13516_/Y _13520_/Y _12558_/B vssd1 vssd1 vccd1 vccd1 hold844/A sky130_fd_sc_hd__a21oi_1
X_22719_ _18958_/A _25837_/Q _22717_/Y _22718_/Y vssd1 vssd1 vccd1 vccd1 _22720_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23699_ hold2072/X _25972_/Q _23754_/S vssd1 vssd1 vccd1 vccd1 _23699_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16240_ _16240_/A _16245_/A vssd1 vssd1 vccd1 vccd1 _16240_/Y sky130_fd_sc_hd__nand2_1
X_13452_ _13522_/A _13450_/X _23629_/B _13451_/X vssd1 vssd1 vccd1 vccd1 _13452_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25438_ _26047_/CLK _25438_/D vssd1 vssd1 vccd1 vccd1 _25438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16171_ _16171_/A _16171_/B vssd1 vssd1 vccd1 vccd1 _16216_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_152_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13383_ _13383_/A vssd1 vssd1 vccd1 vccd1 _19744_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25369_ _26193_/CLK hold262/X vssd1 vssd1 vccd1 vccd1 hold260/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15122_ _15122_/A vssd1 vssd1 vccd1 vccd1 _16712_/A sky130_fd_sc_hd__inv_2
XFILLER_0_51_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15053_ _15270_/A _15068_/B _15052_/X vssd1 vssd1 vccd1 vccd1 _15055_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_120_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19930_ _19923_/X _19929_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19930_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_160_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14004_ _26298_/Q _13988_/X _13981_/X _14003_/Y vssd1 vssd1 vccd1 vccd1 _14005_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19861_ _19862_/B _19862_/A vssd1 vssd1 vccd1 vccd1 _19861_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18812_ _18954_/A _25766_/Q vssd1 vssd1 vccd1 vccd1 _18814_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19792_ _19793_/B _19793_/A vssd1 vssd1 vccd1 vccd1 _19792_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18743_ _18741_/Y _18742_/Y _18539_/X vssd1 vssd1 vccd1 vccd1 _25681_/D sky130_fd_sc_hd__a21oi_1
X_15955_ _15953_/B _16000_/B _15954_/Y vssd1 vssd1 vccd1 vccd1 _15955_/X sky130_fd_sc_hd__a21o_1
X_14906_ _14906_/A vssd1 vssd1 vccd1 vccd1 _25412_/D sky130_fd_sc_hd__inv_2
X_18674_ _18674_/A _18674_/B _18674_/C vssd1 vssd1 vccd1 vccd1 _22372_/A sky130_fd_sc_hd__nand3_1
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15886_ _15956_/A hold461/X vssd1 vssd1 vccd1 vccd1 hold462/A sky130_fd_sc_hd__nand2_1
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17625_ _17623_/X _17528_/X _17624_/X vssd1 vssd1 vccd1 vccd1 _17626_/A sky130_fd_sc_hd__a21o_1
X_14837_ _25853_/Q _12527_/A _14836_/Y _14696_/Y vssd1 vssd1 vccd1 vccd1 _14837_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17556_ _17556_/A _17556_/B vssd1 vssd1 vccd1 vccd1 _17556_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_59_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14768_ _14900_/A _14768_/B vssd1 vssd1 vccd1 vccd1 _14768_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16507_ _16505_/X hold746/X _16343_/X vssd1 vssd1 vccd1 vccd1 hold747/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_175_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13719_ _25750_/Q vssd1 vssd1 vccd1 vccd1 _18489_/B sky130_fd_sc_hd__inv_2
XFILLER_0_156_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17487_ _17485_/X _17241_/X _17486_/X vssd1 vssd1 vccd1 vccd1 _17488_/A sky130_fd_sc_hd__a21o_1
X_14699_ _14696_/Y _15621_/A _16702_/A vssd1 vssd1 vccd1 vccd1 _14899_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_156_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19226_ _19220_/X _18879_/X _19225_/X vssd1 vssd1 vccd1 vccd1 _19227_/A sky130_fd_sc_hd__a21o_1
X_16438_ _16438_/A _16438_/B vssd1 vssd1 vccd1 vccd1 _16461_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_117_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19157_ _19157_/A _19980_/B _19157_/C vssd1 vssd1 vccd1 vccd1 _19157_/X sky130_fd_sc_hd__and3_1
X_16369_ _22796_/B _16369_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _16371_/A sky130_fd_sc_hd__and3_1
XFILLER_0_14_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18108_ _18106_/X _17528_/X _18107_/X vssd1 vssd1 vccd1 vccd1 _18109_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19088_ _21749_/A _20023_/B vssd1 vssd1 vccd1 vccd1 _19088_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18039_ _21835_/B _25604_/Q vssd1 vssd1 vccd1 vccd1 _18041_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21050_ _21050_/A _25867_/Q vssd1 vssd1 vccd1 vccd1 _21054_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20001_ _20004_/A _20004_/C vssd1 vssd1 vccd1 vccd1 _20003_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21952_ _21952_/A _22715_/B vssd1 vssd1 vccd1 vccd1 _21953_/B sky130_fd_sc_hd__nand2_1
X_24740_ hold2648/X hold2625/X _24740_/S vssd1 vssd1 vccd1 vccd1 _24741_/A sky130_fd_sc_hd__mux2_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20903_ _21042_/A _20903_/B _20902_/X vssd1 vssd1 vccd1 vccd1 _20904_/B sky130_fd_sc_hd__or3b_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24671_ hold2652/X hold2591/X _24740_/S vssd1 vssd1 vccd1 vccd1 _24672_/A sky130_fd_sc_hd__mux2_1
X_21883_ _21883_/A _22662_/B vssd1 vssd1 vccd1 vccd1 _21884_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_68_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23622_ hold1991/X _25947_/Q _23677_/S vssd1 vssd1 vccd1 vccd1 _23622_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_49_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20834_ _20836_/B _20836_/C vssd1 vssd1 vccd1 vccd1 _20835_/A sky130_fd_sc_hd__nand2_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26341_ _26341_/CLK _26341_/D vssd1 vssd1 vccd1 vccd1 _26341_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23553_ _23550_/Y _23552_/Y _24946_/A vssd1 vssd1 vccd1 vccd1 _23553_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_147_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20765_ _21400_/C _21676_/B vssd1 vssd1 vccd1 vccd1 _20767_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_175_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22504_ _22504_/A _22504_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22506_/A sky130_fd_sc_hd__or3_1
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26272_ _26273_/CLK _26272_/D vssd1 vssd1 vccd1 vccd1 _26272_/Q sky130_fd_sc_hd__dfxtp_1
X_23484_ _23484_/A _23484_/B vssd1 vssd1 vccd1 vccd1 _23484_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_162_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20696_ _20696_/A _20696_/B vssd1 vssd1 vccd1 vccd1 _20697_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_162_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25223_ _25807_/CLK hold514/X vssd1 vssd1 vccd1 vccd1 hold512/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22435_ _22435_/A _25890_/Q vssd1 vssd1 vccd1 vccd1 _22435_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_18_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25154_ _26286_/CLK hold493/X vssd1 vssd1 vccd1 vccd1 hold491/A sky130_fd_sc_hd__dfxtp_1
X_22366_ _22366_/A _22387_/B vssd1 vssd1 vccd1 vccd1 _22366_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_116_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24105_ hold2124/X _26102_/Q _24126_/S vssd1 vssd1 vccd1 vccd1 _24105_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21317_ _21678_/B _21370_/A vssd1 vssd1 vccd1 vccd1 _21319_/A sky130_fd_sc_hd__nand2_1
X_25085_ _26299_/CLK _25085_/D vssd1 vssd1 vccd1 vccd1 _25085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22297_ _25820_/Q _22297_/B vssd1 vssd1 vccd1 vccd1 _22297_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_130_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24036_ _24036_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24037_/A sky130_fd_sc_hd__and2_1
Xhold370 hold370/A vssd1 vssd1 vccd1 vccd1 hold370/X sky130_fd_sc_hd__dlygate4sd3_1
X_21248_ _21627_/C _21675_/C vssd1 vssd1 vccd1 vccd1 _21249_/B sky130_fd_sc_hd__nand2_1
Xhold381 hold381/A vssd1 vssd1 vccd1 vccd1 hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 hold392/A vssd1 vssd1 vccd1 vccd1 hold392/X sky130_fd_sc_hd__dlygate4sd3_1
X_21179_ _21179_/A _21179_/B vssd1 vssd1 vccd1 vccd1 _21180_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25987_ _25991_/CLK _25987_/D vssd1 vssd1 vccd1 vccd1 _25987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15740_ _23124_/B _15812_/B vssd1 vssd1 vccd1 vccd1 _16638_/B sky130_fd_sc_hd__nand2_1
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24938_ _24946_/A _24935_/X _24958_/B _24937_/Y vssd1 vssd1 vccd1 vccd1 _24938_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _12891_/X _14413_/A _12909_/X _25621_/Q vssd1 vssd1 vccd1 vccd1 _12952_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_172_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1070 _12970_/X vssd1 vssd1 vccd1 vccd1 _25044_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1081 _25085_/Q vssd1 vssd1 vccd1 vccd1 _18415_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1092 _13108_/X vssd1 vssd1 vccd1 vccd1 _25070_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15671_ _16585_/A _15778_/B vssd1 vssd1 vccd1 vccd1 _16923_/A sky130_fd_sc_hd__nand2_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24869_ _24852_/X _24868_/X _25912_/Q vssd1 vssd1 vccd1 vccd1 _24870_/A sky130_fd_sc_hd__mux2_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _26111_/Q _12748_/X _12882_/X vssd1 vssd1 vccd1 vccd1 _12883_/X sky130_fd_sc_hd__a21o_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _21291_/B _25876_/Q _25812_/Q vssd1 vssd1 vccd1 vccd1 _17411_/B sky130_fd_sc_hd__mux2_2
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _14620_/Y hold234/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold235/A sky130_fd_sc_hd__a21oi_1
X_18390_ _18390_/A _21210_/A vssd1 vssd1 vccd1 vccd1 _18738_/A sky130_fd_sc_hd__xor2_4
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17341_ _17535_/A _17586_/A vssd1 vssd1 vccd1 vccd1 _17342_/B sky130_fd_sc_hd__xnor2_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14553_ _14551_/Y hold99/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold100/A sky130_fd_sc_hd__a21oi_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _13522_/A hold739/X vssd1 vssd1 vccd1 vccd1 hold740/A sky130_fd_sc_hd__nand2_1
XFILLER_0_83_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17272_ _17272_/A _17272_/B vssd1 vssd1 vccd1 vccd1 _17272_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_181_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14484_ _14482_/Y hold60/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__a21oi_1
X_19011_ _19060_/A _19011_/B vssd1 vssd1 vccd1 vccd1 _19011_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_82_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16223_ _16223_/A vssd1 vssd1 vccd1 vccd1 _16238_/B sky130_fd_sc_hd__inv_2
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13435_ _26207_/Q _13426_/X _13434_/X vssd1 vssd1 vccd1 vccd1 _13435_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_126_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16154_ _16212_/A hold861/X vssd1 vssd1 vccd1 vccd1 _16154_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13366_ _26324_/Q _19701_/A vssd1 vssd1 vccd1 vccd1 _14638_/A sky130_fd_sc_hd__xor2_1
X_15105_ _15103_/X _15104_/Y _15090_/X vssd1 vssd1 vccd1 vccd1 _15105_/Y sky130_fd_sc_hd__a21oi_1
X_16085_ _16071_/B _16084_/B _16070_/A vssd1 vssd1 vccd1 vccd1 _16107_/A sky130_fd_sc_hd__o21ai_1
X_13297_ _13220_/X _14605_/A _13242_/X _19546_/A vssd1 vssd1 vccd1 vccd1 _13297_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15036_ _15000_/X _15032_/A _15035_/X vssd1 vssd1 vccd1 vccd1 _15037_/B sky130_fd_sc_hd__a21oi_1
X_19913_ _19914_/B _19914_/A vssd1 vssd1 vccd1 vccd1 _19913_/X sky130_fd_sc_hd__or2_1
XFILLER_0_139_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19844_ _19844_/A _20712_/B vssd1 vssd1 vccd1 vccd1 _19844_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19775_ _20517_/A _22436_/B _25634_/Q vssd1 vssd1 vccd1 vccd1 _20522_/C sky130_fd_sc_hd__nand3_1
X_16987_ _20285_/B _25845_/Q _25781_/Q vssd1 vssd1 vccd1 vccd1 _16988_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_78_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18726_ _20518_/B _19774_/A vssd1 vssd1 vccd1 vccd1 _18727_/B sky130_fd_sc_hd__nand2_1
X_15938_ _15956_/A hold443/X vssd1 vssd1 vccd1 vccd1 hold444/A sky130_fd_sc_hd__nand2_1
XFILLER_0_155_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18657_ _18657_/A _18657_/B vssd1 vssd1 vccd1 vccd1 _18657_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_189_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15869_ _15869_/A _15869_/B vssd1 vssd1 vccd1 vccd1 _15895_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_149_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17608_ _17608_/A _17608_/B vssd1 vssd1 vccd1 vccd1 _17608_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_114_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18588_ _18793_/A _25755_/Q _18894_/C vssd1 vssd1 vccd1 vccd1 _18589_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_175_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17539_ _17605_/A _17539_/B vssd1 vssd1 vccd1 vccd1 _17539_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20550_ _25852_/Q vssd1 vssd1 vccd1 vccd1 _22195_/B sky130_fd_sc_hd__inv_2
XFILLER_0_184_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19209_ _19220_/A _19294_/B vssd1 vssd1 vccd1 vccd1 _19211_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_61_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20481_ _20481_/A _25889_/Q vssd1 vssd1 vccd1 vccd1 _20487_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22220_ _18037_/A _25789_/Q _22218_/Y _22219_/Y vssd1 vssd1 vccd1 vccd1 _22221_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22151_ _22151_/A _22151_/B vssd1 vssd1 vccd1 vccd1 _22151_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_100_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21102_ _21102_/A _21102_/B vssd1 vssd1 vccd1 vccd1 _21105_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22082_ _22082_/A _22082_/B vssd1 vssd1 vccd1 vccd1 _23058_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_11_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25910_ _26002_/CLK _25910_/D vssd1 vssd1 vccd1 vccd1 _25910_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_61_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21033_ _21033_/A _21033_/B _21033_/C vssd1 vssd1 vccd1 vccd1 _21037_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_10_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25841_ _25860_/CLK _25841_/D vssd1 vssd1 vccd1 vccd1 _25841_/Q sky130_fd_sc_hd__dfxtp_4
X_22984_ _22984_/A _23001_/B _22984_/C vssd1 vssd1 vccd1 vccd1 _22984_/X sky130_fd_sc_hd__and3_1
X_25772_ _26275_/CLK _25772_/D vssd1 vssd1 vccd1 vccd1 _25772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24723_ _24723_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24724_/A sky130_fd_sc_hd__and2_1
X_21935_ _21933_/X _14270_/A _21934_/Y _14759_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _21936_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_96_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21866_ _21864_/X _14270_/A _21865_/Y _14740_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _21867_/A sky130_fd_sc_hd__a32o_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24654_ _24654_/A vssd1 vssd1 vccd1 vccd1 _26280_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23605_ _23605_/A _23629_/B vssd1 vssd1 vccd1 vccd1 _23606_/A sky130_fd_sc_hd__and2_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20817_ _20817_/A _21801_/B vssd1 vssd1 vccd1 vccd1 _20818_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_148_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21797_ _21797_/A _22145_/B vssd1 vssd1 vccd1 vccd1 _21797_/Y sky130_fd_sc_hd__nand2_1
X_24585_ _24585_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24586_/A sky130_fd_sc_hd__and2_1
XFILLER_0_38_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26324_ _26324_/CLK _26324_/D vssd1 vssd1 vccd1 vccd1 _26324_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_147_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20748_ _20747_/B _20748_/B _20748_/C vssd1 vssd1 vccd1 vccd1 _20749_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_65_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23536_ _24942_/S hold368/A _23535_/X vssd1 vssd1 vccd1 vccd1 _23536_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_181_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23467_ _24956_/S hold224/A _23466_/X vssd1 vssd1 vccd1 vccd1 _23467_/Y sky130_fd_sc_hd__o21ai_1
X_26255_ _26267_/CLK _26255_/D vssd1 vssd1 vccd1 vccd1 _26255_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_163_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20679_ _20681_/B vssd1 vssd1 vccd1 vccd1 _20680_/B sky130_fd_sc_hd__inv_2
XFILLER_0_52_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ _13220_/A vssd1 vssd1 vccd1 vccd1 _13220_/X sky130_fd_sc_hd__buf_8
XFILLER_0_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22418_ _22418_/A _22418_/B vssd1 vssd1 vccd1 vccd1 _22419_/B sky130_fd_sc_hd__nand2_1
X_25206_ _26289_/CLK hold744/X vssd1 vssd1 vccd1 vccd1 hold742/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23398_ hold281/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23398_/X sky130_fd_sc_hd__or2b_1
X_26186_ _26190_/CLK _26186_/D vssd1 vssd1 vccd1 vccd1 _26186_/Q sky130_fd_sc_hd__dfxtp_1
X_13151_ _13109_/X _13149_/X _13096_/X _13150_/X vssd1 vssd1 vccd1 vccd1 _13151_/X
+ sky130_fd_sc_hd__o211a_1
X_22349_ _18655_/A _25822_/Q _22347_/Y _22348_/Y vssd1 vssd1 vccd1 vccd1 _22350_/B
+ sky130_fd_sc_hd__a31o_1
X_25137_ _26152_/CLK hold770/X vssd1 vssd1 vccd1 vccd1 hold768/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25068_ _26152_/CLK _25068_/D vssd1 vssd1 vccd1 vccd1 _25068_/Q sky130_fd_sc_hd__dfxtp_1
X_13082_ _13082_/A vssd1 vssd1 vccd1 vccd1 _21749_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16910_ _16911_/B _16911_/A vssd1 vssd1 vccd1 vccd1 _16910_/X sky130_fd_sc_hd__or2_1
X_24019_ _24019_/A vssd1 vssd1 vccd1 vccd1 _26074_/D sky130_fd_sc_hd__clkbuf_1
X_17890_ _18611_/A _17895_/B vssd1 vssd1 vccd1 vccd1 _17893_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16841_ _25881_/Q _13468_/X _16774_/Y vssd1 vssd1 vccd1 vccd1 _16841_/Y sky130_fd_sc_hd__a21oi_1
X_19560_ _19560_/A _21265_/B vssd1 vssd1 vccd1 vccd1 _19560_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_176_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16772_ _16770_/Y _16771_/Y _16594_/X vssd1 vssd1 vccd1 vccd1 _16772_/Y sky130_fd_sc_hd__a21oi_1
X_13984_ _26295_/Q _13801_/X _13981_/X _13983_/Y vssd1 vssd1 vccd1 vccd1 _13985_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18511_ _20106_/C _22151_/A vssd1 vssd1 vccd1 vccd1 _20098_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_137_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15723_ _15723_/A _15810_/B vssd1 vssd1 vccd1 vccd1 _15724_/B sky130_fd_sc_hd__nand2_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ _12930_/X _12933_/X _12917_/X _12934_/X vssd1 vssd1 vccd1 vccd1 _12935_/X
+ sky130_fd_sc_hd__o211a_1
X_19491_ _19509_/B _19579_/B vssd1 vssd1 vccd1 vccd1 _19493_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ _21291_/B _19574_/A vssd1 vssd1 vccd1 vccd1 _18443_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_186_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15654_ _15654_/A vssd1 vssd1 vccd1 vccd1 _15656_/A sky130_fd_sc_hd__inv_2
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12866_ _26236_/Q _25605_/Q vssd1 vssd1 vccd1 vccd1 _14361_/A sky130_fd_sc_hd__xor2_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14605_ _14605_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14605_/Y sky130_fd_sc_hd__nand2_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18373_ _18535_/A _18373_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _18373_/X sky130_fd_sc_hd__and3_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15585_ _15795_/A _16520_/B vssd1 vssd1 vccd1 vccd1 _15588_/A sky130_fd_sc_hd__nor2_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12797_ _12746_/X _12795_/X _14910_/B _12796_/X vssd1 vssd1 vccd1 vccd1 _12797_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _17324_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17324_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_55_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14536_ _14536_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14536_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17255_ _17485_/A _17255_/B vssd1 vssd1 vccd1 vccd1 _17255_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_37_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14467_ _14464_/Y hold480/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold481/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16206_ _16206_/A _16206_/B vssd1 vssd1 vccd1 vccd1 _16207_/A sky130_fd_sc_hd__and2_1
XFILLER_0_10_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13418_ _13315_/X _13416_/X _23629_/B _13417_/X vssd1 vssd1 vccd1 vccd1 _13418_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17186_ _17448_/A _17186_/B vssd1 vssd1 vccd1 vccd1 _17186_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_113_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14398_ _14404_/A hold284/X vssd1 vssd1 vccd1 vccd1 hold285/A sky130_fd_sc_hd__nand2_1
XFILLER_0_144_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16137_ _22386_/B _16691_/B vssd1 vssd1 vccd1 vccd1 _16139_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_144_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13349_ _13220_/X _14629_/A _13242_/X _19659_/A vssd1 vssd1 vccd1 vccd1 _13349_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16068_ _16069_/B _16069_/A vssd1 vssd1 vccd1 vccd1 _16070_/A sky130_fd_sc_hd__or2_1
XFILLER_0_121_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15019_ _15019_/A _15029_/A vssd1 vssd1 vccd1 vccd1 _15019_/Y sky130_fd_sc_hd__nand2_1
Xhold2507 _26047_/Q vssd1 vssd1 vccd1 vccd1 hold2507/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2518 _12636_/X vssd1 vssd1 vccd1 vccd1 _12637_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2529 _25696_/Q vssd1 vssd1 vccd1 vccd1 _13383_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1806 _25862_/Q vssd1 vssd1 vccd1 vccd1 _22460_/B sky130_fd_sc_hd__dlygate4sd3_1
X_19827_ _26263_/Q hold847/X vssd1 vssd1 vccd1 vccd1 _19827_/Y sky130_fd_sc_hd__nand2_1
Xhold1817 _25906_/Q vssd1 vssd1 vccd1 vccd1 _23211_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1828 _22143_/Y vssd1 vssd1 vccd1 vccd1 _25850_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1839 _25905_/Q vssd1 vssd1 vccd1 vccd1 _17674_/A sky130_fd_sc_hd__buf_1
XFILLER_0_159_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19758_ _19758_/A _20479_/B vssd1 vssd1 vccd1 vccd1 _19758_/Y sky130_fd_sc_hd__nor2_1
X_18709_ _18792_/A _18713_/B vssd1 vssd1 vccd1 vccd1 _18711_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19689_ _20272_/A _19687_/Y _20277_/C vssd1 vssd1 vccd1 vccd1 _19779_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_149_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21720_ _21718_/Y _21719_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21720_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21651_ _21650_/Y _21203_/X _20986_/A _20957_/A vssd1 vssd1 vccd1 vccd1 _21651_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20602_ _20605_/A _20605_/C vssd1 vssd1 vccd1 vccd1 _20604_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24370_ _24370_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24371_/A sky130_fd_sc_hd__and2_1
XFILLER_0_157_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21582_ _21582_/A _21599_/B vssd1 vssd1 vccd1 vccd1 _21587_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_117_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23321_ _23321_/A _23377_/B _23321_/C vssd1 vssd1 vccd1 vccd1 _23321_/X sky130_fd_sc_hd__and3_1
XFILLER_0_89_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20533_ _21305_/B _21579_/A vssd1 vssd1 vccd1 vccd1 _20534_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_172_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23252_ _24949_/S vssd1 vssd1 vccd1 vccd1 _24959_/C sky130_fd_sc_hd__inv_2
X_26040_ _26040_/CLK _26040_/D vssd1 vssd1 vccd1 vccd1 _26040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20464_ _20660_/A _20464_/B vssd1 vssd1 vccd1 vccd1 _20464_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_171_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22203_ _22653_/A _22203_/B vssd1 vssd1 vccd1 vccd1 _22203_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23183_ _23183_/A _23183_/B vssd1 vssd1 vccd1 vccd1 _23185_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20395_ _20397_/B _20397_/C vssd1 vssd1 vccd1 vccd1 _20396_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22134_ _19206_/A _22133_/A _22133_/Y vssd1 vssd1 vccd1 vccd1 _22136_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22065_ _25812_/Q _22065_/B vssd1 vssd1 vccd1 vccd1 _22065_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_101_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21016_ _21042_/A _21016_/B _21015_/X vssd1 vssd1 vccd1 vccd1 _21017_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_173_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25824_ _25838_/CLK _25824_/D vssd1 vssd1 vccd1 vccd1 _25824_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_96_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25755_ _25756_/CLK _25755_/D vssd1 vssd1 vccd1 vccd1 _25755_/Q sky130_fd_sc_hd__dfxtp_1
X_22967_ _22967_/A _23001_/B _22967_/C vssd1 vssd1 vccd1 vccd1 _22967_/X sky130_fd_sc_hd__and3_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12720_ _14270_/B _23193_/B vssd1 vssd1 vccd1 vccd1 _17009_/B sky130_fd_sc_hd__nand2_4
X_24706_ _24706_/A vssd1 vssd1 vccd1 vccd1 _26297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21918_ _21918_/A _22689_/B vssd1 vssd1 vccd1 vccd1 _21919_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25686_ _25689_/CLK _25686_/D vssd1 vssd1 vccd1 vccd1 _25686_/Q sky130_fd_sc_hd__dfxtp_1
X_22898_ _22898_/A _23001_/B _22898_/C vssd1 vssd1 vccd1 vccd1 _22898_/X sky130_fd_sc_hd__and3_1
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12651_ _12651_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _12651_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_155_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24637_ _24637_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24638_/A sky130_fd_sc_hd__and2_1
X_21849_ _21849_/A _22637_/B vssd1 vssd1 vccd1 vccd1 _21850_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_66_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15370_ _16356_/A _16711_/A vssd1 vssd1 vccd1 vccd1 _16810_/A sky130_fd_sc_hd__nand2_2
X_12582_ _12582_/A _23924_/A vssd1 vssd1 vccd1 vccd1 _12582_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24568_ _24568_/A vssd1 vssd1 vccd1 vccd1 _26252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14321_ _14319_/Y hold189/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold190/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26307_ _26308_/CLK _26307_/D vssd1 vssd1 vccd1 vccd1 _26307_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_80_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23519_ _23513_/X _23518_/X _24958_/B vssd1 vssd1 vccd1 vccd1 _23519_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24499_ _24499_/A _24557_/B vssd1 vssd1 vccd1 vccd1 _24500_/A sky130_fd_sc_hd__and2_1
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17040_ _25625_/Q vssd1 vssd1 vccd1 vccd1 _20163_/B sky130_fd_sc_hd__inv_2
X_26238_ _26239_/CLK _26238_/D vssd1 vssd1 vccd1 vccd1 _26238_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_52_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14252_ _14264_/A _14252_/B vssd1 vssd1 vccd1 vccd1 _14252_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13203_ _13049_/X _14557_/A _13067_/X _19331_/A vssd1 vssd1 vccd1 vccd1 _13203_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_180_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14183_ _25824_/Q vssd1 vssd1 vccd1 vccd1 _18694_/B sky130_fd_sc_hd__inv_2
X_26169_ _26171_/CLK _26169_/D vssd1 vssd1 vccd1 vccd1 _26169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13134_ _13109_/X _13132_/X _13096_/X _13133_/X vssd1 vssd1 vccd1 vccd1 _13134_/X
+ sky130_fd_sc_hd__o211a_1
X_18991_ _18989_/X _18879_/X _18990_/X vssd1 vssd1 vccd1 vccd1 _18992_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_21_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17942_ _17942_/A _25787_/Q _17942_/C vssd1 vssd1 vccd1 vccd1 _20513_/B sky130_fd_sc_hd__nand3_2
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _14262_/B vssd1 vssd1 vccd1 vccd1 _13065_/X sky130_fd_sc_hd__buf_12
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17873_ _17873_/A _17873_/B _20114_/A vssd1 vssd1 vccd1 vccd1 _17883_/A sky130_fd_sc_hd__and3_1
XFILLER_0_136_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16824_ _16824_/A _16824_/B vssd1 vssd1 vccd1 vccd1 _16824_/Y sky130_fd_sc_hd__nand2_1
X_19612_ _26248_/Q _19483_/X hold401/X vssd1 vssd1 vccd1 vccd1 _19612_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19543_ _26243_/Q hold629/X vssd1 vssd1 vccd1 vccd1 _19543_/Y sky130_fd_sc_hd__nand2_1
X_16755_ _16753_/X _16711_/X _16754_/Y _25868_/Q _14170_/X vssd1 vssd1 vccd1 vccd1
+ _16756_/A sky130_fd_sc_hd__a32o_1
X_13967_ _13962_/Y _13966_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold854/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15706_ _15706_/A _15774_/B vssd1 vssd1 vccd1 vccd1 _15707_/B sky130_fd_sc_hd__nand2_1
X_12918_ _17424_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12918_/X sky130_fd_sc_hd__or2_1
X_19474_ _21101_/A _21844_/B _25613_/Q vssd1 vssd1 vccd1 vccd1 _21105_/C sky130_fd_sc_hd__nand3_1
X_16686_ _16686_/A _16686_/B _16695_/A vssd1 vssd1 vccd1 vccd1 _16686_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13898_ _13941_/A _13898_/B vssd1 vssd1 vccd1 vccd1 _13898_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18425_ _18445_/A _18429_/B vssd1 vssd1 vccd1 vccd1 _18427_/A sky130_fd_sc_hd__nand2_1
X_15637_ _15637_/A vssd1 vssd1 vccd1 vccd1 _16561_/A sky130_fd_sc_hd__inv_2
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12849_ _17282_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12849_/X sky130_fd_sc_hd__or2_1
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18356_ _18641_/A _19257_/A vssd1 vssd1 vccd1 vccd1 _18356_/Y sky130_fd_sc_hd__nand2_1
X_15568_ _15568_/A vssd1 vssd1 vccd1 vccd1 _16510_/A sky130_fd_sc_hd__inv_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17307_ _17563_/A _17644_/A vssd1 vssd1 vccd1 vccd1 _17308_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14519_ _14525_/A hold8/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__nand2_1
XFILLER_0_83_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18287_ _18952_/A _18287_/B _18952_/C vssd1 vssd1 vccd1 vccd1 _18288_/C sky130_fd_sc_hd__nand3_1
X_15499_ _15500_/B _15500_/A vssd1 vssd1 vccd1 vccd1 _15499_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17238_ _17527_/A _17607_/A vssd1 vssd1 vccd1 vccd1 _17239_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold903 hold903/A vssd1 vssd1 vccd1 vccd1 hold903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 hold914/A vssd1 vssd1 vccd1 vccd1 hold914/X sky130_fd_sc_hd__dlygate4sd3_1
X_17169_ _25634_/Q vssd1 vssd1 vccd1 vccd1 _20518_/B sky130_fd_sc_hd__inv_2
Xhold925 hold925/A vssd1 vssd1 vccd1 vccd1 hold925/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold936 hold936/A vssd1 vssd1 vccd1 vccd1 hold936/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold947 hold947/A vssd1 vssd1 vccd1 vccd1 hold947/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 hold958/A vssd1 vssd1 vccd1 vccd1 hold958/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_20180_ _20180_/A _20180_/B _20180_/C vssd1 vssd1 vccd1 vccd1 _20181_/B sky130_fd_sc_hd__nand3_1
Xhold969 hold969/A vssd1 vssd1 vccd1 vccd1 hold969/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2304 _25432_/Q vssd1 vssd1 vccd1 vccd1 _15065_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2315 _24984_/Q vssd1 vssd1 vccd1 vccd1 _12659_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2326 _26084_/Q vssd1 vssd1 vccd1 vccd1 hold2326/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2337 _25418_/Q vssd1 vssd1 vccd1 vccd1 _14945_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1603 _17387_/Y vssd1 vssd1 vccd1 vccd1 _25610_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2348 _25672_/Q vssd1 vssd1 vccd1 vccd1 _13233_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1614 _25613_/Q vssd1 vssd1 vccd1 vccd1 _17417_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2359 _25670_/Q vssd1 vssd1 vccd1 vccd1 _13221_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1625 _20388_/Y vssd1 vssd1 vccd1 vccd1 _25783_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1636 _21704_/Y vssd1 vssd1 vccd1 vccd1 _25836_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23870_ _23870_/A vssd1 vssd1 vccd1 vccd1 _26027_/D sky130_fd_sc_hd__clkbuf_1
Xhold1647 _25648_/Q vssd1 vssd1 vccd1 vccd1 _17917_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1658 _17347_/Y vssd1 vssd1 vccd1 vccd1 _25606_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1669 _25605_/Q vssd1 vssd1 vccd1 vccd1 _17336_/B sky130_fd_sc_hd__dlygate4sd3_1
X_22821_ _22937_/A _22821_/B vssd1 vssd1 vccd1 vccd1 _22821_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25540_ _26047_/CLK _25540_/D vssd1 vssd1 vccd1 vccd1 _25540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22752_ _22752_/A _23001_/B _22752_/C vssd1 vssd1 vccd1 vccd1 _22752_/X sky130_fd_sc_hd__and3_1
XFILLER_0_17_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21703_ _22058_/A _21703_/B vssd1 vssd1 vccd1 vccd1 _21703_/Y sky130_fd_sc_hd__nand2_1
X_25471_ _25532_/CLK _25471_/D vssd1 vssd1 vccd1 vccd1 _25471_/Q sky130_fd_sc_hd__dfxtp_1
X_22683_ _22683_/A _22683_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22685_/A sky130_fd_sc_hd__or3_1
XFILLER_0_48_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24422_ _24422_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24423_/A sky130_fd_sc_hd__and2_1
X_21634_ _26335_/Q hold383/X vssd1 vssd1 vccd1 vccd1 _21634_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_35_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24353_ hold2392/X _26183_/Q _24356_/S vssd1 vssd1 vccd1 vccd1 _24353_/X sky130_fd_sc_hd__mux2_1
X_21565_ _21565_/A _21565_/B vssd1 vssd1 vccd1 vccd1 _21566_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23304_ hold986/X _23303_/Y _12702_/A vssd1 vssd1 vccd1 vccd1 hold987/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20516_ _21305_/B vssd1 vssd1 vccd1 vccd1 _21302_/C sky130_fd_sc_hd__inv_2
XFILLER_0_127_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24284_ _24560_/A vssd1 vssd1 vccd1 vccd1 _24373_/B sky130_fd_sc_hd__buf_6
X_21496_ _21498_/A _21547_/A vssd1 vssd1 vccd1 vccd1 _21497_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_90_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23235_ _23235_/A vssd1 vssd1 vccd1 vccd1 _25910_/D sky130_fd_sc_hd__clkbuf_1
X_26023_ _26023_/CLK _26023_/D vssd1 vssd1 vccd1 vccd1 _26023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20447_ _20447_/A _20447_/B _20447_/C vssd1 vssd1 vccd1 vccd1 _20448_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_160_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23166_ _23164_/X _23165_/Y _12702_/A vssd1 vssd1 vccd1 vccd1 _23166_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20378_ _20378_/A _21117_/B _20378_/C vssd1 vssd1 vccd1 vccd1 _20379_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_101_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22117_ _22115_/X _15839_/B _22116_/Y _14813_/B _21725_/X vssd1 vssd1 vccd1 vccd1
+ _22118_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_63_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23097_ _23097_/A _23193_/B _23097_/C vssd1 vssd1 vccd1 vccd1 _23097_/X sky130_fd_sc_hd__and3_1
XFILLER_0_101_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22048_ _22048_/A _22759_/A vssd1 vssd1 vccd1 vccd1 _22055_/A sky130_fd_sc_hd__nand2_1
X_14870_ _25857_/Q _12527_/A _15058_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14870_/X
+ sky130_fd_sc_hd__a22o_1
X_13821_ _18813_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13821_/Y sky130_fd_sc_hd__nor2_1
X_25807_ _25807_/CLK _25807_/D vssd1 vssd1 vccd1 vccd1 _25807_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_98_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23999_ _23999_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _24000_/A sky130_fd_sc_hd__and2_1
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16540_ _16538_/X _16539_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 _16540_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25738_ _25738_/CLK _25738_/D vssd1 vssd1 vccd1 vccd1 _25738_/Q sky130_fd_sc_hd__dfxtp_1
X_13752_ _13823_/A _13752_/B vssd1 vssd1 vccd1 vccd1 _13752_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12703_ hold997/X _12704_/A _12702_/Y vssd1 vssd1 vccd1 vccd1 hold998/A sky130_fd_sc_hd__o21a_1
X_16471_ _16480_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16471_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_167_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25669_ _26299_/CLK _25669_/D vssd1 vssd1 vccd1 vccd1 _25669_/Q sky130_fd_sc_hd__dfxtp_1
X_13683_ _18367_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13683_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18210_ _21791_/A vssd1 vssd1 vccd1 vccd1 _18579_/B sky130_fd_sc_hd__clkbuf_8
X_15422_ _15422_/A vssd1 vssd1 vccd1 vccd1 _16401_/A sky130_fd_sc_hd__inv_2
X_12634_ _12654_/A vssd1 vssd1 vccd1 vccd1 _12636_/A sky130_fd_sc_hd__inv_2
XFILLER_0_38_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19190_ _19211_/B _19280_/B vssd1 vssd1 vccd1 vccd1 _19191_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18141_ _18141_/A _20908_/A vssd1 vssd1 vccd1 vccd1 _18514_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_108_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15353_ _15353_/A vssd1 vssd1 vccd1 vccd1 _16346_/A sky130_fd_sc_hd__inv_2
X_12565_ _12570_/A _24836_/B _12565_/C vssd1 vssd1 vccd1 vccd1 _12566_/A sky130_fd_sc_hd__and3_1
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14304_ _14304_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14304_/Y sky130_fd_sc_hd__nand2_1
X_18072_ _18074_/A _18074_/C vssd1 vssd1 vccd1 vccd1 _18073_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15284_ _15284_/A _15810_/B vssd1 vssd1 vccd1 vccd1 _15285_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12496_ _12496_/A vssd1 vssd1 vccd1 vccd1 _23199_/C sky130_fd_sc_hd__inv_2
XFILLER_0_123_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17023_ _25654_/Q _17023_/B vssd1 vssd1 vccd1 vccd1 _17413_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14235_ hold384/X _14234_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold385/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14166_ _26324_/Q _13988_/X _13981_/X _14165_/Y vssd1 vssd1 vccd1 vccd1 _14167_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _26155_/Q _13065_/X _13116_/X vssd1 vssd1 vccd1 vccd1 _13117_/X sky130_fd_sc_hd__a21o_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _26313_/Q _13988_/X _13981_/X _14096_/Y vssd1 vssd1 vccd1 vccd1 _14098_/B
+ sky130_fd_sc_hd__a22o_1
X_18974_ _18974_/A _19045_/A vssd1 vssd1 vccd1 vccd1 _18975_/B sky130_fd_sc_hd__xnor2_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _13018_/X _13046_/X _13005_/X _13047_/X vssd1 vssd1 vccd1 vccd1 _13048_/X
+ sky130_fd_sc_hd__o211a_1
X_17925_ _17925_/A _17925_/B vssd1 vssd1 vccd1 vccd1 _17927_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_147_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17856_ _17856_/A _25785_/Q _17856_/C vssd1 vssd1 vccd1 vccd1 _20434_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_179_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16807_ _16805_/Y _16806_/Y _16791_/X vssd1 vssd1 vccd1 vccd1 _16807_/Y sky130_fd_sc_hd__a21oi_1
X_17787_ _22786_/A _17763_/Y _17780_/B _17784_/B vssd1 vssd1 vccd1 vccd1 _18153_/C
+ sky130_fd_sc_hd__o211ai_4
X_14999_ _14981_/B _14998_/B _14990_/B vssd1 vssd1 vccd1 vccd1 _14999_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_152_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16738_ _16980_/A _16743_/B vssd1 vssd1 vccd1 vccd1 _16740_/B sky130_fd_sc_hd__nand2_1
X_19526_ _19723_/A _19526_/B vssd1 vssd1 vccd1 vccd1 _19526_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_92_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19457_ _19454_/Y _19457_/B _19980_/B vssd1 vssd1 vccd1 vccd1 _19457_/X sky130_fd_sc_hd__and3b_1
X_16669_ _16669_/A vssd1 vssd1 vccd1 vccd1 _16670_/B sky130_fd_sc_hd__inv_2
XFILLER_0_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18408_ _18793_/A _18408_/B _18894_/C vssd1 vssd1 vccd1 vccd1 _18409_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19388_ _19388_/A _20936_/B vssd1 vssd1 vccd1 vccd1 _19388_/Y sky130_fd_sc_hd__nor2_1
X_18339_ _21913_/B _25615_/Q vssd1 vssd1 vccd1 vccd1 _18341_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_189_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21350_ _21401_/A _21707_/C vssd1 vssd1 vccd1 vccd1 _21351_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_25_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20301_ _26284_/Q _20078_/X hold736/X vssd1 vssd1 vccd1 vccd1 _20304_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_170_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold700 hold700/A vssd1 vssd1 vccd1 vccd1 hold700/X sky130_fd_sc_hd__dlygate4sd3_1
X_21281_ _21281_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _21286_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_141_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold711 hold711/A vssd1 vssd1 vccd1 vccd1 hold711/X sky130_fd_sc_hd__dlygate4sd3_1
X_23020_ _23011_/Y _23019_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _23020_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_124_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold722 hold722/A vssd1 vssd1 vccd1 vccd1 hold722/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20232_ _20232_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _20232_/Y sky130_fd_sc_hd__nand2_1
Xhold733 hold733/A vssd1 vssd1 vccd1 vccd1 hold733/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 hold744/A vssd1 vssd1 vccd1 vccd1 hold744/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 hold755/A vssd1 vssd1 vccd1 vccd1 hold755/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold766 hold766/A vssd1 vssd1 vccd1 vccd1 hold766/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 hold777/A vssd1 vssd1 vccd1 vccd1 hold777/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 hold788/A vssd1 vssd1 vccd1 vccd1 hold788/X sky130_fd_sc_hd__dlygate4sd3_1
X_20163_ _20163_/A _20163_/B vssd1 vssd1 vccd1 vccd1 _20167_/A sky130_fd_sc_hd__nand2_1
Xhold799 hold799/A vssd1 vssd1 vccd1 vccd1 hold799/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2101 _25948_/Q vssd1 vssd1 vccd1 vccd1 hold2101/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2112 _25927_/Q vssd1 vssd1 vccd1 vccd1 _23324_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2123 _26007_/Q vssd1 vssd1 vccd1 vccd1 hold2123/X sky130_fd_sc_hd__dlygate4sd3_1
X_24971_ _25420_/CLK _24971_/D vssd1 vssd1 vccd1 vccd1 _24971_/Q sky130_fd_sc_hd__dfxtp_1
X_20094_ _20094_/A _20094_/B vssd1 vssd1 vccd1 vccd1 _20096_/A sky130_fd_sc_hd__nand2_1
Xhold2134 _26088_/Q vssd1 vssd1 vccd1 vccd1 hold2134/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2145 _26107_/Q vssd1 vssd1 vccd1 vccd1 hold2145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1400 _19354_/Y vssd1 vssd1 vccd1 vccd1 _25726_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1411 _25560_/Q vssd1 vssd1 vccd1 vccd1 _16842_/B sky130_fd_sc_hd__buf_1
Xhold2156 _25990_/Q vssd1 vssd1 vccd1 vccd1 hold2156/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2167 _26019_/Q vssd1 vssd1 vccd1 vccd1 hold2167/X sky130_fd_sc_hd__dlygate4sd3_1
X_23922_ _23922_/A vssd1 vssd1 vccd1 vccd1 _26044_/D sky130_fd_sc_hd__clkbuf_1
Xhold1422 _12839_/X vssd1 vssd1 vccd1 vccd1 _25019_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1433 _25104_/Q vssd1 vssd1 vccd1 vccd1 _18799_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2178 _26062_/Q vssd1 vssd1 vccd1 vccd1 hold2178/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1444 _16915_/Y vssd1 vssd1 vccd1 vccd1 _25570_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2189 _26129_/Q vssd1 vssd1 vccd1 vccd1 hold2189/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 _25399_/Q vssd1 vssd1 vccd1 vccd1 _14795_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1466 _13007_/X vssd1 vssd1 vccd1 vccd1 _25051_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23853_ hold2070/X hold2039/X _23907_/S vssd1 vssd1 vccd1 vccd1 _23854_/A sky130_fd_sc_hd__mux2_1
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1477 _25389_/Q vssd1 vssd1 vccd1 vccd1 _14703_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1488 _13270_/X vssd1 vssd1 vccd1 vccd1 _25097_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 _25896_/Q vssd1 vssd1 vccd1 vccd1 _23117_/B sky130_fd_sc_hd__buf_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22804_ _22795_/Y _22803_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22804_/X sky130_fd_sc_hd__a21o_1
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23784_ _23784_/A vssd1 vssd1 vccd1 vccd1 _25999_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20996_ _20996_/A _25865_/Q vssd1 vssd1 vccd1 vccd1 _21002_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_95_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25523_ _25534_/CLK _25523_/D vssd1 vssd1 vccd1 vccd1 _25523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22735_ _22734_/A _22454_/X _22734_/B vssd1 vssd1 vccd1 vccd1 _22736_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25454_ _26060_/CLK _25454_/D vssd1 vssd1 vccd1 vccd1 _25454_/Q sky130_fd_sc_hd__dfxtp_1
X_22666_ _18917_/A _25835_/Q _22664_/Y _22665_/Y vssd1 vssd1 vccd1 vccd1 _22667_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_94_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24405_ _24405_/A vssd1 vssd1 vccd1 vccd1 _26199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21617_ _26334_/Q _19130_/X hold566/X vssd1 vssd1 vccd1 vccd1 _21620_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25385_ _26336_/CLK hold352/X vssd1 vssd1 vccd1 vccd1 hold350/A sky130_fd_sc_hd__dfxtp_1
X_22597_ _23104_/B vssd1 vssd1 vccd1 vccd1 _23103_/B sky130_fd_sc_hd__inv_2
XFILLER_0_118_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24336_ _24336_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24337_/A sky130_fd_sc_hd__and2_1
XFILLER_0_133_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21548_ _21548_/A _21548_/B _21548_/C vssd1 vssd1 vccd1 vccd1 _21549_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24267_ hold2221/X hold2201/X _24279_/S vssd1 vssd1 vccd1 vccd1 _24268_/A sky130_fd_sc_hd__mux2_1
X_21479_ _21530_/A _21482_/A vssd1 vssd1 vccd1 vccd1 _21480_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_121_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26006_ _26073_/CLK _26006_/D vssd1 vssd1 vccd1 vccd1 _26006_/Q sky130_fd_sc_hd__dfxtp_1
X_14020_ _14118_/A hold635/X vssd1 vssd1 vccd1 vccd1 hold636/A sky130_fd_sc_hd__nand2_1
X_23218_ _23278_/B _24956_/S vssd1 vssd1 vccd1 vccd1 _23220_/A sky130_fd_sc_hd__or2_1
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24198_ _24198_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24199_/A sky130_fd_sc_hd__and2_1
X_23149_ _23197_/A _23149_/B vssd1 vssd1 vccd1 vccd1 _23149_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15971_ _15971_/A _15971_/B vssd1 vssd1 vccd1 vccd1 _15972_/B sky130_fd_sc_hd__nand2_1
X_17710_ _17759_/C _17738_/A vssd1 vssd1 vccd1 vccd1 _17737_/A sky130_fd_sc_hd__nand2_1
X_14922_ _14923_/B _14923_/A vssd1 vssd1 vccd1 vccd1 _14924_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_101_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18690_ _18952_/A _25760_/Q _18891_/C vssd1 vssd1 vccd1 vccd1 _18691_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2690 _26218_/Q vssd1 vssd1 vccd1 vccd1 hold2690/X sky130_fd_sc_hd__dlygate4sd3_1
X_17641_ _17641_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _17641_/Y sky130_fd_sc_hd__nand2_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
X_14853_ _22262_/B _15543_/B vssd1 vssd1 vccd1 vccd1 _14854_/A sky130_fd_sc_hd__nand2_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
X_13804_ _26266_/Q _13801_/X _13793_/X _13803_/Y vssd1 vssd1 vccd1 vccd1 _13805_/B
+ sky130_fd_sc_hd__a22o_1
X_17572_ _17624_/A _17572_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17572_/X sky130_fd_sc_hd__and3_1
X_14784_ _25847_/Q _13466_/A _14783_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14785_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19311_ _19452_/A _19311_/B vssd1 vssd1 vccd1 vccd1 _19311_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16523_ _16537_/B _16523_/B vssd1 vssd1 vccd1 vccd1 _16541_/A sky130_fd_sc_hd__and2_1
XFILLER_0_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13735_ hold381/X _13734_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold382/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_168_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19242_ _19452_/A hold922/X vssd1 vssd1 vccd1 vccd1 hold923/A sky130_fd_sc_hd__nand2_1
X_16454_ _16437_/B _16437_/A _16447_/C vssd1 vssd1 vccd1 vccd1 _16456_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13666_ _13703_/A _13666_/B vssd1 vssd1 vccd1 vccd1 _13666_/Y sky130_fd_sc_hd__nand2_1
X_15405_ _15405_/A _15405_/B vssd1 vssd1 vccd1 vccd1 _15406_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _12618_/B _12618_/A vssd1 vssd1 vccd1 vccd1 _12624_/A sky130_fd_sc_hd__or2_1
XFILLER_0_27_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19173_ _19172_/Y _19130_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19175_/A
+ sky130_fd_sc_hd__a211o_1
X_16385_ _16337_/X _16380_/A _16384_/X vssd1 vssd1 vccd1 vccd1 _16393_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_115_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13597_ hold456/X _13596_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold457/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_171_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18124_ _18124_/A _18124_/B vssd1 vssd1 vccd1 vccd1 _18126_/A sky130_fd_sc_hd__nand2_1
X_15336_ _22747_/B _16369_/B vssd1 vssd1 vccd1 vccd1 _16329_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12548_ _13465_/A _24871_/B _12548_/C vssd1 vssd1 vccd1 vccd1 _17742_/A sky130_fd_sc_hd__and3_4
XFILLER_0_42_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18055_ _18055_/A _20855_/A vssd1 vssd1 vccd1 vccd1 _18474_/A sky130_fd_sc_hd__xor2_4
X_15267_ _15267_/A vssd1 vssd1 vccd1 vccd1 _15268_/A sky130_fd_sc_hd__inv_2
XFILLER_0_151_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_2 _21007_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17006_ _17393_/A hold77/X _19994_/B vssd1 vssd1 vccd1 vccd1 _17006_/X sky130_fd_sc_hd__and3_1
XFILLER_0_151_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14218_ _14236_/A hold398/X vssd1 vssd1 vccd1 vccd1 hold399/A sky130_fd_sc_hd__nand2_1
XFILLER_0_123_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15198_ _15198_/A _16740_/A vssd1 vssd1 vccd1 vccd1 _15199_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14149_ hold435/X _14148_/Y _14037_/X vssd1 vssd1 vccd1 vccd1 hold436/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18957_ _20094_/B _22720_/A vssd1 vssd1 vccd1 vccd1 _20087_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17908_ _18529_/A _17908_/B _18083_/C vssd1 vssd1 vccd1 vccd1 _17909_/C sky130_fd_sc_hd__nand3_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18888_ _18888_/A _18888_/B vssd1 vssd1 vccd1 vccd1 _22639_/A sky130_fd_sc_hd__or2_1
X_17839_ _20702_/B _19289_/A vssd1 vssd1 vccd1 vccd1 _17840_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_89_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20850_ _21042_/A _20850_/B _20849_/X vssd1 vssd1 vccd1 vccd1 _20851_/B sky130_fd_sc_hd__or3b_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19509_ _19509_/A _19509_/B vssd1 vssd1 vccd1 vccd1 _19509_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20781_ _20784_/A _20784_/C vssd1 vssd1 vccd1 vccd1 _20782_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22520_ _23056_/B vssd1 vssd1 vccd1 vccd1 _23055_/B sky130_fd_sc_hd__inv_2
XFILLER_0_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22451_ _26045_/Q vssd1 vssd1 vccd1 vccd1 _22453_/A sky130_fd_sc_hd__inv_2
XFILLER_0_135_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21402_ _21402_/A _21450_/A vssd1 vssd1 vccd1 vccd1 _21403_/C sky130_fd_sc_hd__nand2_1
X_22382_ _22380_/X _22381_/Y _22900_/B vssd1 vssd1 vccd1 vccd1 _22382_/Y sky130_fd_sc_hd__a21oi_1
X_25170_ _25759_/CLK hold926/X vssd1 vssd1 vccd1 vccd1 hold925/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24121_ _24121_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24122_/A sky130_fd_sc_hd__and2_1
X_21333_ _21694_/B _21386_/A vssd1 vssd1 vccd1 vccd1 _21335_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_143_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24052_ _24835_/S vssd1 vssd1 vccd1 vccd1 _24126_/S sky130_fd_sc_hd__clkbuf_16
Xhold530 hold530/A vssd1 vssd1 vccd1 vccd1 hold530/X sky130_fd_sc_hd__dlygate4sd3_1
X_21264_ _21264_/A _22040_/B vssd1 vssd1 vccd1 vccd1 _21265_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold541 hold541/A vssd1 vssd1 vccd1 vccd1 hold541/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 hold552/A vssd1 vssd1 vccd1 vccd1 hold552/X sky130_fd_sc_hd__dlygate4sd3_1
X_23003_ _23003_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _23003_/Y sky130_fd_sc_hd__nand2_1
Xhold563 hold563/A vssd1 vssd1 vccd1 vccd1 hold563/X sky130_fd_sc_hd__dlygate4sd3_1
X_20215_ _20217_/B _20217_/C vssd1 vssd1 vccd1 vccd1 _20216_/A sky130_fd_sc_hd__nand2_1
Xhold574 hold574/A vssd1 vssd1 vccd1 vccd1 hold574/X sky130_fd_sc_hd__dlygate4sd3_1
X_21195_ _21195_/A _21195_/B _21195_/C vssd1 vssd1 vccd1 vccd1 _21199_/A sky130_fd_sc_hd__nand3_1
Xhold585 hold585/A vssd1 vssd1 vccd1 vccd1 hold585/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold596 hold596/A vssd1 vssd1 vccd1 vccd1 hold596/X sky130_fd_sc_hd__dlygate4sd3_1
X_20146_ _21418_/A _21033_/C vssd1 vssd1 vccd1 vccd1 _20151_/A sky130_fd_sc_hd__nand2_1
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24954_ _24951_/X _24957_/S _24958_/B _24953_/X vssd1 vssd1 vccd1 vccd1 _24954_/X
+ sky130_fd_sc_hd__a211o_2
X_20077_ _20077_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20083_/A sky130_fd_sc_hd__nand2_2
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1230 _25793_/Q vssd1 vssd1 vccd1 vccd1 _20777_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1241 _19853_/Y vssd1 vssd1 vccd1 vccd1 _25761_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23905_ _23905_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23906_/A sky130_fd_sc_hd__and2_1
Xhold1252 _25087_/Q vssd1 vssd1 vccd1 vccd1 _18455_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24885_ _24885_/A _24946_/A vssd1 vssd1 vccd1 vccd1 _24885_/Y sky130_fd_sc_hd__nand2_1
Xhold1263 _19797_/Y vssd1 vssd1 vccd1 vccd1 _25757_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 _25543_/Q vssd1 vssd1 vccd1 vccd1 _16729_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1285 _19326_/Y vssd1 vssd1 vccd1 vccd1 _25724_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1296 _25794_/Q vssd1 vssd1 vccd1 vccd1 _20815_/B sky130_fd_sc_hd__buf_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23836_ _23836_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23837_/A sky130_fd_sc_hd__and2_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23767_ _14806_/B _25994_/Q _23831_/S vssd1 vssd1 vccd1 vccd1 _23767_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_94_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20979_ _21464_/C _21516_/B vssd1 vssd1 vccd1 vccd1 _20981_/A sky130_fd_sc_hd__nand2_1
X_25506_ _25510_/CLK hold890/X vssd1 vssd1 vccd1 vccd1 hold889/A sky130_fd_sc_hd__dfxtp_1
X_13520_ _13583_/A _13520_/B vssd1 vssd1 vccd1 vccd1 _13520_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22718_ _25837_/Q _22718_/B vssd1 vssd1 vccd1 vccd1 _22718_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_83_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23698_ _23698_/A vssd1 vssd1 vccd1 vccd1 _25971_/D sky130_fd_sc_hd__clkbuf_1
X_25437_ _25501_/CLK _25437_/D vssd1 vssd1 vccd1 vccd1 _25437_/Q sky130_fd_sc_hd__dfxtp_1
X_13451_ _19068_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13451_/X sky130_fd_sc_hd__or2_1
X_22649_ _22991_/B _23136_/B vssd1 vssd1 vccd1 vccd1 _22650_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16170_ _16172_/B vssd1 vssd1 vccd1 vccd1 _16189_/B sky130_fd_sc_hd__inv_2
X_13382_ _13315_/X _13380_/X _13300_/X _13381_/X vssd1 vssd1 vccd1 vccd1 _13382_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25368_ _26193_/CLK hold151/X vssd1 vssd1 vccd1 vccd1 hold149/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15121_ hold931/X vssd1 vssd1 vccd1 vccd1 _15123_/A sky130_fd_sc_hd__inv_2
XFILLER_0_140_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24319_ _24319_/A vssd1 vssd1 vccd1 vccd1 _26171_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25299_ _25716_/CLK hold409/X vssd1 vssd1 vccd1 vccd1 hold407/A sky130_fd_sc_hd__dfxtp_1
X_15052_ _15028_/B _15051_/B _15043_/B vssd1 vssd1 vccd1 vccd1 _15052_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_142_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14003_ _18003_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14003_/Y sky130_fd_sc_hd__nor2_1
X_19860_ _19937_/A _19875_/B vssd1 vssd1 vccd1 vccd1 _19862_/A sky130_fd_sc_hd__xnor2_1
X_18811_ _18811_/A _25830_/Q _18811_/C vssd1 vssd1 vccd1 vccd1 _20681_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19791_ _19807_/B _19875_/B vssd1 vssd1 vccd1 vccd1 _19793_/A sky130_fd_sc_hd__xnor2_1
X_15954_ _15961_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _15954_/Y sky130_fd_sc_hd__nand2_1
X_18742_ _18986_/A _19532_/A vssd1 vssd1 vccd1 vccd1 _18742_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14905_ _23245_/A _14905_/B _14909_/B vssd1 vssd1 vccd1 vccd1 _14905_/X sky130_fd_sc_hd__or3_1
X_18673_ _18793_/A _18673_/B _18894_/C vssd1 vssd1 vccd1 vccd1 _18674_/C sky130_fd_sc_hd__nand3_1
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15885_ _15883_/X _15884_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _15885_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_196_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _26117_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14836_ _15021_/B vssd1 vssd1 vccd1 vccd1 _14836_/Y sky130_fd_sc_hd__inv_2
X_17624_ _17624_/A _17624_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _17624_/X sky130_fd_sc_hd__and3_1
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ _17555_/A _17607_/A vssd1 vssd1 vccd1 vccd1 _17556_/B sky130_fd_sc_hd__xnor2_1
X_14767_ _14767_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14767_/Y sky130_fd_sc_hd__nand2_1
X_16506_ _16698_/A hold745/X vssd1 vssd1 vccd1 vccd1 hold746/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13718_ _13760_/A hold925/X vssd1 vssd1 vccd1 vccd1 _13718_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17486_ _17624_/A _17486_/B _17572_/C vssd1 vssd1 vccd1 vccd1 _17486_/X sky130_fd_sc_hd__and3_1
X_14698_ _25838_/Q _13466_/A _14697_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14701_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16437_ _16437_/A _16437_/B vssd1 vssd1 vccd1 vccd1 _16438_/B sky130_fd_sc_hd__and2_1
X_19225_ _19225_/A _19994_/B _19225_/C vssd1 vssd1 vccd1 vccd1 _19225_/X sky130_fd_sc_hd__and3_1
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13649_ _14125_/A vssd1 vssd1 vccd1 vccd1 _13760_/A sky130_fd_sc_hd__buf_6
XFILLER_0_183_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19156_ _26216_/Q _19134_/X hold413/X vssd1 vssd1 vccd1 vccd1 _19157_/C sky130_fd_sc_hd__a21o_1
X_16368_ _16366_/Y _16367_/Y _16343_/X vssd1 vssd1 vccd1 vccd1 hold951/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18107_ _18535_/A _18107_/B _18393_/C vssd1 vssd1 vccd1 vccd1 _18107_/X sky130_fd_sc_hd__and3_1
X_15319_ _15320_/B _16787_/A vssd1 vssd1 vccd1 vccd1 _15321_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19087_ _19084_/Y _19085_/Y _19086_/X vssd1 vssd1 vccd1 vccd1 _25709_/D sky130_fd_sc_hd__a21oi_1
X_16299_ _16299_/A _16309_/B vssd1 vssd1 vccd1 vccd1 _16299_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_152_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_120_clk clkbuf_4_14__f_clk/X vssd1 vssd1 vccd1 vccd1 _26330_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_160_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18038_ _19345_/A vssd1 vssd1 vccd1 vccd1 _21835_/B sky130_fd_sc_hd__inv_2
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20000_ _20000_/A _20000_/B vssd1 vssd1 vccd1 vccd1 _20004_/A sky130_fd_sc_hd__nand2_1
X_19989_ _19989_/A _19989_/B vssd1 vssd1 vccd1 vccd1 _19990_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21951_ _22715_/B _21952_/A vssd1 vssd1 vccd1 vccd1 _21953_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_187_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _25781_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20902_ _20901_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20902_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_179_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24670_ _24670_/A vssd1 vssd1 vccd1 vccd1 _26285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21882_ _25870_/Q _21883_/A vssd1 vssd1 vccd1 vccd1 _21884_/A sky130_fd_sc_hd__or2_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23621_ _23621_/A vssd1 vssd1 vccd1 vccd1 _25946_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20833_ _20833_/A _22645_/B _20833_/C vssd1 vssd1 vccd1 vccd1 _20836_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26340_ _26340_/CLK _26340_/D vssd1 vssd1 vccd1 vccd1 _26340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23552_ _24942_/S hold260/A _23551_/X vssd1 vssd1 vccd1 vccd1 _23552_/Y sky130_fd_sc_hd__o21ai_1
X_20764_ _20764_/A _20764_/B _21354_/B vssd1 vssd1 vccd1 vccd1 _20768_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22503_ _26047_/Q vssd1 vssd1 vccd1 vccd1 _22504_/A sky130_fd_sc_hd__inv_2
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26271_ _26273_/CLK _26271_/D vssd1 vssd1 vccd1 vccd1 _26271_/Q sky130_fd_sc_hd__dfxtp_2
X_23483_ _24870_/B _23432_/X _23482_/X vssd1 vssd1 vccd1 vccd1 _23484_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_119_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20695_ _21042_/A _20695_/B _20694_/X vssd1 vssd1 vccd1 vccd1 _20696_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_80_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25222_ _25678_/CLK hold484/X vssd1 vssd1 vccd1 vccd1 hold482/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22434_ _22431_/X _22432_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22434_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25153_ _26286_/CLK hold601/X vssd1 vssd1 vccd1 vccd1 hold599/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22365_ _22653_/A _22365_/B vssd1 vssd1 vccd1 vccd1 _22365_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_111_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _25991_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_115_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24104_ _24104_/A vssd1 vssd1 vccd1 vccd1 _26101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21316_ _21314_/Y _21315_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21316_/Y sky130_fd_sc_hd__a21oi_1
X_25084_ _26299_/CLK _25084_/D vssd1 vssd1 vccd1 vccd1 _25084_/Q sky130_fd_sc_hd__dfxtp_1
X_22296_ _22296_/A _25884_/Q vssd1 vssd1 vccd1 vccd1 _22296_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_130_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24035_ hold2389/X hold2286/X _24047_/S vssd1 vssd1 vccd1 vccd1 _24036_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_131_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21247_ _21678_/B _21630_/B vssd1 vssd1 vccd1 vccd1 _21249_/A sky130_fd_sc_hd__nand2_1
Xhold360 hold360/A vssd1 vssd1 vccd1 vccd1 hold360/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 hold371/A vssd1 vssd1 vccd1 vccd1 hold371/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold382 hold382/A vssd1 vssd1 vccd1 vccd1 hold382/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 hold393/A vssd1 vssd1 vccd1 vccd1 hold393/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21178_ _21636_/A _21178_/B _21177_/X vssd1 vssd1 vccd1 vccd1 _21179_/B sky130_fd_sc_hd__or3b_1
X_20129_ _20660_/A _20129_/B vssd1 vssd1 vccd1 vccd1 _20129_/Y sky130_fd_sc_hd__nand2_1
X_25986_ _25991_/CLK _25986_/D vssd1 vssd1 vccd1 vccd1 _25986_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24937_ _24946_/A _24937_/B vssd1 vssd1 vccd1 vccd1 _24937_/Y sky130_fd_sc_hd__nor2_1
X_12951_ _26252_/Q _25621_/Q vssd1 vssd1 vccd1 vccd1 _14413_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_172_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_178_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _26286_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1060 _20700_/Y vssd1 vssd1 vccd1 vccd1 _25791_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1071 _25126_/Q vssd1 vssd1 vccd1 vccd1 _19061_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15670_ _15670_/A vssd1 vssd1 vccd1 vccd1 _16585_/A sky130_fd_sc_hd__inv_2
Xhold1082 _13194_/X vssd1 vssd1 vccd1 vccd1 _25085_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24868_ _24859_/X _24867_/X _24949_/S vssd1 vssd1 vccd1 vccd1 _24868_/X sky130_fd_sc_hd__mux2_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1093 _25008_/Q vssd1 vssd1 vccd1 vccd1 _17109_/B sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ _12726_/B _14370_/A _12752_/X _25608_/Q vssd1 vssd1 vccd1 vccd1 _12882_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _14645_/A hold233/X vssd1 vssd1 vccd1 vccd1 hold234/A sky130_fd_sc_hd__nand2_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23819_ hold2105/X hold2032/X _23831_/S vssd1 vssd1 vccd1 vccd1 _23820_/A sky130_fd_sc_hd__mux2_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24799_ hold2722/X hold2714/X _24817_/S vssd1 vssd1 vccd1 vccd1 _24800_/A sky130_fd_sc_hd__mux2_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _19473_/A _17340_/B vssd1 vssd1 vccd1 vccd1 _17586_/A sky130_fd_sc_hd__xor2_4
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14585_/A hold98/X vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13503_ hold531/X _13502_/Y _12558_/B vssd1 vssd1 vccd1 vccd1 hold532/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17271_ _17271_/A _17444_/B vssd1 vssd1 vccd1 vccd1 _17271_/Y sky130_fd_sc_hd__nand2_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14483_ _14525_/A hold59/X vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__nand2_1
XFILLER_0_181_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19010_ _19010_/A _19080_/B vssd1 vssd1 vccd1 vccd1 _19011_/B sky130_fd_sc_hd__xnor2_1
X_16222_ _16224_/B _16224_/A vssd1 vssd1 vccd1 vccd1 _16223_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_153_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13434_ _13220_/A _14672_/A _13242_/A _25704_/Q vssd1 vssd1 vccd1 vccd1 _13434_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16153_ _16151_/X _16152_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _16153_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_102_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _25939_/CLK sky130_fd_sc_hd__clkbuf_16
X_13365_ _13365_/A vssd1 vssd1 vccd1 vccd1 _19701_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_183_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15104_ _15104_/A _15106_/B vssd1 vssd1 vccd1 vccd1 _15104_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16084_ _16084_/A _16084_/B vssd1 vssd1 vccd1 vccd1 _16104_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_11_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13296_ _26313_/Q _19546_/A vssd1 vssd1 vccd1 vccd1 _14605_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_146_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15035_ _15021_/A _14836_/Y _15016_/Y _15030_/B _15034_/Y vssd1 vssd1 vccd1 vccd1
+ _15035_/X sky130_fd_sc_hd__a221o_1
X_19912_ _19981_/A _19928_/B vssd1 vssd1 vccd1 vccd1 _19914_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19843_ _19840_/Y _19843_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19843_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_78_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19774_ _19774_/A _20518_/B vssd1 vssd1 vccd1 vccd1 _19774_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16986_ _25589_/Q vssd1 vssd1 vccd1 vccd1 _20285_/B sky130_fd_sc_hd__inv_2
X_18725_ _22436_/B _25634_/Q vssd1 vssd1 vccd1 vccd1 _18727_/A sky130_fd_sc_hd__nand2_1
X_15937_ _15935_/X _15936_/Y _15233_/X vssd1 vssd1 vccd1 vccd1 _15937_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_169_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _25793_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_155_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15868_ _15894_/A vssd1 vssd1 vccd1 vccd1 _15874_/B sky130_fd_sc_hd__inv_2
X_18656_ _18858_/A _18974_/A vssd1 vssd1 vccd1 vccd1 _18657_/B sky130_fd_sc_hd__xnor2_1
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14819_ _25851_/Q _12527_/A _15006_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14819_/X
+ sky130_fd_sc_hd__a22o_1
X_17607_ _17607_/A _17607_/B vssd1 vssd1 vccd1 vccd1 _17608_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15799_ _15799_/A _16974_/A vssd1 vssd1 vccd1 vccd1 _15800_/B sky130_fd_sc_hd__nor2_1
X_18587_ _18792_/A _18591_/B vssd1 vssd1 vccd1 vccd1 _18589_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_114_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17538_ _17538_/A _17582_/B vssd1 vssd1 vccd1 vccd1 _17538_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_175_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17469_ _17519_/A _17637_/B vssd1 vssd1 vccd1 vccd1 _17470_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19208_ _20467_/A _19206_/Y _20472_/C vssd1 vssd1 vccd1 vccd1 _19294_/B sky130_fd_sc_hd__o21a_4
X_20480_ _20483_/A _20483_/C vssd1 vssd1 vccd1 vccd1 _20481_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19139_ _19138_/C _17923_/B _20143_/A vssd1 vssd1 vccd1 vccd1 _19972_/B sky130_fd_sc_hd__a21boi_4
XFILLER_0_113_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22150_ _18512_/A _25815_/Q _22148_/Y _22149_/Y vssd1 vssd1 vccd1 vccd1 _22151_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21101_ _21101_/A _21844_/B vssd1 vssd1 vccd1 vccd1 _21102_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_140_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22081_ _22081_/A _22081_/B vssd1 vssd1 vccd1 vccd1 _22082_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21032_ _21500_/B _21548_/B vssd1 vssd1 vccd1 vccd1 _21033_/B sky130_fd_sc_hd__nand2_1
X_25840_ _25864_/CLK _25840_/D vssd1 vssd1 vccd1 vccd1 _25840_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_129_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25771_ _26275_/CLK _25771_/D vssd1 vssd1 vccd1 vccd1 _25771_/Q sky130_fd_sc_hd__dfxtp_1
X_22983_ _22982_/A _22849_/X _22982_/B vssd1 vssd1 vccd1 vccd1 _22984_/C sky130_fd_sc_hd__o21ai_1
X_24722_ hold2704/X hold2103/X _24740_/S vssd1 vssd1 vccd1 vccd1 _24723_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_97_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21934_ _21934_/A _22145_/B vssd1 vssd1 vccd1 vccd1 _21934_/Y sky130_fd_sc_hd__nand2_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24653_ _24653_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24654_/A sky130_fd_sc_hd__and2_1
XFILLER_0_179_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21865_ _21865_/A _22145_/B vssd1 vssd1 vccd1 vccd1 _21865_/Y sky130_fd_sc_hd__nand2_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23604_ input3/X hold2283/X _23677_/S vssd1 vssd1 vccd1 vccd1 _23605_/A sky130_fd_sc_hd__mux2_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20816_ _20814_/Y _20815_/Y _20465_/X vssd1 vssd1 vccd1 vccd1 _20816_/Y sky130_fd_sc_hd__a21oi_1
X_24584_ hold2701/X hold2575/X _24587_/S vssd1 vssd1 vccd1 vccd1 _24585_/A sky130_fd_sc_hd__mux2_1
X_21796_ _22653_/A _21796_/B vssd1 vssd1 vccd1 vccd1 _21796_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26323_ _26325_/CLK _26323_/D vssd1 vssd1 vccd1 vccd1 _26323_/Q sky130_fd_sc_hd__dfxtp_2
X_23535_ hold44/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23535_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_167_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20747_ _20747_/A _20747_/B vssd1 vssd1 vccd1 vccd1 _20749_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26254_ _26267_/CLK _26254_/D vssd1 vssd1 vccd1 vccd1 _26254_/Q sky130_fd_sc_hd__dfxtp_4
X_23466_ hold29/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23466_/X sky130_fd_sc_hd__or2b_1
X_20678_ _20681_/A _20681_/C vssd1 vssd1 vccd1 vccd1 _20680_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25205_ _25785_/CLK hold487/X vssd1 vssd1 vccd1 vccd1 hold485/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22417_ _22841_/A _22992_/B vssd1 vssd1 vccd1 vccd1 _22418_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26185_ _26190_/CLK _26185_/D vssd1 vssd1 vccd1 vccd1 _26185_/Q sky130_fd_sc_hd__dfxtp_1
X_23397_ _24942_/S hold257/A _23396_/X vssd1 vssd1 vccd1 vccd1 _23397_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13150_ _18270_/B _13320_/B vssd1 vssd1 vccd1 vccd1 _13150_/X sky130_fd_sc_hd__or2_1
X_25136_ _26122_/CLK hold741/X vssd1 vssd1 vccd1 vccd1 hold739/A sky130_fd_sc_hd__dfxtp_1
X_22348_ _25822_/Q _22348_/B vssd1 vssd1 vccd1 vccd1 _22348_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_27_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25067_ _26151_/CLK _25067_/D vssd1 vssd1 vccd1 vccd1 _25067_/Q sky130_fd_sc_hd__dfxtp_1
X_13081_ _13018_/X _13079_/X _13005_/X _13080_/X vssd1 vssd1 vccd1 vccd1 _13081_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22279_ _17816_/A _25791_/Q _22277_/Y _22278_/Y vssd1 vssd1 vccd1 vccd1 _22280_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_130_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24018_ _24018_/A _24096_/B vssd1 vssd1 vccd1 vccd1 _24019_/A sky130_fd_sc_hd__and2_1
XFILLER_0_104_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold190 hold190/A vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ _22848_/B _16773_/A _16836_/Y _16839_/Y _12702_/A vssd1 vssd1 vccd1 vccd1
+ _16840_/Y sky130_fd_sc_hd__a221oi_1
X_16771_ _16858_/A _16771_/B vssd1 vssd1 vccd1 vccd1 _16771_/Y sky130_fd_sc_hd__nand2_1
X_25969_ _26041_/CLK _25969_/D vssd1 vssd1 vccd1 vccd1 _25969_/Q sky130_fd_sc_hd__dfxtp_1
X_13983_ _17847_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13983_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_176_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15722_ _26039_/Q _25975_/Q _15809_/S vssd1 vssd1 vccd1 vccd1 _15723_/A sky130_fd_sc_hd__mux2_1
X_18510_ _18510_/A _18510_/B _18510_/C vssd1 vssd1 vccd1 vccd1 _22151_/A sky130_fd_sc_hd__nand3_2
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12934_ _17449_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12934_/X sky130_fd_sc_hd__or2_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ _21128_/A _19488_/Y _21132_/C vssd1 vssd1 vccd1 vccd1 _19579_/B sky130_fd_sc_hd__o21a_2
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15653_ _15654_/A _15655_/A vssd1 vssd1 vccd1 vccd1 _15657_/A sky130_fd_sc_hd__nor2_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18441_ _22065_/B _25620_/Q vssd1 vssd1 vccd1 vccd1 _18443_/A sky130_fd_sc_hd__nand2_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ _12840_/X _12863_/X _12827_/X _12864_/X vssd1 vssd1 vccd1 vccd1 _12865_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14604_ _14602_/Y hold45/X _14586_/X vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__a21oi_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18372_ _18372_/A _18372_/B vssd1 vssd1 vccd1 vccd1 _18372_/X sky130_fd_sc_hd__xor2_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15584_ _22979_/B _16369_/B vssd1 vssd1 vccd1 vccd1 _16520_/B sky130_fd_sc_hd__nand2_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _17148_/B _14264_/A vssd1 vssd1 vccd1 vccd1 _12796_/X sky130_fd_sc_hd__or2_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17323_ _17321_/X _17241_/X _17322_/X vssd1 vssd1 vccd1 vccd1 _17324_/A sky130_fd_sc_hd__a21o_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14535_ _14533_/Y hold105/X _14526_/X vssd1 vssd1 vccd1 vccd1 hold106/A sky130_fd_sc_hd__a21oi_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17254_ _17535_/A _17615_/A vssd1 vssd1 vccd1 vccd1 _17255_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_183_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14466_ _15464_/A vssd1 vssd1 vccd1 vccd1 _14466_/X sky130_fd_sc_hd__buf_8
X_16205_ _16205_/A hold912/X vssd1 vssd1 vccd1 vccd1 _16206_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13417_ _19026_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13417_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17185_ _17499_/A _17577_/A vssd1 vssd1 vccd1 vccd1 _17186_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14397_ _14397_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14397_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_141_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16136_ hold964/X vssd1 vssd1 vccd1 vccd1 _16139_/B sky130_fd_sc_hd__inv_2
X_13348_ _26321_/Q _19659_/A vssd1 vssd1 vccd1 vccd1 _14629_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_110_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16067_ _22262_/B _16401_/C vssd1 vssd1 vccd1 vccd1 _16069_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_122_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13279_ _13220_/X _14596_/A _13242_/X _19504_/A vssd1 vssd1 vccd1 vccd1 _13279_/X
+ sky130_fd_sc_hd__a22o_1
X_15018_ _15029_/A _15019_/A vssd1 vssd1 vccd1 vccd1 _15018_/X sky130_fd_sc_hd__or2_1
Xhold2508 _26325_/Q vssd1 vssd1 vccd1 vccd1 hold2508/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2519 _25904_/Q vssd1 vssd1 vccd1 vccd1 _17685_/A sky130_fd_sc_hd__buf_1
X_19826_ _26263_/Q _19134_/X hold847/X vssd1 vssd1 vccd1 vccd1 _19826_/Y sky130_fd_sc_hd__a21oi_1
Xhold1807 _22461_/Y vssd1 vssd1 vccd1 vccd1 _25862_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1818 _23211_/X vssd1 vssd1 vccd1 vccd1 _23212_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1829 _25622_/Q vssd1 vssd1 vccd1 vccd1 _17489_/B sky130_fd_sc_hd__dlygate4sd3_1
X_19757_ _19754_/Y _19757_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19757_/X sky130_fd_sc_hd__and3b_1
X_16969_ _16969_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16969_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_155_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18708_ _25889_/Q _22407_/A vssd1 vssd1 vccd1 vccd1 _18716_/A sky130_fd_sc_hd__or2_2
XFILLER_0_91_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19688_ _20272_/A _22297_/B _25628_/Q vssd1 vssd1 vccd1 vccd1 _20277_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_78_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18639_ _18637_/X _18269_/X _18638_/X vssd1 vssd1 vccd1 vccd1 _18640_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_177_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21650_ _26336_/Q hold632/X vssd1 vssd1 vccd1 vccd1 _21650_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20601_ _20601_/A _22493_/B _20601_/C vssd1 vssd1 vccd1 vccd1 _20605_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_117_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21581_ _21581_/A _21581_/B vssd1 vssd1 vccd1 vccd1 _21582_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23320_ _23320_/A _23320_/B vssd1 vssd1 vccd1 vccd1 _23320_/Y sky130_fd_sc_hd__nand2_1
X_20532_ _21302_/C _21578_/A vssd1 vssd1 vccd1 vccd1 _20534_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_89_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23251_ _23581_/B vssd1 vssd1 vccd1 vccd1 _23484_/B sky130_fd_sc_hd__inv_2
XFILLER_0_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20463_ _20463_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _20463_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_160_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22202_ _22200_/Y _22201_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _22202_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23182_ _23180_/X _23181_/Y _12702_/A vssd1 vssd1 vccd1 vccd1 _23182_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20394_ _20394_/A _22081_/B _20394_/C vssd1 vssd1 vccd1 vccd1 _20397_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_70_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22133_ _22133_/A _22133_/B vssd1 vssd1 vccd1 vccd1 _22133_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_101_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22064_ _22064_/A _25876_/Q vssd1 vssd1 vccd1 vccd1 _22064_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21015_ _21014_/Y _20192_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21015_/X
+ sky130_fd_sc_hd__a211o_1
X_25823_ _25838_/CLK _25823_/D vssd1 vssd1 vccd1 vccd1 _25823_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25754_ _25756_/CLK _25754_/D vssd1 vssd1 vccd1 vccd1 _25754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22966_ _22965_/A _22849_/X _22965_/B vssd1 vssd1 vccd1 vccd1 _22967_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_186_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24705_ _24705_/A _24741_/B vssd1 vssd1 vccd1 vccd1 _24706_/A sky130_fd_sc_hd__and2_1
XFILLER_0_179_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21917_ _22689_/B _21918_/A vssd1 vssd1 vccd1 vccd1 _21919_/A sky130_fd_sc_hd__or2_1
XFILLER_0_69_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25685_ _25687_/CLK _25685_/D vssd1 vssd1 vccd1 vccd1 _25685_/Q sky130_fd_sc_hd__dfxtp_1
X_22897_ _22896_/A _22454_/X _22896_/B vssd1 vssd1 vccd1 vccd1 _22898_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_168_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12650_ _12654_/B _12651_/A vssd1 vssd1 vccd1 vccd1 _12652_/A sky130_fd_sc_hd__or2_1
XFILLER_0_66_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24636_ hold2720/X hold2663/X _24664_/S vssd1 vssd1 vccd1 vccd1 _24637_/A sky130_fd_sc_hd__mux2_1
X_21848_ _22637_/B _21849_/A vssd1 vssd1 vccd1 vccd1 _21850_/A sky130_fd_sc_hd__or2_1
XFILLER_0_66_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12581_ _23377_/B vssd1 vssd1 vccd1 vccd1 _14910_/B sky130_fd_sc_hd__clkbuf_16
X_24567_ _24567_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24568_/A sky130_fd_sc_hd__and2_1
XFILLER_0_182_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21779_ _21779_/A _21779_/B vssd1 vssd1 vccd1 vccd1 _22575_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_33_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ _14344_/A hold188/X vssd1 vssd1 vccd1 vccd1 hold189/A sky130_fd_sc_hd__nand2_1
X_26306_ _26306_/CLK _26306_/D vssd1 vssd1 vccd1 vccd1 _26306_/Q sky130_fd_sc_hd__dfxtp_2
X_23518_ _23515_/Y _23517_/Y _24858_/S vssd1 vssd1 vccd1 vccd1 _23518_/X sky130_fd_sc_hd__mux2_1
X_24498_ hold2611/X hold2559/X _24510_/S vssd1 vssd1 vccd1 vccd1 _24499_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_92_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26237_ _26239_/CLK _26237_/D vssd1 vssd1 vccd1 vccd1 _26237_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_68_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14251_ _26338_/Q _13518_/B _14170_/X _14250_/Y vssd1 vssd1 vccd1 vccd1 _14252_/B
+ sky130_fd_sc_hd__a22o_1
X_23449_ _24922_/S hold299/A _23448_/X vssd1 vssd1 vccd1 vccd1 _23449_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13202_ _26298_/Q _19331_/A vssd1 vssd1 vccd1 vccd1 _14557_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14182_ _14236_/A hold823/X vssd1 vssd1 vccd1 vccd1 _14182_/Y sky130_fd_sc_hd__nand2_1
X_26168_ _26299_/CLK _26168_/D vssd1 vssd1 vccd1 vccd1 _26168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25119_ _26330_/CLK hold996/X vssd1 vssd1 vccd1 vccd1 hold995/A sky130_fd_sc_hd__dfxtp_1
X_13133_ _18208_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13133_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18990_ _19026_/A _18990_/B _22786_/A vssd1 vssd1 vccd1 vccd1 _18990_/X sky130_fd_sc_hd__and3_1
X_26099_ _26103_/CLK _26099_/D vssd1 vssd1 vccd1 vccd1 _26099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941_ _18612_/A _25723_/Q _18083_/C vssd1 vssd1 vccd1 vccd1 _17942_/C sky130_fd_sc_hd__nand3_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _13018_/X _13062_/X _13005_/X _13063_/X vssd1 vssd1 vccd1 vccd1 _13064_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17872_ _25840_/Q vssd1 vssd1 vccd1 vccd1 _20114_/A sky130_fd_sc_hd__inv_2
XFILLER_0_139_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19611_ _19609_/Y _19610_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19611_/Y sky130_fd_sc_hd__a21oi_1
X_16823_ _16824_/B _16824_/A vssd1 vssd1 vccd1 vccd1 _16823_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19542_ _26243_/Q _19483_/X hold629/X vssd1 vssd1 vccd1 vccd1 _19542_/Y sky130_fd_sc_hd__a21oi_1
X_16754_ _16754_/A _16754_/B vssd1 vssd1 vccd1 vccd1 _16754_/Y sky130_fd_sc_hd__nand2_1
X_13966_ _14061_/A _13966_/B vssd1 vssd1 vccd1 vccd1 _13966_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15705_ _26038_/Q _25974_/Q _15773_/S vssd1 vssd1 vccd1 vccd1 _15706_/A sky130_fd_sc_hd__mux2_1
X_12917_ _23377_/B vssd1 vssd1 vccd1 vccd1 _12917_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16685_ _16685_/A _16685_/B vssd1 vssd1 vccd1 vccd1 _16695_/A sky130_fd_sc_hd__nand2_1
X_19473_ _19473_/A _21102_/B vssd1 vssd1 vccd1 vccd1 _19473_/Y sky130_fd_sc_hd__nor2_1
X_13897_ _26281_/Q _13801_/X _13793_/X _13896_/Y vssd1 vssd1 vccd1 vccd1 _13898_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18424_ _25875_/Q _22039_/A vssd1 vssd1 vccd1 vccd1 _18432_/A sky130_fd_sc_hd__or2_2
X_15636_ _23028_/B _15812_/B vssd1 vssd1 vccd1 vccd1 _15637_/A sky130_fd_sc_hd__nand2_1
X_12848_ _26104_/Q _12748_/X _12847_/X vssd1 vssd1 vccd1 vccd1 _12848_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15567_ _22962_/B _15812_/B vssd1 vssd1 vccd1 vccd1 _15568_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18355_ _18355_/A _18579_/B vssd1 vssd1 vccd1 vccd1 _18355_/Y sky130_fd_sc_hd__nand2_1
X_12779_ _12726_/B _14307_/A _12752_/X _25588_/Q vssd1 vssd1 vccd1 vccd1 _12779_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17306_ _25708_/Q _17306_/B vssd1 vssd1 vccd1 vccd1 _17644_/A sky130_fd_sc_hd__xor2_4
X_14518_ _14518_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14518_/Y sky130_fd_sc_hd__nand2_1
X_15498_ _15470_/X _15502_/B _15481_/B vssd1 vssd1 vccd1 vccd1 _15500_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18286_ _18529_/A vssd1 vssd1 vccd1 vccd1 _18952_/A sky130_fd_sc_hd__buf_8
XFILLER_0_142_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17237_ _19844_/A _17237_/B vssd1 vssd1 vccd1 vccd1 _17607_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_47_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14449_ _14449_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _14449_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_114_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold904 hold904/A vssd1 vssd1 vccd1 vccd1 hold904/X sky130_fd_sc_hd__dlygate4sd3_1
X_17168_ _19289_/A _17168_/B vssd1 vssd1 vccd1 vccd1 _17492_/A sky130_fd_sc_hd__xor2_4
Xhold915 hold915/A vssd1 vssd1 vccd1 vccd1 hold915/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold926 hold926/A vssd1 vssd1 vccd1 vccd1 hold926/X sky130_fd_sc_hd__dlygate4sd3_1
X_16119_ _16117_/X hold429/X _16076_/X vssd1 vssd1 vccd1 vccd1 hold430/A sky130_fd_sc_hd__a21oi_1
Xhold937 hold937/A vssd1 vssd1 vccd1 vccd1 hold937/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 hold948/A vssd1 vssd1 vccd1 vccd1 hold948/X sky130_fd_sc_hd__buf_1
XFILLER_0_122_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold959 hold959/A vssd1 vssd1 vccd1 vccd1 hold959/X sky130_fd_sc_hd__dlygate4sd3_1
X_17099_ _20248_/B _25844_/Q _25780_/Q vssd1 vssd1 vccd1 vccd1 _17100_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_110_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2305 _15073_/Y vssd1 vssd1 vccd1 vccd1 hold2305/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2316 _12660_/Y vssd1 vssd1 vccd1 vccd1 _12662_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2327 _24047_/X vssd1 vssd1 vccd1 vccd1 _24048_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2338 _14952_/Y vssd1 vssd1 vccd1 vccd1 hold2338/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1604 _25604_/Q vssd1 vssd1 vccd1 vccd1 _17325_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2349 _25675_/Q vssd1 vssd1 vccd1 vccd1 _13253_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1615 _17418_/Y vssd1 vssd1 vccd1 vccd1 _25613_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1626 _25889_/Q vssd1 vssd1 vccd1 vccd1 _23005_/B sky130_fd_sc_hd__buf_1
X_19809_ _19801_/X _19808_/Y _19766_/X vssd1 vssd1 vccd1 vccd1 _19809_/Y sky130_fd_sc_hd__o21ai_1
Xhold1637 _25640_/Q vssd1 vssd1 vccd1 vccd1 _17620_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1648 _17918_/Y vssd1 vssd1 vccd1 vccd1 _25648_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1659 _25829_/Q vssd1 vssd1 vccd1 vccd1 _21590_/B sky130_fd_sc_hd__dlygate4sd3_1
X_22820_ _22811_/Y _22819_/Y _22534_/X vssd1 vssd1 vccd1 vccd1 _22820_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22751_ _22750_/A _22454_/X _22750_/B vssd1 vssd1 vccd1 vccd1 _22752_/C sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_91_clk clkbuf_leaf_95_clk/A vssd1 vssd1 vccd1 vccd1 _26341_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21702_ _21702_/A _22902_/B vssd1 vssd1 vccd1 vccd1 _21702_/Y sky130_fd_sc_hd__nand2_1
X_25470_ _25532_/CLK hold884/X vssd1 vssd1 vccd1 vccd1 hold883/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22682_ _26054_/Q vssd1 vssd1 vccd1 vccd1 _22683_/A sky130_fd_sc_hd__inv_2
XFILLER_0_176_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24421_ hold2328/X hold2214/X _24433_/S vssd1 vssd1 vccd1 vccd1 _24422_/A sky130_fd_sc_hd__mux2_1
X_21633_ _26335_/Q _19130_/X hold383/X vssd1 vssd1 vccd1 vccd1 _21636_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24352_ _24352_/A vssd1 vssd1 vccd1 vccd1 _26182_/D sky130_fd_sc_hd__clkbuf_1
X_21564_ _21564_/A _21564_/B _21564_/C vssd1 vssd1 vccd1 vccd1 _21565_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23303_ _23303_/A _23303_/B vssd1 vssd1 vccd1 vccd1 _23303_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_160_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20515_ _20515_/A _20515_/B vssd1 vssd1 vccd1 vccd1 _21305_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24283_ hold2309/X hold1909/X _24356_/S vssd1 vssd1 vccd1 vccd1 _24285_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_132_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21495_ _21546_/A _21499_/A vssd1 vssd1 vccd1 vccd1 _21497_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_160_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26022_ _26023_/CLK _26022_/D vssd1 vssd1 vccd1 vccd1 _26022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23234_ _23234_/A _24836_/B _23238_/A vssd1 vssd1 vccd1 vccd1 _23235_/A sky130_fd_sc_hd__and3_1
X_20446_ _20446_/A _20446_/B vssd1 vssd1 vccd1 vccd1 _20448_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23165_ _23197_/A _23165_/B vssd1 vssd1 vccd1 vccd1 _23165_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_141_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20377_ _21195_/C _21515_/A vssd1 vssd1 vccd1 vccd1 _20378_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_113_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22116_ _22116_/A _22145_/B vssd1 vssd1 vccd1 vccd1 _22116_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23096_ _23095_/A _22849_/X _23095_/B vssd1 vssd1 vccd1 vccd1 _23097_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22047_ _22758_/B vssd1 vssd1 vccd1 vccd1 _22759_/A sky130_fd_sc_hd__inv_2
X_13820_ _25766_/Q vssd1 vssd1 vccd1 vccd1 _18813_/B sky130_fd_sc_hd__inv_2
X_25806_ _25807_/CLK _25806_/D vssd1 vssd1 vccd1 vccd1 _25806_/Q sky130_fd_sc_hd__dfxtp_1
X_23998_ _26067_/Q hold2437/X _24001_/S vssd1 vssd1 vccd1 vccd1 _23998_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_187_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25737_ _25740_/CLK _25737_/D vssd1 vssd1 vccd1 vccd1 _25737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13751_ _26258_/Q _13612_/X _13605_/X _13750_/Y vssd1 vssd1 vccd1 vccd1 _13752_/B
+ sky130_fd_sc_hd__a22o_1
X_22949_ _22948_/A _22849_/X _22948_/B vssd1 vssd1 vccd1 vccd1 _22950_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_82_clk clkbuf_leaf_82_clk/A vssd1 vssd1 vccd1 vccd1 _26004_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12702_ _12702_/A _12702_/B vssd1 vssd1 vccd1 vccd1 _12702_/Y sky130_fd_sc_hd__nor2_1
X_16470_ _16470_/A _16470_/B vssd1 vssd1 vccd1 vccd1 _16480_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_39_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25668_ _26302_/CLK _25668_/D vssd1 vssd1 vccd1 vccd1 _25668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13682_ _25744_/Q vssd1 vssd1 vccd1 vccd1 _18367_/B sky130_fd_sc_hd__inv_2
X_15421_ _22828_/B _15776_/B vssd1 vssd1 vccd1 vccd1 _15422_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_128_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12633_ _12635_/B _12635_/A vssd1 vssd1 vccd1 vccd1 _12654_/A sky130_fd_sc_hd__nor2_1
X_24619_ _24619_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24620_/A sky130_fd_sc_hd__and2_1
X_25599_ _26109_/CLK _25599_/D vssd1 vssd1 vccd1 vccd1 _25599_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15352_ _22763_/B _16369_/B vssd1 vssd1 vccd1 vccd1 _15353_/A sky130_fd_sc_hd__nand2_1
X_18140_ _20915_/B _21906_/A vssd1 vssd1 vccd1 vccd1 _20908_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_183_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12564_ _12564_/A _23597_/C vssd1 vssd1 vccd1 vccd1 _12565_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_109_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14303_ _14301_/Y hold237/X _14280_/X vssd1 vssd1 vccd1 vccd1 hold238/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18071_ _18071_/A _25716_/Q _18118_/A vssd1 vssd1 vccd1 vccd1 _18074_/C sky130_fd_sc_hd__nand3_2
X_15283_ _26014_/Q _25950_/Q _15773_/S vssd1 vssd1 vccd1 vccd1 _15284_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_108_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12495_ input7/X vssd1 vssd1 vccd1 vccd1 _14345_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17022_ _20310_/B _25846_/Q _25782_/Q vssd1 vssd1 vccd1 vccd1 _17023_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_34_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14234_ _14264_/A _14234_/B vssd1 vssd1 vccd1 vccd1 _14234_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_151_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14165_ _18633_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _14165_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13116_ _13049_/X _14509_/A _13067_/X _25652_/Q vssd1 vssd1 vccd1 vccd1 _13116_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _18409_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14096_/Y sky130_fd_sc_hd__nor2_1
X_18973_ _18971_/Y _18972_/Y _18924_/X vssd1 vssd1 vccd1 vccd1 _25693_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _17609_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13047_/X sky130_fd_sc_hd__or2_1
X_17924_ _17924_/A _17924_/B vssd1 vssd1 vccd1 vccd1 _17925_/A sky130_fd_sc_hd__or2_1
X_17855_ _18612_/A _25721_/Q _18083_/C vssd1 vssd1 vccd1 vccd1 _17856_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_79_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16806_ _16858_/A _16806_/B vssd1 vssd1 vccd1 vccd1 _16806_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17786_ _18118_/A _18153_/B _18118_/B vssd1 vssd1 vccd1 vccd1 _18122_/C sky130_fd_sc_hd__nand3_4
XFILLER_0_178_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14998_ _14998_/A _14998_/B vssd1 vssd1 vccd1 vccd1 _15032_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_152_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19525_ _19517_/X _19524_/Y _19496_/X vssd1 vssd1 vccd1 vccd1 _19525_/Y sky130_fd_sc_hd__o21ai_1
X_16737_ _16735_/Y _16736_/Y _16594_/X vssd1 vssd1 vccd1 vccd1 _16737_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13949_ hold743/X _13948_/Y _13917_/X vssd1 vssd1 vccd1 vccd1 hold744/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_163_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_73_clk _25759_/CLK vssd1 vssd1 vccd1 vccd1 _25883_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19456_ _19455_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19457_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_186_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16668_ _16668_/A _16668_/B vssd1 vssd1 vccd1 vccd1 _16680_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18407_ _18529_/C vssd1 vssd1 vccd1 vccd1 _18894_/C sky130_fd_sc_hd__buf_6
X_15619_ _23015_/B _15619_/B vssd1 vssd1 vccd1 vccd1 _23012_/B sky130_fd_sc_hd__xor2_1
X_19387_ _19384_/Y _19387_/B _19980_/B vssd1 vssd1 vccd1 vccd1 _19387_/X sky130_fd_sc_hd__and3b_1
X_16599_ _16599_/A _16599_/B vssd1 vssd1 vccd1 vccd1 _16602_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18338_ _19504_/A vssd1 vssd1 vccd1 vccd1 _21913_/B sky130_fd_sc_hd__inv_2
XFILLER_0_127_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18269_ _22704_/A vssd1 vssd1 vccd1 vccd1 _18269_/X sky130_fd_sc_hd__buf_8
XFILLER_0_4_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20300_ _20300_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20305_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_142_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21280_ _21280_/A _21280_/B vssd1 vssd1 vccd1 vccd1 _21281_/A sky130_fd_sc_hd__nand2_1
Xhold701 hold701/A vssd1 vssd1 vccd1 vccd1 hold701/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 hold712/A vssd1 vssd1 vccd1 vccd1 hold712/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold723 hold723/A vssd1 vssd1 vccd1 vccd1 hold723/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20231_ _20231_/A _20231_/B vssd1 vssd1 vccd1 vccd1 _20232_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold734 hold734/A vssd1 vssd1 vccd1 vccd1 hold734/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 hold745/A vssd1 vssd1 vccd1 vccd1 hold745/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 hold756/A vssd1 vssd1 vccd1 vccd1 hold756/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 hold767/A vssd1 vssd1 vccd1 vccd1 hold767/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 hold778/A vssd1 vssd1 vccd1 vccd1 hold778/X sky130_fd_sc_hd__dlygate4sd3_1
X_20162_ _20162_/A _22208_/B vssd1 vssd1 vccd1 vccd1 _20163_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_110_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold789 hold789/A vssd1 vssd1 vccd1 vccd1 hold789/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2102 _23625_/X vssd1 vssd1 vccd1 vccd1 _23626_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2113 _23323_/X vssd1 vssd1 vccd1 vccd1 _23325_/A sky130_fd_sc_hd__dlygate4sd3_1
X_24970_ _25420_/CLK _24970_/D vssd1 vssd1 vccd1 vccd1 _24970_/Q sky130_fd_sc_hd__dfxtp_1
X_20093_ _20095_/B _20095_/C vssd1 vssd1 vccd1 vccd1 _20094_/A sky130_fd_sc_hd__nand2_1
Xhold2124 _26101_/Q vssd1 vssd1 vccd1 vccd1 hold2124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2135 _26111_/Q vssd1 vssd1 vccd1 vccd1 hold2135/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1401 _25103_/Q vssd1 vssd1 vccd1 vccd1 _18779_/B sky130_fd_sc_hd__dlygate4sd3_1
X_23921_ _23921_/A _24002_/B vssd1 vssd1 vccd1 vccd1 _23922_/A sky130_fd_sc_hd__and2_1
Xhold2146 _24123_/X vssd1 vssd1 vccd1 vccd1 _24124_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1412 _16845_/Y vssd1 vssd1 vccd1 vccd1 _25560_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2157 _26125_/Q vssd1 vssd1 vccd1 vccd1 hold2157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2168 _25932_/Q vssd1 vssd1 vccd1 vccd1 _23345_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1423 _25076_/Q vssd1 vssd1 vccd1 vccd1 _18229_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2179 _23983_/X vssd1 vssd1 vccd1 vccd1 _23984_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 _13314_/X vssd1 vssd1 vccd1 vccd1 _25104_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1445 _25770_/Q vssd1 vssd1 vccd1 vccd1 _19964_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1456 _14796_/Y vssd1 vssd1 vccd1 vccd1 _25399_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23852_ _23852_/A vssd1 vssd1 vccd1 vccd1 _26021_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1467 _25400_/Q vssd1 vssd1 vccd1 vccd1 _14804_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1478 _14704_/Y vssd1 vssd1 vccd1 vccd1 _25389_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1489 _25755_/Q vssd1 vssd1 vccd1 vccd1 _19768_/B sky130_fd_sc_hd__dlygate4sd3_1
X_22803_ _22803_/A _23099_/B vssd1 vssd1 vccd1 vccd1 _22803_/Y sky130_fd_sc_hd__nand2_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23783_ _23783_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23784_/A sky130_fd_sc_hd__and2_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20995_ _20998_/A _20998_/C vssd1 vssd1 vccd1 vccd1 _20996_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_64_clk _25472_/CLK vssd1 vssd1 vccd1 vccd1 _25450_/CLK sky130_fd_sc_hd__clkbuf_16
X_25522_ _25534_/CLK hold971/X vssd1 vssd1 vccd1 vccd1 hold970/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22734_ _22734_/A _22734_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22736_/A sky130_fd_sc_hd__or3_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25453_ _26057_/CLK _25453_/D vssd1 vssd1 vccd1 vccd1 _25453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22665_ _25835_/Q _22665_/B vssd1 vssd1 vccd1 vccd1 _22665_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_153_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24404_ _24404_/A _24465_/B vssd1 vssd1 vccd1 vccd1 _24405_/A sky130_fd_sc_hd__and2_1
XFILLER_0_34_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21616_ _21616_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _21621_/A sky130_fd_sc_hd__nand2_1
X_25384_ _26207_/CLK hold232/X vssd1 vssd1 vccd1 vccd1 hold230/A sky130_fd_sc_hd__dfxtp_1
X_22596_ _22596_/A _22596_/B vssd1 vssd1 vccd1 vccd1 _23104_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24335_ hold2412/X hold2404/X _24356_/S vssd1 vssd1 vccd1 vccd1 _24336_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_63_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21547_ _21547_/A _21596_/A vssd1 vssd1 vccd1 vccd1 _21548_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_16_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24266_ _24266_/A vssd1 vssd1 vccd1 vccd1 _26154_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21478_ _21481_/A _21531_/A vssd1 vssd1 vccd1 vccd1 _21480_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_133_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26005_ _26073_/CLK _26005_/D vssd1 vssd1 vccd1 vccd1 _26005_/Q sky130_fd_sc_hd__dfxtp_1
X_23217_ _24945_/S vssd1 vssd1 vccd1 vccd1 _24956_/S sky130_fd_sc_hd__buf_12
XFILLER_0_160_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20429_ _20429_/A _20429_/B vssd1 vssd1 vccd1 vccd1 _20432_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24197_ hold1831/X hold2110/X _24203_/S vssd1 vssd1 vccd1 vccd1 _24198_/A sky130_fd_sc_hd__mux2_1
X_23148_ _23139_/Y _23147_/Y _19199_/A vssd1 vssd1 vccd1 vccd1 _23148_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15970_ _15971_/B _15971_/A vssd1 vssd1 vccd1 vccd1 _15987_/B sky130_fd_sc_hd__or2_1
X_23079_ _23079_/A _23079_/B _23191_/C vssd1 vssd1 vccd1 vccd1 _23081_/A sky130_fd_sc_hd__or3_1
XFILLER_0_101_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14921_ _14921_/A vssd1 vssd1 vccd1 vccd1 _25414_/D sky130_fd_sc_hd__inv_2
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2680 _25475_/Q vssd1 vssd1 vccd1 vccd1 _15807_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
X_17640_ _17638_/X _17528_/X _17639_/X vssd1 vssd1 vccd1 vccd1 _17641_/A sky130_fd_sc_hd__a21o_1
X_14852_ _14852_/A _22263_/A vssd1 vssd1 vccd1 vccd1 _22262_/B sky130_fd_sc_hd__xnor2_2
Xhold2691 _26326_/Q vssd1 vssd1 vccd1 vccd1 hold2691/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1990 _24415_/X vssd1 vssd1 vccd1 vccd1 _24416_/A sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ _18753_/B _13876_/B vssd1 vssd1 vccd1 vccd1 _13803_/Y sky130_fd_sc_hd__nor2_1
X_14783_ _25847_/Q _12527_/A _14972_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14783_/X
+ sky130_fd_sc_hd__a22o_1
X_17571_ _17571_/A _17571_/B vssd1 vssd1 vccd1 vccd1 _17571_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_187_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_55_clk _25472_/CLK vssd1 vssd1 vccd1 vccd1 _26064_/CLK sky130_fd_sc_hd__clkbuf_16
X_19310_ _19302_/X _19309_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19310_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16522_ _16522_/A _16522_/B vssd1 vssd1 vccd1 vccd1 _16523_/B sky130_fd_sc_hd__nand2_1
X_13734_ _13823_/A _13734_/B vssd1 vssd1 vccd1 vccd1 _13734_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19241_ _19241_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _19241_/Y sky130_fd_sc_hd__nand2_1
X_16453_ _16461_/B vssd1 vssd1 vccd1 vccd1 _16456_/B sky130_fd_sc_hd__inv_2
XFILLER_0_151_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13665_ _26244_/Q _13612_/X _13605_/X _13664_/Y vssd1 vssd1 vccd1 vccd1 _13666_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _15404_/A _15403_/Y vssd1 vssd1 vccd1 vccd1 _15443_/A sky130_fd_sc_hd__or2b_1
XFILLER_0_156_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12616_ _12616_/A vssd1 vssd1 vccd1 vccd1 _12618_/B sky130_fd_sc_hd__inv_2
X_16384_ _16362_/X _16379_/A _16383_/Y vssd1 vssd1 vccd1 vccd1 _16384_/X sky130_fd_sc_hd__a21o_1
X_19172_ _26217_/Q hold766/X vssd1 vssd1 vccd1 vccd1 _19172_/Y sky130_fd_sc_hd__nand2_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _13703_/A _13596_/B vssd1 vssd1 vccd1 vccd1 _13596_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15335_ _22750_/B _15335_/B vssd1 vssd1 vccd1 vccd1 _22747_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_137_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18123_ _18125_/A _18125_/B vssd1 vssd1 vccd1 vccd1 _18124_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12547_ _13220_/A _21203_/A vssd1 vssd1 vccd1 vccd1 _13465_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_42_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15266_ _15266_/A _15266_/B vssd1 vssd1 vccd1 vccd1 _15267_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_152_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18054_ _20862_/B _21837_/A vssd1 vssd1 vccd1 vccd1 _20855_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_83_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_3 _20158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14217_ hold752/X _14216_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold753/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17005_ _22786_/A vssd1 vssd1 vccd1 vccd1 _19994_/B sky130_fd_sc_hd__buf_8
X_15197_ _15197_/A vssd1 vssd1 vccd1 vccd1 _16740_/A sky130_fd_sc_hd__inv_2
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14148_ _14180_/A _14148_/B vssd1 vssd1 vccd1 vccd1 _14148_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18956_ _18956_/A _18956_/B _18956_/C vssd1 vssd1 vccd1 vccd1 _22720_/A sky130_fd_sc_hd__nand3_2
X_14079_ _26310_/Q _13988_/X _13981_/X _14078_/Y vssd1 vssd1 vccd1 vccd1 _14080_/B
+ sky130_fd_sc_hd__a22o_1
X_17907_ _18528_/A _25729_/Q vssd1 vssd1 vccd1 vccd1 _17909_/A sky130_fd_sc_hd__nand2_1
X_18887_ _25642_/Q _22640_/B vssd1 vssd1 vccd1 vccd1 _18888_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_179_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17838_ _22308_/B _25600_/Q vssd1 vssd1 vccd1 vccd1 _17840_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17769_ _17771_/B vssd1 vssd1 vccd1 vccd1 _17783_/C sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_46_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _26023_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19508_ _19509_/B _19509_/A vssd1 vssd1 vccd1 vccd1 _19508_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20780_ _20780_/A _20780_/B vssd1 vssd1 vccd1 vccd1 _20784_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_147_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19439_ _19437_/Y _19438_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19439_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22450_ _15116_/B _22387_/B _14273_/X vssd1 vssd1 vccd1 vccd1 _22450_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21401_ _21401_/A _21449_/A vssd1 vssd1 vccd1 vccd1 _21403_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22381_ _22381_/A _23087_/A _22381_/C vssd1 vssd1 vccd1 vccd1 _22381_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_127_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24120_ hold2451/X hold2145/X _24126_/S vssd1 vssd1 vccd1 vccd1 _24121_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_60_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21332_ _21330_/Y _21331_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21332_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24051_ _24743_/A vssd1 vssd1 vccd1 vccd1 _24835_/S sky130_fd_sc_hd__clkbuf_16
Xhold520 hold520/A vssd1 vssd1 vccd1 vccd1 hold520/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21263_ _21260_/Y _21262_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21263_/Y sky130_fd_sc_hd__a21oi_1
Xhold531 hold531/A vssd1 vssd1 vccd1 vccd1 hold531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 hold542/A vssd1 vssd1 vccd1 vccd1 hold542/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_23002_ _16900_/B _22421_/X _22996_/X _22997_/Y _23001_/X vssd1 vssd1 vccd1 vccd1
+ _23003_/A sky130_fd_sc_hd__a221o_1
Xhold553 hold553/A vssd1 vssd1 vccd1 vccd1 hold553/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20214_ _20214_/A _20214_/B _20214_/C vssd1 vssd1 vccd1 vccd1 _20217_/C sky130_fd_sc_hd__nand3_1
Xhold564 hold564/A vssd1 vssd1 vccd1 vccd1 hold564/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 hold575/A vssd1 vssd1 vccd1 vccd1 hold575/X sky130_fd_sc_hd__dlygate4sd3_1
X_21194_ _21597_/B _21643_/C vssd1 vssd1 vccd1 vccd1 _21195_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold586 hold586/A vssd1 vssd1 vccd1 vccd1 hold586/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold597 hold597/A vssd1 vssd1 vccd1 vccd1 hold597/X sky130_fd_sc_hd__dlygate4sd3_1
X_20145_ _20145_/A _20145_/B vssd1 vssd1 vccd1 vccd1 _21033_/C sky130_fd_sc_hd__xor2_4
XFILLER_0_110_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24953_ _24956_/S hold871/X _24946_/A _24952_/Y vssd1 vssd1 vccd1 vccd1 _24953_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20076_ _20076_/A _20076_/B vssd1 vssd1 vccd1 vccd1 _20077_/A sky130_fd_sc_hd__nand2_1
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1220 _19724_/Y vssd1 vssd1 vccd1 vccd1 _25752_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1231 _20778_/Y vssd1 vssd1 vccd1 vccd1 _25793_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1242 _25576_/Q vssd1 vssd1 vccd1 vccd1 _16956_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_23904_ hold1963/X _26039_/Q _23907_/S vssd1 vssd1 vccd1 vccd1 _23904_/X sky130_fd_sc_hd__mux2_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24884_ _16113_/B _16123_/B _24956_/S vssd1 vssd1 vccd1 vccd1 _24885_/A sky130_fd_sc_hd__mux2_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1253 _13206_/X vssd1 vssd1 vccd1 vccd1 _25087_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1264 _25397_/Q vssd1 vssd1 vccd1 vccd1 _14777_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1275 _16730_/Y vssd1 vssd1 vccd1 vccd1 _25543_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23835_ hold2120/X _26016_/Q _23907_/S vssd1 vssd1 vccd1 vccd1 _23835_/X sky130_fd_sc_hd__mux2_1
Xhold1286 _25405_/Q vssd1 vssd1 vccd1 vccd1 _14844_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1297 _20816_/Y vssd1 vssd1 vccd1 vccd1 _25794_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_37_clk _25184_/CLK vssd1 vssd1 vccd1 vccd1 _26273_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23766_ _23766_/A vssd1 vssd1 vccd1 vccd1 _25993_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20978_ _20978_/A _20978_/B _20978_/C vssd1 vssd1 vccd1 vccd1 _20982_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25505_ _25510_/CLK _25505_/D vssd1 vssd1 vccd1 vccd1 hold972/A sky130_fd_sc_hd__dfxtp_1
X_22717_ _22717_/A _25901_/Q vssd1 vssd1 vccd1 vccd1 _22717_/Y sky130_fd_sc_hd__nand2_1
X_23697_ _23697_/A _23721_/B vssd1 vssd1 vccd1 vccd1 _23698_/A sky130_fd_sc_hd__and2_1
XFILLER_0_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25436_ _25501_/CLK hold932/X vssd1 vssd1 vccd1 vccd1 hold931/A sky130_fd_sc_hd__dfxtp_1
X_13450_ _26210_/Q _13426_/X _13449_/X vssd1 vssd1 vccd1 vccd1 _13450_/X sky130_fd_sc_hd__a21o_1
X_22648_ _23135_/B _22992_/B vssd1 vssd1 vccd1 vccd1 _22650_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13381_ _18983_/B _13944_/A vssd1 vssd1 vccd1 vccd1 _13381_/X sky130_fd_sc_hd__or2_1
X_25367_ _26190_/CLK hold472/X vssd1 vssd1 vccd1 vccd1 hold470/A sky130_fd_sc_hd__dfxtp_1
X_22579_ _26050_/Q vssd1 vssd1 vccd1 vccd1 _22580_/A sky130_fd_sc_hd__inv_2
XFILLER_0_180_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15120_ hold931/X _15122_/A vssd1 vssd1 vccd1 vccd1 _15124_/A sky130_fd_sc_hd__nor2_1
X_24318_ _24318_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24319_/A sky130_fd_sc_hd__and2_1
XFILLER_0_161_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25298_ _26249_/CLK hold331/X vssd1 vssd1 vccd1 vccd1 hold329/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15051_ _15051_/A _15051_/B vssd1 vssd1 vccd1 vccd1 _15068_/B sky130_fd_sc_hd__nor2_1
X_24249_ hold2153/X _26149_/Q _24279_/S vssd1 vssd1 vccd1 vccd1 _24249_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14002_ _14120_/A vssd1 vssd1 vccd1 vccd1 _14114_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18810_ _18952_/A _25766_/Q _18891_/C vssd1 vssd1 vccd1 vccd1 _18811_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_101_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19790_ _20557_/A _19788_/Y _20562_/C vssd1 vssd1 vccd1 vccd1 _19875_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18741_ _18741_/A _18963_/B vssd1 vssd1 vccd1 vccd1 _18741_/Y sky130_fd_sc_hd__nand2_1
X_15953_ _16000_/B _15953_/B vssd1 vssd1 vccd1 vccd1 _15961_/A sky130_fd_sc_hd__or2_1
X_14904_ _14904_/A vssd1 vssd1 vccd1 vccd1 _14909_/B sky130_fd_sc_hd__inv_2
X_18672_ _18792_/A _19824_/B vssd1 vssd1 vccd1 vccd1 _18674_/A sky130_fd_sc_hd__nand2_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ _15894_/B _15884_/B _15884_/C vssd1 vssd1 vccd1 vccd1 _15884_/Y sky130_fd_sc_hd__nand3b_1
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17623_ _17623_/A _17623_/B vssd1 vssd1 vccd1 vccd1 _17623_/X sky130_fd_sc_hd__xor2_1
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14835_ _22203_/B _15778_/B vssd1 vssd1 vccd1 vccd1 _15021_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_clk _25759_/CLK vssd1 vssd1 vccd1 vccd1 _25773_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _17552_/Y _17553_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _17554_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14766_ _25845_/Q _13466_/A _14765_/X _14270_/A vssd1 vssd1 vccd1 vccd1 _14767_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16505_ _16503_/B _16524_/A _16504_/Y vssd1 vssd1 vccd1 vccd1 _16505_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13717_ hold543/X _13716_/Y _13679_/X vssd1 vssd1 vccd1 vccd1 hold544/A sky130_fd_sc_hd__a21oi_1
X_14697_ _25838_/Q _12527_/A _14903_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14697_/X
+ sky130_fd_sc_hd__a22o_1
X_17485_ _17485_/A _17485_/B vssd1 vssd1 vccd1 vccd1 _17485_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_160_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19224_ _26220_/Q _19483_/A hold768/X vssd1 vssd1 vccd1 vccd1 _19225_/C sky130_fd_sc_hd__a21o_1
X_16436_ _16437_/B _16437_/A vssd1 vssd1 vccd1 vccd1 _16438_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_144_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13648_ hold597/X _13647_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold598/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_183_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ _22786_/A vssd1 vssd1 vccd1 vccd1 _19980_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16367_ _16473_/A hold950/X vssd1 vssd1 vccd1 vccd1 _16367_/Y sky130_fd_sc_hd__nand2_1
X_13579_ _13642_/A hold464/X vssd1 vssd1 vccd1 vccd1 hold465/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18106_ _19060_/A _18106_/B vssd1 vssd1 vccd1 vccd1 _18106_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_87_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15318_ _22731_/B _16369_/B _15778_/B vssd1 vssd1 vccd1 vccd1 _16787_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_26_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16298_ _16309_/B _16299_/A vssd1 vssd1 vccd1 vccd1 _16298_/X sky130_fd_sc_hd__or2_1
X_19086_ _21099_/A vssd1 vssd1 vccd1 vccd1 _19086_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_152_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18037_ _18037_/A _20585_/A vssd1 vssd1 vccd1 vccd1 _19073_/A sky130_fd_sc_hd__xor2_4
X_15249_ _15266_/A vssd1 vssd1 vccd1 vccd1 _15252_/B sky130_fd_sc_hd__inv_2
XFILLER_0_169_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19988_ _19985_/Y _19987_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _19988_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18939_ _19024_/A _19073_/B vssd1 vssd1 vccd1 vccd1 _18940_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21950_ _19518_/A _21949_/A _21949_/Y vssd1 vssd1 vccd1 vccd1 _21952_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20901_ _26300_/Q hold503/X vssd1 vssd1 vccd1 vccd1 _20901_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_55_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21881_ _19488_/A _21880_/A _21880_/Y vssd1 vssd1 vccd1 vccd1 _21883_/A sky130_fd_sc_hd__o21ai_2
Xclkbuf_leaf_19_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _26152_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23620_ _23620_/A _23629_/B vssd1 vssd1 vccd1 vccd1 _23621_/A sky130_fd_sc_hd__and2_1
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20832_ _23149_/B vssd1 vssd1 vccd1 vccd1 _22645_/B sky130_fd_sc_hd__inv_2
XFILLER_0_166_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23551_ hold143/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23551_/X sky130_fd_sc_hd__or2b_1
X_20763_ _21676_/B _21403_/B vssd1 vssd1 vccd1 vccd1 _20764_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_175_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22502_ _15154_/B _22387_/B _14273_/X vssd1 vssd1 vccd1 vccd1 _22502_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26270_ _26273_/CLK _26270_/D vssd1 vssd1 vccd1 vccd1 _26270_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_174_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23482_ _23457_/X _24959_/A _23256_/B _23481_/X vssd1 vssd1 vccd1 vccd1 _23482_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20694_ _20693_/Y _20192_/X _19236_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _20694_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25221_ _26306_/CLK hold373/X vssd1 vssd1 vccd1 vccd1 hold371/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22433_ _23245_/A vssd1 vssd1 vccd1 vccd1 _22433_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25152_ _26286_/CLK hold643/X vssd1 vssd1 vccd1 vccd1 hold641/A sky130_fd_sc_hd__dfxtp_1
X_22364_ _22362_/Y _22363_/Y _21897_/X vssd1 vssd1 vccd1 vccd1 _22364_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24103_ _24103_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24104_/A sky130_fd_sc_hd__and2_1
X_21315_ _21573_/A _21315_/B vssd1 vssd1 vccd1 vccd1 _21315_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_102_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25083_ _26167_/CLK _25083_/D vssd1 vssd1 vccd1 vccd1 _25083_/Q sky130_fd_sc_hd__dfxtp_1
X_22295_ _22295_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _22295_/X sky130_fd_sc_hd__and2_1
X_24034_ _24034_/A vssd1 vssd1 vccd1 vccd1 _26079_/D sky130_fd_sc_hd__clkbuf_1
Xhold350 hold350/A vssd1 vssd1 vccd1 vccd1 hold350/X sky130_fd_sc_hd__dlygate4sd3_1
X_21246_ _21675_/C vssd1 vssd1 vccd1 vccd1 _21678_/B sky130_fd_sc_hd__inv_2
Xhold361 hold361/A vssd1 vssd1 vccd1 vccd1 hold361/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold372 hold372/A vssd1 vssd1 vccd1 vccd1 hold372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 hold383/A vssd1 vssd1 vccd1 vccd1 hold383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 hold394/A vssd1 vssd1 vccd1 vccd1 hold394/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21177_ _21176_/Y _20192_/X _20986_/X _20957_/X vssd1 vssd1 vccd1 vccd1 _21177_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_102_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20128_ _20128_/A _20503_/B vssd1 vssd1 vccd1 vccd1 _20128_/Y sky130_fd_sc_hd__nand2_1
X_25985_ _25999_/CLK _25985_/D vssd1 vssd1 vccd1 vccd1 _25985_/Q sky130_fd_sc_hd__dfxtp_1
X_12950_ _12930_/X _12948_/X _12917_/X _12949_/X vssd1 vssd1 vccd1 vccd1 _12950_/X
+ sky130_fd_sc_hd__o211a_1
X_24936_ hold882/A hold912/A _24945_/S vssd1 vssd1 vccd1 vccd1 _24937_/B sky130_fd_sc_hd__mux2_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20059_ _20062_/A _20062_/B vssd1 vssd1 vccd1 vccd1 _20061_/A sky130_fd_sc_hd__nand2_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1050 _13462_/X vssd1 vssd1 vccd1 vccd1 _25129_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1061 _25106_/Q vssd1 vssd1 vccd1 vccd1 _18839_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1072 _13447_/X vssd1 vssd1 vccd1 vccd1 _25126_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 _25545_/Q vssd1 vssd1 vccd1 vccd1 _16743_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _26239_/Q _25608_/Q vssd1 vssd1 vccd1 vccd1 _14370_/A sky130_fd_sc_hd__xor2_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24867_ _24862_/X _24866_/X _24867_/S vssd1 vssd1 vccd1 vccd1 _24867_/X sky130_fd_sc_hd__mux2_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 _12782_/X vssd1 vssd1 vccd1 vccd1 _25008_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _14620_/A _14644_/B vssd1 vssd1 vccd1 vccd1 _14620_/Y sky130_fd_sc_hd__nand2_1
X_23818_ _23818_/A vssd1 vssd1 vccd1 vccd1 _26010_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24798_ _24798_/A vssd1 vssd1 vccd1 vccd1 _26327_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _14551_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14551_/Y sky130_fd_sc_hd__nand2_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23749_ _23749_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23750_/A sky130_fd_sc_hd__and2_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _13583_/A _13502_/B vssd1 vssd1 vccd1 vccd1 _13502_/Y sky130_fd_sc_hd__nand2_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17270_ _17268_/X _17241_/X _17269_/X vssd1 vssd1 vccd1 vccd1 _17271_/A sky130_fd_sc_hd__a21o_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _14482_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14482_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16221_ _16676_/A _16221_/B vssd1 vssd1 vccd1 vccd1 _16224_/A sky130_fd_sc_hd__or2_1
XFILLER_0_165_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13433_ _26335_/Q _25704_/Q vssd1 vssd1 vccd1 vccd1 _14672_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_181_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25419_ _25420_/CLK _25419_/D vssd1 vssd1 vccd1 vccd1 _25419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16152_ _16152_/A _16156_/B vssd1 vssd1 vccd1 vccd1 _16152_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_51_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13364_ _13315_/X _13362_/X _13300_/X _13363_/X vssd1 vssd1 vccd1 vccd1 _13364_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15103_ _15106_/B _15104_/A vssd1 vssd1 vccd1 vccd1 _15103_/X sky130_fd_sc_hd__or2_1
X_16083_ _16103_/A vssd1 vssd1 vccd1 vccd1 _16088_/B sky130_fd_sc_hd__inv_2
XFILLER_0_121_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13295_ _13295_/A vssd1 vssd1 vccd1 vccd1 _19546_/A sky130_fd_sc_hd__clkbuf_8
X_15034_ _15034_/A _15034_/B vssd1 vssd1 vccd1 vccd1 _15034_/Y sky130_fd_sc_hd__nor2_1
X_19911_ _20043_/A _18929_/A _20048_/C vssd1 vssd1 vccd1 vccd1 _19981_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_139_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19842_ _19841_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19843_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_177_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19773_ _19770_/Y _19773_/B _21789_/A vssd1 vssd1 vccd1 vccd1 _19773_/X sky130_fd_sc_hd__and3b_1
X_16985_ _21749_/A _16985_/B vssd1 vssd1 vccd1 vccd1 _17608_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_155_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18724_ _19774_/A vssd1 vssd1 vccd1 vccd1 _22436_/B sky130_fd_sc_hd__inv_2
X_15936_ _15936_/A _15940_/B vssd1 vssd1 vccd1 vccd1 _15936_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_189_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18655_ _18655_/A _20361_/A vssd1 vssd1 vccd1 vccd1 _18974_/A sky130_fd_sc_hd__xor2_4
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15867_ _15884_/C _15867_/B vssd1 vssd1 vccd1 vccd1 _15894_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17606_ _17604_/Y _17605_/Y _17568_/X vssd1 vssd1 vccd1 vccd1 _25638_/D sky130_fd_sc_hd__a21oi_1
X_14818_ _14818_/A vssd1 vssd1 vccd1 vccd1 _15006_/A sky130_fd_sc_hd__inv_2
XFILLER_0_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18586_ _25883_/Q _22266_/A vssd1 vssd1 vccd1 vccd1 _18594_/A sky130_fd_sc_hd__or2_2
X_15798_ _15798_/A vssd1 vssd1 vccd1 vccd1 _16974_/A sky130_fd_sc_hd__inv_2
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17537_ _17535_/X _17528_/X _17536_/X vssd1 vssd1 vccd1 vccd1 _17538_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_86_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14749_ _14749_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14749_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17468_ _17466_/Y _17467_/Y _17428_/X vssd1 vssd1 vccd1 vccd1 _17468_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19207_ _20467_/A _22131_/B _25594_/Q vssd1 vssd1 vccd1 vccd1 _20472_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16419_ _16420_/B _16420_/A vssd1 vssd1 vccd1 vccd1 _16421_/A sky130_fd_sc_hd__or2_1
XFILLER_0_183_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17399_ _21265_/B _25875_/Q _25811_/Q vssd1 vssd1 vccd1 vccd1 _17400_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_116_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19138_ _25649_/Q _19138_/B _19138_/C vssd1 vssd1 vccd1 vccd1 _20143_/A sky130_fd_sc_hd__or3_1
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19069_ _19067_/X _18879_/X _19068_/X vssd1 vssd1 vccd1 vccd1 _19070_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _26139_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21100_ _21097_/Y _21098_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21100_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_160_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22080_ _22081_/B _22081_/A vssd1 vssd1 vccd1 vccd1 _22082_/A sky130_fd_sc_hd__or2_1
XFILLER_0_160_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21031_ _21545_/C _21497_/C vssd1 vssd1 vccd1 vccd1 _21033_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22982_ _22982_/A _22982_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22984_/A sky130_fd_sc_hd__or3_1
X_25770_ _25770_/CLK _25770_/D vssd1 vssd1 vccd1 vccd1 _25770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21933_ _22653_/A _21933_/B vssd1 vssd1 vccd1 vccd1 _21933_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24721_ _24721_/A vssd1 vssd1 vccd1 vccd1 _26302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24652_ _24745_/A vssd1 vssd1 vccd1 vccd1 _24741_/B sky130_fd_sc_hd__clkbuf_16
X_21864_ _22653_/A _21864_/B vssd1 vssd1 vccd1 vccd1 _21864_/X sky130_fd_sc_hd__or2_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23603_ _23920_/S vssd1 vssd1 vccd1 vccd1 _23677_/S sky130_fd_sc_hd__clkbuf_16
X_20815_ _21235_/A _20815_/B vssd1 vssd1 vccd1 vccd1 _20815_/Y sky130_fd_sc_hd__nand2_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24583_ _24583_/A vssd1 vssd1 vccd1 vccd1 _26257_/D sky130_fd_sc_hd__clkbuf_1
X_21795_ _22680_/A vssd1 vssd1 vccd1 vccd1 _22653_/A sky130_fd_sc_hd__buf_8
XFILLER_0_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23534_ _24922_/S hold386/A _23533_/X vssd1 vssd1 vccd1 vccd1 _23534_/Y sky130_fd_sc_hd__o21ai_1
X_26322_ _26325_/CLK _26322_/D vssd1 vssd1 vccd1 vccd1 _26322_/Q sky130_fd_sc_hd__dfxtp_2
X_20746_ _20748_/B _20748_/C vssd1 vssd1 vccd1 vccd1 _20747_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26253_ _26267_/CLK _26253_/D vssd1 vssd1 vccd1 vccd1 _26253_/Q sky130_fd_sc_hd__dfxtp_4
X_23465_ _24956_/S hold341/A _23464_/X vssd1 vssd1 vccd1 vccd1 _23465_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20677_ _20677_/A _22544_/B _20677_/C vssd1 vssd1 vccd1 vccd1 _20681_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_135_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25204_ _25794_/CLK hold688/X vssd1 vssd1 vccd1 vccd1 hold686/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22416_ _22991_/B _22840_/B vssd1 vssd1 vccd1 vccd1 _22418_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26184_ _26184_/CLK _26184_/D vssd1 vssd1 vccd1 vccd1 _26184_/Q sky130_fd_sc_hd__dfxtp_1
X_23396_ hold203/A _23391_/A vssd1 vssd1 vccd1 vccd1 _23396_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_27_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25135_ _25135_/CLK hold532/X vssd1 vssd1 vccd1 vccd1 hold530/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22347_ _22347_/A _25886_/Q vssd1 vssd1 vccd1 vccd1 _22347_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_21_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13080_ _17653_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13080_/X sky130_fd_sc_hd__or2_1
X_25066_ _25712_/CLK _25066_/D vssd1 vssd1 vccd1 vccd1 _25066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22278_ _25791_/Q _22278_/B vssd1 vssd1 vccd1 vccd1 _22278_/Y sky130_fd_sc_hd__nor2_1
X_24017_ hold2253/X _26074_/Q _24047_/S vssd1 vssd1 vccd1 vccd1 _24017_/X sky130_fd_sc_hd__mux2_1
Xhold180 hold180/A vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__dlygate4sd3_1
X_21229_ _26312_/Q _21228_/X hold569/X vssd1 vssd1 vccd1 vccd1 _21232_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold191 hold191/A vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16770_ _16770_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16770_/Y sky130_fd_sc_hd__nand2_1
X_25968_ _26041_/CLK _25968_/D vssd1 vssd1 vccd1 vccd1 _25968_/Q sky130_fd_sc_hd__dfxtp_1
X_13982_ _25792_/Q vssd1 vssd1 vccd1 vccd1 _17847_/B sky130_fd_sc_hd__inv_2
X_15721_ _16949_/B vssd1 vssd1 vccd1 vccd1 _23111_/B sky130_fd_sc_hd__inv_2
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24919_ _24867_/S _24912_/Y _24914_/Y _24918_/X vssd1 vssd1 vccd1 vccd1 _24919_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ _26120_/Q _12907_/X _12932_/X vssd1 vssd1 vccd1 vccd1 _12933_/X sky130_fd_sc_hd__a21o_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25899_ _26084_/CLK _25899_/D vssd1 vssd1 vccd1 vccd1 _25899_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ _19574_/A vssd1 vssd1 vccd1 vccd1 _22065_/B sky130_fd_sc_hd__inv_2
X_15652_ _15795_/A _16571_/B vssd1 vssd1 vccd1 vccd1 _15655_/A sky130_fd_sc_hd__nor2_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _17322_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12864_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14603_ _14645_/A hold44/X vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ _18576_/A _18718_/A vssd1 vssd1 vccd1 vccd1 _18372_/B sky130_fd_sc_hd__xnor2_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15583_ _22982_/B _15583_/B vssd1 vssd1 vccd1 vccd1 _22979_/B sky130_fd_sc_hd__xor2_1
X_12795_ hold721/X _12748_/X _12794_/X vssd1 vssd1 vccd1 vccd1 _12795_/X sky130_fd_sc_hd__a21o_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17322_ _17393_/A _17322_/B _19994_/B vssd1 vssd1 vccd1 vccd1 _17322_/X sky130_fd_sc_hd__and3_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14534_ _14585_/A hold104/X vssd1 vssd1 vccd1 vccd1 hold105/A sky130_fd_sc_hd__nand2_1
XFILLER_0_138_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17253_ _25704_/Q _17253_/B vssd1 vssd1 vccd1 vccd1 _17615_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14465_ _14465_/A hold479/X vssd1 vssd1 vccd1 vccd1 hold480/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16204_ hold912/X _16205_/A vssd1 vssd1 vccd1 vccd1 _16206_/A sky130_fd_sc_hd__or2_1
XFILLER_0_114_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13416_ _26204_/Q _13239_/X _13415_/X vssd1 vssd1 vccd1 vccd1 _13416_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_113_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17184_ _19788_/A _17184_/B vssd1 vssd1 vccd1 vccd1 _17577_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14396_ _14394_/Y hold354/X _14345_/X vssd1 vssd1 vccd1 vccd1 hold355/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_183_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16135_ _16135_/A _16157_/B vssd1 vssd1 vccd1 vccd1 _16135_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_180_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13347_ _13347_/A vssd1 vssd1 vccd1 vccd1 _19659_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16066_ hold548/X vssd1 vssd1 vccd1 vccd1 _16069_/B sky130_fd_sc_hd__inv_2
X_13278_ _26310_/Q _19504_/A vssd1 vssd1 vccd1 vccd1 _14596_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15017_ _15003_/A _15030_/A _15016_/Y vssd1 vssd1 vccd1 vccd1 _15019_/A sky130_fd_sc_hd__a21o_1
Xhold2509 _24793_/X vssd1 vssd1 vccd1 vccd1 _24794_/A sky130_fd_sc_hd__dlygate4sd3_1
X_19825_ _19823_/Y _19824_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19825_/Y sky130_fd_sc_hd__a21oi_1
Xhold1808 _25858_/Q vssd1 vssd1 vccd1 vccd1 _22363_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1819 _25627_/Q vssd1 vssd1 vccd1 vccd1 _17524_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19756_ _19755_/Y _19483_/A _19104_/X _19105_/X vssd1 vssd1 vccd1 vccd1 _19757_/B
+ sky130_fd_sc_hd__a211o_1
X_16968_ _16966_/X _16711_/A _16967_/Y _25899_/Q _14170_/A vssd1 vssd1 vccd1 vccd1
+ _16969_/A sky130_fd_sc_hd__a32o_1
X_18707_ _18707_/A _18707_/B vssd1 vssd1 vccd1 vccd1 _22407_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15919_ _15934_/B _15919_/B vssd1 vssd1 vccd1 vccd1 _15940_/A sky130_fd_sc_hd__nand2_1
X_19687_ _19687_/A _20273_/B vssd1 vssd1 vccd1 vccd1 _19687_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_155_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16899_ _16899_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16899_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_188_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18638_ _19026_/A _18638_/B _18976_/C vssd1 vssd1 vccd1 vccd1 _18638_/X sky130_fd_sc_hd__and3_1
XFILLER_0_91_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18569_ _18569_/A _21412_/B _18569_/C vssd1 vssd1 vccd1 vccd1 _20208_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_75_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20600_ _23053_/B vssd1 vssd1 vccd1 vccd1 _22493_/B sky130_fd_sc_hd__inv_2
XFILLER_0_47_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21580_ _21580_/A _21580_/B _21580_/C vssd1 vssd1 vccd1 vccd1 _21581_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_144_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20531_ _20531_/A _20531_/B _21222_/C vssd1 vssd1 vccd1 vccd1 _20535_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23250_ _23248_/X hold1916/X _12702_/A vssd1 vssd1 vccd1 vccd1 _23250_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20462_ _20462_/A _20462_/B vssd1 vssd1 vccd1 vccd1 _20463_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_172_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22201_ _22561_/A _22201_/B vssd1 vssd1 vccd1 vccd1 _22201_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_127_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23181_ _23197_/A _23181_/B vssd1 vssd1 vccd1 vccd1 _23181_/Y sky130_fd_sc_hd__nand2_1
X_20393_ _25848_/Q vssd1 vssd1 vccd1 vccd1 _22081_/B sky130_fd_sc_hd__inv_2
XFILLER_0_42_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22132_ _17898_/A _25786_/Q _22130_/Y _22131_/Y vssd1 vssd1 vccd1 vccd1 _22133_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22063_ _22063_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _22063_/X sky130_fd_sc_hd__and2_1
X_21014_ _26304_/Q hold371/X vssd1 vssd1 vccd1 vccd1 _21014_/Y sky130_fd_sc_hd__nand2_1
X_25822_ _25822_/CLK _25822_/D vssd1 vssd1 vccd1 vccd1 _25822_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_173_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22965_ _22965_/A _22965_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22967_/A sky130_fd_sc_hd__or3_1
X_25753_ _25756_/CLK _25753_/D vssd1 vssd1 vccd1 vccd1 _25753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24704_ hold2674/X hold2580/X _24740_/S vssd1 vssd1 vccd1 vccd1 _24705_/A sky130_fd_sc_hd__mux2_1
X_21916_ _19504_/A _21915_/A _21915_/Y vssd1 vssd1 vccd1 vccd1 _21918_/A sky130_fd_sc_hd__o21ai_2
X_22896_ _22896_/A _22896_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22898_/A sky130_fd_sc_hd__or3_1
X_25684_ _26317_/CLK _25684_/D vssd1 vssd1 vccd1 vccd1 _25684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21847_ _19473_/A _21846_/A _21846_/Y vssd1 vssd1 vccd1 vccd1 _21849_/A sky130_fd_sc_hd__o21ai_2
X_24635_ _24635_/A vssd1 vssd1 vccd1 vccd1 _26274_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12580_ _24745_/A vssd1 vssd1 vccd1 vccd1 _23377_/B sky130_fd_sc_hd__buf_12
XFILLER_0_66_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24566_ hold2639/X _26252_/Q _24587_/S vssd1 vssd1 vccd1 vccd1 _24566_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_154_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21778_ _21778_/A _22587_/B vssd1 vssd1 vccd1 vccd1 _21779_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26305_ _26305_/CLK _26305_/D vssd1 vssd1 vccd1 vccd1 _26305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23517_ _24944_/S hold212/A _23516_/X vssd1 vssd1 vccd1 vccd1 _23517_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20729_ _20729_/A _20729_/B vssd1 vssd1 vccd1 vccd1 _20730_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_136_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24497_ _24497_/A vssd1 vssd1 vccd1 vccd1 _26229_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14250_ _18915_/B _14262_/B vssd1 vssd1 vccd1 vccd1 _14250_/Y sky130_fd_sc_hd__nor2_1
X_26236_ _26236_/CLK _26236_/D vssd1 vssd1 vccd1 vccd1 _26236_/Q sky130_fd_sc_hd__dfxtp_2
X_23448_ hold215/A _24945_/S vssd1 vssd1 vccd1 vccd1 _23448_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13201_ _13201_/A vssd1 vssd1 vccd1 vccd1 _19331_/A sky130_fd_sc_hd__buf_4
XFILLER_0_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14181_ hold699/X _14180_/Y _14155_/X vssd1 vssd1 vccd1 vccd1 hold700/A sky130_fd_sc_hd__a21oi_1
X_23379_ hold476/X _23380_/A vssd1 vssd1 vccd1 vccd1 _23379_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_26167_ _26167_/CLK _26167_/D vssd1 vssd1 vccd1 vccd1 _26167_/Q sky130_fd_sc_hd__dfxtp_1
X_13132_ _26158_/Q _13065_/X _13131_/X vssd1 vssd1 vccd1 vccd1 _13132_/X sky130_fd_sc_hd__a21o_1
X_25118_ _26200_/CLK _25118_/D vssd1 vssd1 vccd1 vccd1 _25118_/Q sky130_fd_sc_hd__dfxtp_1
X_26098_ _26103_/CLK _26098_/D vssd1 vssd1 vccd1 vccd1 _26098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17940_ _18611_/A _17944_/B vssd1 vssd1 vccd1 vccd1 _17942_/A sky130_fd_sc_hd__nand2_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25049_ _26135_/CLK _25049_/D vssd1 vssd1 vccd1 vccd1 _25049_/Q sky130_fd_sc_hd__dfxtp_1
X_13063_ _17632_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13063_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17871_ _21821_/A _25584_/Q vssd1 vssd1 vccd1 vccd1 _17873_/B sky130_fd_sc_hd__nand2_1
X_19610_ _19723_/A _19610_/B vssd1 vssd1 vccd1 vccd1 _19610_/Y sky130_fd_sc_hd__nand2_1
X_16822_ _16935_/A _16827_/B vssd1 vssd1 vccd1 vccd1 _16824_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19541_ _19539_/Y _19540_/Y _19382_/X vssd1 vssd1 vccd1 vccd1 _19541_/Y sky130_fd_sc_hd__a21oi_1
X_16753_ _16754_/B _16754_/A vssd1 vssd1 vccd1 vccd1 _16753_/X sky130_fd_sc_hd__or2_1
X_13965_ _26292_/Q _13801_/X _13793_/X _13964_/Y vssd1 vssd1 vccd1 vccd1 _13966_/B
+ sky130_fd_sc_hd__a22o_1
X_15704_ _16940_/B vssd1 vssd1 vccd1 vccd1 _23095_/B sky130_fd_sc_hd__inv_2
X_12916_ _26117_/Q _12907_/X _12915_/X vssd1 vssd1 vccd1 vccd1 _12916_/X sky130_fd_sc_hd__a21o_1
X_19472_ _19469_/Y _19472_/B _19980_/B vssd1 vssd1 vccd1 vccd1 _19472_/X sky130_fd_sc_hd__and3b_1
X_16684_ _16685_/B _16685_/A vssd1 vssd1 vccd1 vccd1 _16686_/A sky130_fd_sc_hd__or2_1
X_13896_ _17976_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13896_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_88_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18423_ _18423_/A _18423_/B vssd1 vssd1 vccd1 vccd1 _22039_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15635_ _23031_/B _15635_/B vssd1 vssd1 vccd1 vccd1 _23028_/B sky130_fd_sc_hd__xor2_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _12726_/B _14348_/A _12752_/X _25601_/Q vssd1 vssd1 vccd1 vccd1 _12847_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _18352_/X _18269_/X _18353_/X vssd1 vssd1 vccd1 vccd1 _18355_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_56_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15566_ _22965_/B _15566_/B vssd1 vssd1 vccd1 vccd1 _22962_/B sky130_fd_sc_hd__xor2_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12778_ _26219_/Q _25588_/Q vssd1 vssd1 vccd1 vccd1 _14307_/A sky130_fd_sc_hd__xor2_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17305_ _20044_/B _25900_/Q _25836_/Q vssd1 vssd1 vccd1 vccd1 _17306_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_185_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14517_ _14515_/Y hold180/X _14466_/X vssd1 vssd1 vccd1 vccd1 hold181/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18285_ _18951_/A _19554_/B vssd1 vssd1 vccd1 vccd1 _18288_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15497_ _15502_/A vssd1 vssd1 vccd1 vccd1 _15500_/B sky130_fd_sc_hd__inv_2
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17236_ _20712_/B _25895_/Q _25831_/Q vssd1 vssd1 vccd1 vccd1 _17237_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14448_ _14446_/Y hold273/X _14406_/X vssd1 vssd1 vccd1 vccd1 hold274/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17167_ _20702_/B _25856_/Q _25792_/Q vssd1 vssd1 vccd1 vccd1 _17168_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold905 hold905/A vssd1 vssd1 vccd1 vccd1 hold905/X sky130_fd_sc_hd__dlygate4sd3_1
X_14379_ _14379_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14379_/Y sky130_fd_sc_hd__nand2_1
Xhold916 hold916/A vssd1 vssd1 vccd1 vccd1 hold916/X sky130_fd_sc_hd__buf_1
Xhold927 hold927/A vssd1 vssd1 vccd1 vccd1 hold927/X sky130_fd_sc_hd__buf_1
X_16118_ _16212_/A hold428/X vssd1 vssd1 vccd1 vccd1 hold429/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold938 hold938/A vssd1 vssd1 vccd1 vccd1 hold938/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 hold949/A vssd1 vssd1 vccd1 vccd1 hold949/X sky130_fd_sc_hd__dlygate4sd3_1
X_17098_ _25588_/Q vssd1 vssd1 vccd1 vccd1 _20248_/B sky130_fd_sc_hd__inv_2
X_16049_ _16049_/A _16049_/B vssd1 vssd1 vccd1 vccd1 _16050_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2306 _15074_/Y vssd1 vssd1 vccd1 vccd1 _25432_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2317 _12662_/X vssd1 vssd1 vccd1 vccd1 _12663_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2328 _26204_/Q vssd1 vssd1 vccd1 vccd1 hold2328/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2339 _14953_/Y vssd1 vssd1 vccd1 vccd1 _25418_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1605 _17326_/Y vssd1 vssd1 vccd1 vccd1 _25604_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1616 _25601_/Q vssd1 vssd1 vccd1 vccd1 _17286_/B sky130_fd_sc_hd__dlygate4sd3_1
X_19808_ _19806_/X _19807_/Y _19764_/X vssd1 vssd1 vccd1 vccd1 _19808_/Y sky130_fd_sc_hd__a21oi_1
Xhold1627 _23006_/Y vssd1 vssd1 vccd1 vccd1 _25889_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1638 _17621_/Y vssd1 vssd1 vccd1 vccd1 _25640_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1649 _25590_/Q vssd1 vssd1 vccd1 vccd1 _17138_/B sky130_fd_sc_hd__clkbuf_2
X_19739_ _19736_/Y _19738_/Y _19653_/X vssd1 vssd1 vccd1 vccd1 _19739_/Y sky130_fd_sc_hd__a21oi_1
X_22750_ _22750_/A _22750_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22752_/A sky130_fd_sc_hd__or3_1
XFILLER_0_56_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21701_ _21701_/A _21701_/B vssd1 vssd1 vccd1 vccd1 _21702_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_176_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22681_ _15285_/B _22680_/X _14273_/X vssd1 vssd1 vccd1 vccd1 _22681_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_1253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24420_ _24420_/A vssd1 vssd1 vccd1 vccd1 _26204_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21632_ _21632_/A _22892_/B vssd1 vssd1 vccd1 vccd1 _21637_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24351_ _24351_/A _24373_/B vssd1 vssd1 vccd1 vccd1 _24352_/A sky130_fd_sc_hd__and2_1
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21563_ _21563_/A _21612_/A vssd1 vssd1 vccd1 vccd1 _21564_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_173_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23302_ hold985/X vssd1 vssd1 vccd1 vccd1 _23303_/B sky130_fd_sc_hd__inv_2
XFILLER_0_117_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20514_ _20513_/B _20514_/B _20514_/C vssd1 vssd1 vccd1 vccd1 _20515_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_172_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24282_ _24835_/S vssd1 vssd1 vccd1 vccd1 _24356_/S sky130_fd_sc_hd__clkbuf_16
X_21494_ _21491_/Y _21492_/Y _21493_/X vssd1 vssd1 vccd1 vccd1 _21494_/Y sky130_fd_sc_hd__a21oi_1
X_23233_ _23240_/A _24958_/B vssd1 vssd1 vccd1 vccd1 _23238_/A sky130_fd_sc_hd__nand2_1
X_26021_ _26021_/CLK _26021_/D vssd1 vssd1 vccd1 vccd1 _26021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20445_ _20447_/B vssd1 vssd1 vccd1 vccd1 _20446_/B sky130_fd_sc_hd__inv_2
XFILLER_0_63_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23164_ _23155_/Y _23163_/Y _19199_/A vssd1 vssd1 vccd1 vccd1 _23164_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20376_ _21198_/B _21514_/A vssd1 vssd1 vccd1 vccd1 _20378_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22115_ _22653_/A _22115_/B vssd1 vssd1 vccd1 vccd1 _22115_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23095_ _23095_/A _23095_/B _23191_/C vssd1 vssd1 vccd1 vccd1 _23097_/A sky130_fd_sc_hd__or3_1
XFILLER_0_30_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22046_ _22046_/A _22046_/B vssd1 vssd1 vccd1 vccd1 _22758_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_138_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25805_ _25808_/CLK _25805_/D vssd1 vssd1 vccd1 vccd1 _25805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23997_ _23997_/A vssd1 vssd1 vccd1 vccd1 _26067_/D sky130_fd_sc_hd__clkbuf_1
X_25736_ _25802_/CLK _25736_/D vssd1 vssd1 vccd1 vccd1 _25736_/Q sky130_fd_sc_hd__dfxtp_1
X_13750_ _18591_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13750_/Y sky130_fd_sc_hd__nor2_1
X_22948_ _22948_/A _22948_/B _22999_/C vssd1 vssd1 vccd1 vccd1 _22950_/A sky130_fd_sc_hd__or3_1
XFILLER_0_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12701_ _12701_/A hold997/X _24991_/Q vssd1 vssd1 vccd1 vccd1 _12702_/B sky130_fd_sc_hd__and3_1
XFILLER_0_97_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25667_ _26164_/CLK _25667_/D vssd1 vssd1 vccd1 vccd1 _25667_/Q sky130_fd_sc_hd__dfxtp_1
X_13681_ _13760_/A hold614/X vssd1 vssd1 vccd1 vccd1 hold615/A sky130_fd_sc_hd__nand2_1
X_22879_ _23188_/A _22879_/B vssd1 vssd1 vccd1 vccd1 _22879_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15420_ _22832_/B _15420_/B vssd1 vssd1 vccd1 vccd1 _22828_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_155_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12632_ _12632_/A vssd1 vssd1 vccd1 vccd1 _12635_/B sky130_fd_sc_hd__inv_2
XFILLER_0_39_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24618_ hold2646/X hold2608/X _24664_/S vssd1 vssd1 vccd1 vccd1 _24619_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_149_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25598_ _26109_/CLK _25598_/D vssd1 vssd1 vccd1 vccd1 _25598_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_109_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15351_ _22766_/B _15351_/B vssd1 vssd1 vccd1 vccd1 _22763_/B sky130_fd_sc_hd__xor2_1
X_12563_ _23597_/C _12564_/A vssd1 vssd1 vccd1 vccd1 _12570_/A sky130_fd_sc_hd__or2_1
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24549_ _24549_/A vssd1 vssd1 vccd1 vccd1 _26246_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14302_ _14344_/A hold236/X vssd1 vssd1 vccd1 vccd1 hold237/A sky130_fd_sc_hd__nand2_1
XFILLER_0_109_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18070_ _18070_/A _18070_/B vssd1 vssd1 vccd1 vccd1 _18074_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15282_ _16776_/B vssd1 vssd1 vccd1 vccd1 _22683_/B sky130_fd_sc_hd__inv_2
X_12494_ _13220_/A vssd1 vssd1 vccd1 vccd1 _12726_/B sky130_fd_sc_hd__buf_12
XFILLER_0_25_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17021_ _25590_/Q vssd1 vssd1 vccd1 vccd1 _20310_/B sky130_fd_sc_hd__inv_2
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26219_ _26219_/CLK _26219_/D vssd1 vssd1 vccd1 vccd1 _26219_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14233_ _26335_/Q _13518_/B _14170_/X _14232_/Y vssd1 vssd1 vccd1 vccd1 _14234_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14164_ _25821_/Q vssd1 vssd1 vccd1 vccd1 _18633_/B sky130_fd_sc_hd__inv_2
XFILLER_0_33_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13115_ _26283_/Q _25652_/Q vssd1 vssd1 vccd1 vccd1 _14509_/A sky130_fd_sc_hd__xor2_1
X_14095_ _25810_/Q vssd1 vssd1 vccd1 vccd1 _18409_/B sky130_fd_sc_hd__inv_2
X_18972_ _18986_/A _19701_/A vssd1 vssd1 vccd1 vccd1 _18972_/Y sky130_fd_sc_hd__nand2_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ _17923_/A _17923_/B _20144_/A vssd1 vssd1 vccd1 vccd1 _17933_/A sky130_fd_sc_hd__and3_1
X_13046_ _26142_/Q _12907_/X _13045_/X vssd1 vssd1 vccd1 vccd1 _13046_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_147_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17854_ _18611_/A _17858_/B vssd1 vssd1 vccd1 vccd1 _17856_/A sky130_fd_sc_hd__nand2_1
X_16805_ _16805_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16805_/Y sky130_fd_sc_hd__nand2_1
X_17785_ _18119_/B vssd1 vssd1 vccd1 vccd1 _18153_/B sky130_fd_sc_hd__inv_2
XFILLER_0_89_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14997_ _14997_/A _14997_/B vssd1 vssd1 vccd1 vccd1 _15015_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_163_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19524_ _19522_/X _19523_/Y _19494_/X vssd1 vssd1 vccd1 vccd1 _19524_/Y sky130_fd_sc_hd__a21oi_1
X_16736_ _16858_/A _16736_/B vssd1 vssd1 vccd1 vccd1 _16736_/Y sky130_fd_sc_hd__nand2_1
X_13948_ _14061_/A _13948_/B vssd1 vssd1 vccd1 vccd1 _13948_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19455_ _26237_/Q hold491/X vssd1 vssd1 vccd1 vccd1 _19455_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16667_ _16667_/A _16667_/B vssd1 vssd1 vccd1 vccd1 _16668_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13879_ hold603/X _13878_/Y _13798_/X vssd1 vssd1 vccd1 vccd1 hold604/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18406_ _18792_/A _25746_/Q vssd1 vssd1 vccd1 vccd1 _18409_/A sky130_fd_sc_hd__nand2_1
X_15618_ _15618_/A _15810_/B vssd1 vssd1 vccd1 vccd1 _15619_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_29_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19386_ _19385_/Y _19272_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19387_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16598_ _16598_/A _16598_/B vssd1 vssd1 vccd1 vccd1 _16599_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_174_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18337_ _18335_/Y _18336_/Y _18112_/X vssd1 vssd1 vccd1 vccd1 _25661_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15549_ _15549_/A vssd1 vssd1 vccd1 vccd1 _15577_/B sky130_fd_sc_hd__inv_2
XFILLER_0_155_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18268_ _19052_/A _18268_/B vssd1 vssd1 vccd1 vccd1 _18268_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_114_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17219_ _25604_/Q vssd1 vssd1 vccd1 vccd1 _20856_/B sky130_fd_sc_hd__inv_2
XFILLER_0_53_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18199_ _18446_/A _25736_/Q _18952_/C vssd1 vssd1 vccd1 vccd1 _18200_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_102_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold702 hold702/A vssd1 vssd1 vccd1 vccd1 hold702/X sky130_fd_sc_hd__dlygate4sd3_1
X_20230_ _21042_/A _20230_/B _20229_/X vssd1 vssd1 vccd1 vccd1 _20231_/B sky130_fd_sc_hd__or3b_1
Xhold713 hold713/A vssd1 vssd1 vccd1 vccd1 hold713/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 hold724/A vssd1 vssd1 vccd1 vccd1 hold724/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold735 hold735/A vssd1 vssd1 vccd1 vccd1 hold735/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 hold746/A vssd1 vssd1 vccd1 vccd1 hold746/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 hold757/A vssd1 vssd1 vccd1 vccd1 hold757/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold768 hold768/A vssd1 vssd1 vccd1 vccd1 hold768/X sky130_fd_sc_hd__dlygate4sd3_1
X_20161_ _20159_/Y _20160_/Y _19918_/X vssd1 vssd1 vccd1 vccd1 _20161_/Y sky130_fd_sc_hd__a21oi_1
Xhold779 hold779/A vssd1 vssd1 vccd1 vccd1 hold779/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2103 _26303_/Q vssd1 vssd1 vccd1 vccd1 hold2103/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2114 _23325_/X vssd1 vssd1 vccd1 vccd1 _23326_/A sky130_fd_sc_hd__dlygate4sd3_1
X_20092_ _20092_/A _23197_/B _20092_/C vssd1 vssd1 vccd1 vccd1 _20095_/C sky130_fd_sc_hd__nand3_1
Xhold2125 _24105_/X vssd1 vssd1 vccd1 vccd1 _24106_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2136 _26033_/Q vssd1 vssd1 vccd1 vccd1 hold2136/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_205_clk _26093_/CLK vssd1 vssd1 vccd1 vccd1 _26096_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2147 _25434_/Q vssd1 vssd1 vccd1 vccd1 _15083_/B sky130_fd_sc_hd__dlygate4sd3_1
X_23920_ _26043_/Q hold1976/X _23920_/S vssd1 vssd1 vccd1 vccd1 _23920_/X sky130_fd_sc_hd__mux2_1
Xhold1402 _13308_/X vssd1 vssd1 vccd1 vccd1 _25103_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1413 _25893_/Q vssd1 vssd1 vccd1 vccd1 _23069_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2158 _24178_/X vssd1 vssd1 vccd1 vccd1 _24179_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1424 _13140_/X vssd1 vssd1 vccd1 vccd1 _25076_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2169 _23347_/Y vssd1 vssd1 vccd1 vccd1 _23348_/C sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1435 _25110_/Q vssd1 vssd1 vccd1 vccd1 _18920_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1446 _19965_/Y vssd1 vssd1 vccd1 vccd1 _25770_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23851_ _23851_/A _23905_/B vssd1 vssd1 vccd1 vccd1 _23852_/A sky130_fd_sc_hd__and2_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1457 _25778_/Q vssd1 vssd1 vccd1 vccd1 _20197_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1468 _14805_/Y vssd1 vssd1 vccd1 vccd1 _25400_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1479 _25052_/Q vssd1 vssd1 vccd1 vccd1 _17557_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22802_ _16820_/B _22421_/X _22796_/X _22797_/Y _22801_/X vssd1 vssd1 vccd1 vccd1
+ _22803_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_170_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23782_ _14851_/B _14859_/B _23831_/S vssd1 vssd1 vccd1 vccd1 _23783_/A sky130_fd_sc_hd__mux2_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20994_ _20994_/A _20994_/B vssd1 vssd1 vccd1 vccd1 _20998_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25521_ _25534_/CLK hold936/X vssd1 vssd1 vccd1 vccd1 hold935/A sky130_fd_sc_hd__dfxtp_1
X_22733_ _26056_/Q vssd1 vssd1 vccd1 vccd1 _22734_/A sky130_fd_sc_hd__inv_2
XFILLER_0_48_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_25452_ _25539_/CLK _25452_/D vssd1 vssd1 vccd1 vccd1 _25452_/Q sky130_fd_sc_hd__dfxtp_1
X_22664_ _22664_/A _25899_/Q vssd1 vssd1 vccd1 vccd1 _22664_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_177_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21615_ _22704_/A vssd1 vssd1 vccd1 vccd1 _22892_/B sky130_fd_sc_hd__buf_6
X_24403_ hold2310/X _26199_/Q _24433_/S vssd1 vssd1 vccd1 vccd1 _24403_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25383_ _26334_/CLK hold349/X vssd1 vssd1 vccd1 vccd1 hold347/A sky130_fd_sc_hd__dfxtp_1
X_22595_ _22595_/A _22595_/B vssd1 vssd1 vccd1 vccd1 _22596_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24334_ _24334_/A vssd1 vssd1 vccd1 vccd1 _26176_/D sky130_fd_sc_hd__clkbuf_1
X_21546_ _21546_/A _21595_/A vssd1 vssd1 vccd1 vccd1 _21548_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_106_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24265_ _24265_/A _24280_/B vssd1 vssd1 vccd1 vccd1 _24266_/A sky130_fd_sc_hd__and2_1
XFILLER_0_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21477_ _21475_/Y _21476_/Y _21099_/X vssd1 vssd1 vccd1 vccd1 _21477_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_161_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23216_ _24863_/S vssd1 vssd1 vccd1 vccd1 _24945_/S sky130_fd_sc_hd__buf_12
X_26004_ _26004_/CLK _26004_/D vssd1 vssd1 vccd1 vccd1 _26004_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_31_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20428_ _20428_/A _22106_/A vssd1 vssd1 vccd1 vccd1 _20429_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24196_ _24196_/A vssd1 vssd1 vccd1 vccd1 _26131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23147_ _23147_/A _23195_/B vssd1 vssd1 vccd1 vccd1 _23147_/Y sky130_fd_sc_hd__nand2_1
X_20359_ _20359_/A _20359_/B vssd1 vssd1 vccd1 vccd1 _21195_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_140_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_23078_ _26077_/Q vssd1 vssd1 vccd1 vccd1 _23079_/A sky130_fd_sc_hd__inv_2
XFILLER_0_101_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14920_ _23245_/A _14920_/B _14925_/A vssd1 vssd1 vccd1 vccd1 _14921_/A sky130_fd_sc_hd__or3b_1
X_22029_ _22030_/A _22030_/B _23026_/A vssd1 vssd1 vccd1 vccd1 _22029_/X sky130_fd_sc_hd__a21o_1
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2670 _15325_/Y vssd1 vssd1 vccd1 vccd1 _25447_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2681 _15820_/Y vssd1 vssd1 vccd1 vccd1 hold2681/X sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ _14893_/A _14851_/B vssd1 vssd1 vccd1 vccd1 _22263_/A sky130_fd_sc_hd__nand2_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2692 _24796_/X vssd1 vssd1 vccd1 vccd1 _24797_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13802_ _25763_/Q vssd1 vssd1 vccd1 vccd1 _18753_/B sky130_fd_sc_hd__inv_2
Xhold1980 _26002_/Q vssd1 vssd1 vccd1 vccd1 _14884_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17570_ _17570_/A _17622_/A vssd1 vssd1 vccd1 vccd1 _17571_/B sky130_fd_sc_hd__xnor2_1
Xhold1991 _25946_/Q vssd1 vssd1 vccd1 vccd1 hold1991/X sky130_fd_sc_hd__dlygate4sd3_1
X_14782_ _14782_/A vssd1 vssd1 vccd1 vccd1 _14972_/A sky130_fd_sc_hd__inv_2
XFILLER_0_98_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16521_ _16522_/B _16522_/A vssd1 vssd1 vccd1 vccd1 _16537_/B sky130_fd_sc_hd__or2_1
X_25719_ _26239_/CLK hold893/X vssd1 vssd1 vccd1 vccd1 hold891/A sky130_fd_sc_hd__dfxtp_1
X_13733_ _26255_/Q _13612_/X _13605_/X _13732_/Y vssd1 vssd1 vccd1 vccd1 _13734_/B
+ sky130_fd_sc_hd__a22o_1
X_19240_ _19234_/X _18879_/X _19239_/X vssd1 vssd1 vccd1 vccd1 _19241_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16452_ _16452_/A _16452_/B vssd1 vssd1 vccd1 vccd1 _16461_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_151_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13664_ _18307_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13664_/Y sky130_fd_sc_hd__nor2_1
X_15403_ _16824_/A _15403_/B vssd1 vssd1 vccd1 vccd1 _15403_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ _12615_/A vssd1 vssd1 vccd1 vccd1 _24976_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19171_ _19169_/Y hold816/X _19086_/X vssd1 vssd1 vccd1 vccd1 hold817/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16383_ _16370_/Y _16374_/B _16372_/B vssd1 vssd1 vccd1 vccd1 _16383_/Y sky130_fd_sc_hd__o21ai_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13595_ _26233_/Q _13426_/X _13468_/X _13594_/Y vssd1 vssd1 vccd1 vccd1 _13596_/B
+ sky130_fd_sc_hd__a22o_1
X_18122_ _18122_/A _18122_/B _18122_/C vssd1 vssd1 vccd1 vccd1 _18125_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_81_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15334_ _15334_/A _15812_/B vssd1 vssd1 vccd1 vccd1 _15335_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_53_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12546_ _20957_/A vssd1 vssd1 vccd1 vccd1 _12546_/X sky130_fd_sc_hd__buf_12
XFILLER_0_26_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18053_ _18053_/A _18053_/B _18053_/C vssd1 vssd1 vccd1 vccd1 _21837_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_81_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15265_ _15265_/A vssd1 vssd1 vccd1 vccd1 _15307_/B sky130_fd_sc_hd__inv_2
XANTENNA_4 _22199_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17004_ _17794_/A vssd1 vssd1 vccd1 vccd1 _22786_/A sky130_fd_sc_hd__inv_16
X_14216_ _14264_/A _14216_/B vssd1 vssd1 vccd1 vccd1 _14216_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15196_ hold927/X vssd1 vssd1 vccd1 vccd1 _15198_/A sky130_fd_sc_hd__inv_2
XFILLER_0_111_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14147_ _26321_/Q _13988_/X _13981_/X _14146_/Y vssd1 vssd1 vccd1 vccd1 _14148_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14078_ _18348_/B _14114_/B vssd1 vssd1 vccd1 vccd1 _14078_/Y sky130_fd_sc_hd__nor2_1
X_18955_ _18955_/A _18955_/B _18955_/C vssd1 vssd1 vccd1 vccd1 _18956_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_184_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17906_ _17906_/A _25793_/Q _17906_/C vssd1 vssd1 vccd1 vccd1 _20747_/B sky130_fd_sc_hd__nand3_1
X_13029_ _26267_/Q _25636_/Q vssd1 vssd1 vccd1 vccd1 _14458_/A sky130_fd_sc_hd__xor2_2
X_18886_ _25706_/Q vssd1 vssd1 vccd1 vccd1 _22640_/B sky130_fd_sc_hd__inv_2
X_17837_ _19289_/A vssd1 vssd1 vccd1 vccd1 _22308_/B sky130_fd_sc_hd__inv_2
XFILLER_0_179_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17768_ _17768_/A _17781_/C vssd1 vssd1 vccd1 vccd1 _17771_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_178_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16719_ _16719_/A _16719_/B vssd1 vssd1 vccd1 vccd1 _16719_/Y sky130_fd_sc_hd__nand2_1
X_19507_ _19523_/B _19593_/B vssd1 vssd1 vccd1 vccd1 _19509_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17699_ _17699_/A _17699_/B _17764_/B vssd1 vssd1 vccd1 vccd1 _17705_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_77_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19438_ _19452_/A _19438_/B vssd1 vssd1 vccd1 vccd1 _19438_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_146_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19369_ _26231_/Q _12537_/B hold464/X vssd1 vssd1 vccd1 vccd1 _19369_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21400_ _21400_/A _21400_/B _21400_/C vssd1 vssd1 vccd1 vccd1 _21404_/A sky130_fd_sc_hd__nand3_1
X_22380_ _22381_/A _22381_/C _23087_/A vssd1 vssd1 vccd1 vccd1 _22380_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_128_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21331_ _21573_/A _21331_/B vssd1 vssd1 vccd1 vccd1 _21331_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_115_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24050_ _24050_/A _24050_/B vssd1 vssd1 vccd1 vccd1 _24743_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold510 hold510/A vssd1 vssd1 vccd1 vccd1 hold510/X sky130_fd_sc_hd__dlygate4sd3_1
X_21262_ _21573_/A _21262_/B vssd1 vssd1 vccd1 vccd1 _21262_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold521 hold521/A vssd1 vssd1 vccd1 vccd1 hold521/X sky130_fd_sc_hd__dlygate4sd3_1
X_23001_ _23001_/A _23001_/B _23001_/C vssd1 vssd1 vccd1 vccd1 _23001_/X sky130_fd_sc_hd__and3_1
Xhold532 hold532/A vssd1 vssd1 vccd1 vccd1 hold532/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20213_ _20213_/A _25843_/Q vssd1 vssd1 vccd1 vccd1 _20217_/B sky130_fd_sc_hd__nand2_1
Xhold543 hold543/A vssd1 vssd1 vccd1 vccd1 hold543/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold554 hold554/A vssd1 vssd1 vccd1 vccd1 hold554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 hold565/A vssd1 vssd1 vccd1 vccd1 hold565/X sky130_fd_sc_hd__dlygate4sd3_1
X_21193_ _21646_/B _21594_/C vssd1 vssd1 vccd1 vccd1 _21195_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold576 hold576/A vssd1 vssd1 vccd1 vccd1 hold576/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold587 hold587/A vssd1 vssd1 vccd1 vccd1 hold587/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 hold598/A vssd1 vssd1 vccd1 vccd1 hold598/X sky130_fd_sc_hd__dlygate4sd3_1
X_20144_ _20144_/A _20144_/B vssd1 vssd1 vccd1 vccd1 _20145_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_99_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24952_ _24952_/A _24956_/S vssd1 vssd1 vccd1 vccd1 _24952_/Y sky130_fd_sc_hd__nand2_1
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20075_ _20075_/A _20978_/C _20075_/C vssd1 vssd1 vccd1 vccd1 _20076_/B sky130_fd_sc_hd__nand3_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 _13169_/X vssd1 vssd1 vccd1 vccd1 _25081_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 _25751_/Q vssd1 vssd1 vccd1 vccd1 _19709_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1232 _25573_/Q vssd1 vssd1 vccd1 vccd1 _16933_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_23903_ _23903_/A vssd1 vssd1 vccd1 vccd1 _26038_/D sky130_fd_sc_hd__clkbuf_1
Xhold1243 _16957_/Y vssd1 vssd1 vccd1 vccd1 _25576_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24883_ _24946_/A _24883_/B vssd1 vssd1 vccd1 vccd1 _24883_/X sky130_fd_sc_hd__or2_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1254 _25548_/Q vssd1 vssd1 vccd1 vccd1 _16764_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1265 _14778_/Y vssd1 vssd1 vccd1 vccd1 _25397_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1276 _25544_/Q vssd1 vssd1 vccd1 vccd1 _16736_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1287 _14849_/Y vssd1 vssd1 vccd1 vccd1 _25405_/D sky130_fd_sc_hd__dlygate4sd3_1
X_23834_ _23920_/S vssd1 vssd1 vccd1 vccd1 _23907_/S sky130_fd_sc_hd__clkbuf_16
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1298 _25045_/Q vssd1 vssd1 vccd1 vccd1 _17507_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23765_ _23765_/A _23813_/B vssd1 vssd1 vccd1 vccd1 _23766_/A sky130_fd_sc_hd__and2_1
X_20977_ _21516_/B _21467_/B vssd1 vssd1 vccd1 vccd1 _20978_/B sky130_fd_sc_hd__nand2_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25504_ _25510_/CLK _25504_/D vssd1 vssd1 vccd1 vccd1 hold957/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22716_ _22714_/X _22715_/Y _22433_/X vssd1 vssd1 vccd1 vccd1 _22716_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23696_ hold2111/X hold2072/X _23754_/S vssd1 vssd1 vccd1 vccd1 _23697_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_83_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25435_ _26047_/CLK _25435_/D vssd1 vssd1 vccd1 vccd1 _25435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22647_ _23136_/B vssd1 vssd1 vccd1 vccd1 _23135_/B sky130_fd_sc_hd__inv_2
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13380_ _26198_/Q _13239_/X _13379_/X vssd1 vssd1 vccd1 vccd1 _13380_/X sky130_fd_sc_hd__a21o_1
X_22578_ _15208_/B _22387_/B _14273_/X vssd1 vssd1 vccd1 vccd1 _22578_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25366_ _26193_/CLK hold235/X vssd1 vssd1 vccd1 vccd1 hold233/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_24317_ hold2362/X hold2037/X _24356_/S vssd1 vssd1 vccd1 vccd1 _24318_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21529_ _21529_/A _21529_/B _21529_/C vssd1 vssd1 vccd1 vccd1 _21533_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25297_ _26249_/CLK hold202/X vssd1 vssd1 vccd1 vccd1 hold200/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15050_ _15050_/A _15050_/B vssd1 vssd1 vccd1 vccd1 _15067_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_160_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24248_ _24248_/A vssd1 vssd1 vccd1 vccd1 _26148_/D sky130_fd_sc_hd__clkbuf_1
X_14001_ _25795_/Q vssd1 vssd1 vccd1 vccd1 _18003_/B sky130_fd_sc_hd__inv_2
X_24179_ _24179_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24180_/A sky130_fd_sc_hd__and2_1
XFILLER_0_102_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18740_ _18738_/X _18269_/X _18739_/X vssd1 vssd1 vccd1 vccd1 _18741_/A sky130_fd_sc_hd__a21o_1
X_15952_ _15961_/B _15952_/B vssd1 vssd1 vccd1 vccd1 _16000_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_76_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14903_ _14903_/A _14903_/B vssd1 vssd1 vccd1 vccd1 _14904_/A sky130_fd_sc_hd__nand2_1
X_18671_ _18671_/A _25823_/Q _18671_/C vssd1 vssd1 vccd1 vccd1 _20409_/B sky130_fd_sc_hd__nand3_2
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15883_ _15884_/B _15884_/C _15894_/B vssd1 vssd1 vccd1 vccd1 _15883_/X sky130_fd_sc_hd__a21bo_1
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17622_ _17622_/A _17622_/B vssd1 vssd1 vccd1 vccd1 _17623_/B sky130_fd_sc_hd__xnor2_1
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14834_ hold955/X _22204_/A vssd1 vssd1 vccd1 vccd1 _22203_/B sky130_fd_sc_hd__xnor2_1
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17553_ _17605_/A _17553_/B vssd1 vssd1 vccd1 vccd1 _17553_/Y sky130_fd_sc_hd__nand2_1
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _25845_/Q _12527_/A _14955_/A _14696_/Y vssd1 vssd1 vccd1 vccd1 _14765_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16504_ _16513_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16504_/Y sky130_fd_sc_hd__nand2_1
X_13716_ _13823_/A _13716_/B vssd1 vssd1 vccd1 vccd1 _13716_/Y sky130_fd_sc_hd__nand2_1
X_17484_ _17534_/A _17651_/B vssd1 vssd1 vccd1 vccd1 _17485_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14696_ _22893_/A vssd1 vssd1 vccd1 vccd1 _14696_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19223_ _19221_/Y _21228_/A _19104_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _19225_/A
+ sky130_fd_sc_hd__a211o_1
X_16435_ _16676_/A _16435_/B vssd1 vssd1 vccd1 vccd1 _16437_/A sky130_fd_sc_hd__or2_1
XFILLER_0_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13647_ _13703_/A _13647_/B vssd1 vssd1 vccd1 vccd1 _13647_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_156_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19154_ _19153_/Y _19130_/X _19131_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _19157_/A
+ sky130_fd_sc_hd__a211o_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _16366_/A _16697_/B _16374_/A vssd1 vssd1 vccd1 vccd1 _16366_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_171_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13578_ hold787/X _13577_/Y _13559_/X vssd1 vssd1 vccd1 vccd1 hold788/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18105_ _19080_/A _18494_/A vssd1 vssd1 vccd1 vccd1 _18106_/B sky130_fd_sc_hd__xnor2_2
X_15317_ _22734_/B _15317_/B vssd1 vssd1 vccd1 vccd1 _22731_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12529_ _17008_/B vssd1 vssd1 vccd1 vccd1 _12529_/Y sky130_fd_sc_hd__inv_2
X_19085_ _19186_/A _19085_/B vssd1 vssd1 vccd1 vccd1 _19085_/Y sky130_fd_sc_hd__nand2_1
X_16297_ _16297_/A _16297_/B vssd1 vssd1 vccd1 vccd1 _16299_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18036_ _20592_/B _22221_/A vssd1 vssd1 vccd1 vccd1 _20585_/A sky130_fd_sc_hd__nand2_4
X_15248_ _15248_/A _15248_/B vssd1 vssd1 vccd1 vccd1 _15266_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_23_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15179_ _15184_/A vssd1 vssd1 vccd1 vccd1 _15182_/B sky130_fd_sc_hd__inv_2
X_19987_ _20660_/A _19987_/B vssd1 vssd1 vccd1 vccd1 _19987_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18938_ _18938_/A _20043_/A vssd1 vssd1 vccd1 vccd1 _19073_/B sky130_fd_sc_hd__xor2_4
.ends

