magic
tech sky130A
timestamp 1730450942
<< nwell >>
rect -130 -40 180 340
<< pwell >>
rect -130 -350 180 -70
<< nmos >>
rect 0 -310 120 -110
<< pmos >>
rect 0 0 120 300
<< ndiff >>
rect -40 -120 0 -110
rect -40 -140 -30 -120
rect -10 -140 0 -120
rect -40 -160 0 -140
rect -40 -180 -30 -160
rect -10 -180 0 -160
rect -40 -200 0 -180
rect -40 -220 -30 -200
rect -10 -220 0 -200
rect -40 -240 0 -220
rect -40 -260 -30 -240
rect -10 -260 0 -240
rect -40 -280 0 -260
rect -40 -300 -30 -280
rect -10 -300 0 -280
rect -40 -310 0 -300
rect 120 -120 160 -110
rect 120 -140 130 -120
rect 150 -140 160 -120
rect 120 -160 160 -140
rect 120 -180 130 -160
rect 150 -180 160 -160
rect 120 -200 160 -180
rect 120 -220 130 -200
rect 150 -220 160 -200
rect 120 -240 160 -220
rect 120 -260 130 -240
rect 150 -260 160 -240
rect 120 -280 160 -260
rect 120 -300 130 -280
rect 150 -300 160 -280
rect 120 -310 160 -300
<< pdiff >>
rect -40 290 0 300
rect -40 270 -30 290
rect -10 270 0 290
rect -40 250 0 270
rect -40 230 -30 250
rect -10 230 0 250
rect -40 210 0 230
rect -40 190 -30 210
rect -10 190 0 210
rect -40 170 0 190
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 90 0 110
rect -40 70 -30 90
rect -10 70 0 90
rect -40 50 0 70
rect -40 30 -30 50
rect -10 30 0 50
rect -40 0 0 30
rect 120 290 160 300
rect 120 270 130 290
rect 150 270 160 290
rect 120 250 160 270
rect 120 230 130 250
rect 150 230 160 250
rect 120 210 160 230
rect 120 190 130 210
rect 150 190 160 210
rect 120 170 160 190
rect 120 150 130 170
rect 150 150 160 170
rect 120 130 160 150
rect 120 110 130 130
rect 150 110 160 130
rect 120 90 160 110
rect 120 70 130 90
rect 150 70 160 90
rect 120 50 160 70
rect 120 30 130 50
rect 150 30 160 50
rect 120 0 160 30
<< ndiffc >>
rect -30 -140 -10 -120
rect -30 -180 -10 -160
rect -30 -220 -10 -200
rect -30 -260 -10 -240
rect -30 -300 -10 -280
rect 130 -140 150 -120
rect 130 -180 150 -160
rect 130 -220 150 -200
rect 130 -260 150 -240
rect 130 -300 150 -280
<< pdiffc >>
rect -30 270 -10 290
rect -30 230 -10 250
rect -30 190 -10 210
rect -30 150 -10 170
rect -30 110 -10 130
rect -30 70 -10 90
rect -30 30 -10 50
rect 130 270 150 290
rect 130 230 150 250
rect 130 190 150 210
rect 130 150 150 170
rect 130 110 150 130
rect 130 70 150 90
rect 130 30 150 50
<< psubdiff >>
rect -110 -280 -70 -265
rect -110 -300 -100 -280
rect -80 -300 -70 -280
rect -110 -315 -70 -300
<< nsubdiff >>
rect -110 280 -70 295
rect -110 260 -100 280
rect -80 260 -70 280
rect -110 245 -70 260
<< psubdiffcont >>
rect -100 -300 -80 -280
<< nsubdiffcont >>
rect -100 260 -80 280
<< poly >>
rect 0 300 120 340
rect 0 -110 120 0
rect 0 -350 120 -310
<< locali >>
rect -40 295 0 300
rect -110 290 0 295
rect -110 280 -30 290
rect -110 260 -100 280
rect -80 270 -30 280
rect -10 270 0 290
rect -80 260 0 270
rect -110 250 0 260
rect -110 245 -30 250
rect -40 230 -30 245
rect -10 230 0 250
rect -40 210 0 230
rect -40 190 -30 210
rect -10 190 0 210
rect -40 170 0 190
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 90 0 110
rect -40 70 -30 90
rect -10 70 0 90
rect -40 50 0 70
rect -40 30 -30 50
rect -10 30 0 50
rect -40 0 0 30
rect 120 290 160 300
rect 120 270 130 290
rect 150 270 160 290
rect 120 250 160 270
rect 120 230 130 250
rect 150 230 160 250
rect 120 210 160 230
rect 120 190 130 210
rect 150 190 160 210
rect 120 170 160 190
rect 120 150 130 170
rect 150 150 160 170
rect 120 130 160 150
rect 120 110 130 130
rect 150 110 160 130
rect 120 90 160 110
rect 120 70 130 90
rect 150 70 160 90
rect 120 50 160 70
rect 120 30 130 50
rect 150 30 160 50
rect -40 -120 0 -110
rect -40 -140 -30 -120
rect -10 -140 0 -120
rect -40 -160 0 -140
rect -40 -180 -30 -160
rect -10 -180 0 -160
rect -40 -200 0 -180
rect -40 -220 -30 -200
rect -10 -220 0 -200
rect -40 -240 0 -220
rect -40 -260 -30 -240
rect -10 -260 0 -240
rect -40 -265 0 -260
rect -110 -280 0 -265
rect -110 -300 -100 -280
rect -80 -300 -30 -280
rect -10 -300 0 -280
rect -110 -310 0 -300
rect 120 -120 160 30
rect 120 -140 130 -120
rect 150 -140 160 -120
rect 120 -160 160 -140
rect 120 -180 130 -160
rect 150 -180 160 -160
rect 120 -200 160 -180
rect 120 -220 130 -200
rect 150 -220 160 -200
rect 120 -240 160 -220
rect 120 -260 130 -240
rect 150 -260 160 -240
rect 120 -280 160 -260
rect 120 -300 130 -280
rect 150 -300 160 -280
rect 120 -310 160 -300
rect -110 -315 -70 -310
<< viali >>
rect -100 260 -80 280
rect -100 -300 -80 -280
<< metal1 >>
rect -110 280 -70 295
rect -110 260 -100 280
rect -80 260 -70 280
rect -110 245 -70 260
rect -110 -280 -70 -265
rect -110 -300 -100 -280
rect -80 -300 -70 -280
rect -110 -315 -70 -300
<< labels >>
rlabel poly 0 -55 0 -55 7 A
port 1 w
rlabel locali -20 300 -20 300 1 VDDA
port 3 n
rlabel locali -20 -310 -20 -310 5 VGND
port 4 s
rlabel locali 160 -55 160 -55 3 Y
port 2 e
<< end >>
