magic
tech sky130A
timestamp 1731569169
<< nwell >>
rect 2765 1450 2955 1610
<< pwell >>
rect 2775 1330 2955 1420
<< psubdiff >>
rect 2890 1390 2930 1405
rect 2890 1370 2900 1390
rect 2920 1370 2930 1390
rect 2890 1355 2930 1370
<< nsubdiff >>
rect 2890 1540 2930 1555
rect 2890 1520 2900 1540
rect 2920 1520 2930 1540
rect 2890 1505 2930 1520
<< psubdiffcont >>
rect 2900 1370 2920 1390
<< nsubdiffcont >>
rect 2900 1520 2920 1540
<< locali >>
rect 390 3475 830 3515
rect 3395 1925 4460 1950
rect 3395 1905 4375 1925
rect 4395 1905 4425 1925
rect 4445 1905 4460 1925
rect 3395 1880 4460 1905
rect 2890 1540 2930 1555
rect 2890 1520 2900 1540
rect 2920 1520 2930 1540
rect 2890 1505 2930 1520
rect 2495 1455 2575 1485
rect 2780 1475 2805 1485
rect 2790 1455 2805 1475
rect 2780 1435 2805 1455
rect 2995 1475 3045 1485
rect 2995 1445 3005 1475
rect 3035 1445 3045 1475
rect 2890 1390 2930 1405
rect 2890 1370 2900 1390
rect 2920 1370 2930 1390
rect 2890 1355 2930 1370
rect 2995 190 3045 1445
rect 2995 140 3360 190
<< viali >>
rect 4375 1905 4395 1925
rect 4425 1905 4445 1925
rect 2900 1520 2920 1540
rect 2770 1455 2790 1475
rect 3005 1445 3035 1475
rect 2755 1370 2772 1387
rect 2900 1370 2920 1390
<< metal1 >>
rect 2555 1685 3045 1735
rect 2565 1615 2615 1685
rect 2890 1540 2930 1685
rect 2890 1520 2900 1540
rect 2920 1520 2930 1540
rect 2890 1505 2930 1520
rect 2745 1475 2805 1495
rect 2745 1455 2770 1475
rect 2790 1465 2805 1475
rect 2995 1475 3045 1685
rect 2995 1465 3005 1475
rect 2790 1455 3005 1465
rect 2745 1445 3005 1455
rect 3035 1445 3045 1475
rect 2745 1435 3045 1445
rect 2740 1400 2785 1410
rect 2445 1387 2785 1400
rect 2445 1370 2755 1387
rect 2772 1370 2785 1387
rect 2445 1115 2495 1370
rect 2740 1365 2785 1370
rect 2890 1390 2930 1405
rect 3185 1390 3235 2100
rect 4360 1925 4460 1950
rect 4360 1905 4375 1925
rect 4395 1905 4425 1925
rect 4445 1905 4460 1925
rect 4360 1880 4460 1905
rect 4200 1710 4250 1860
rect 4270 1535 4300 1565
rect 2890 1370 2900 1390
rect 2920 1370 3235 1390
rect 2890 1360 3235 1370
rect 2890 1355 2930 1360
rect 3185 1325 3235 1360
rect 2785 1295 3235 1325
rect 2975 1075 3300 1125
rect 2975 440 3320 490
use sky130_fd_sc_hd__einvp_1  sky130_fd_sc_hd__einvp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 2564 0 1 1319
box -19 -24 249 296
use x5s_cc_osc  x5s_cc_osc_0
timestamp 1731473449
transform 1 0 300 0 1 2100
box -300 -1950 10020 1415
<< labels >>
rlabel locali 2510 1485 2510 1485 1 ENB
port 2 n
rlabel metal1 3065 490 3065 490 1 p[4]
port 3 n
rlabel locali 575 3515 575 3515 1 VDDA
port 4 n
rlabel metal1 3155 1125 3155 1125 1 pn[4]
rlabel metal1 4430 1950 4430 1950 1 Anlg_in
port 1 n
rlabel metal1 4285 1565 4285 1565 1 GND
port 5 n
<< end >>
