magic
tech sky130A
timestamp 1730452893
<< nwell >>
rect 1350 510 1370 530
<< pmos >>
rect 360 600 395 640
<< pdiffc >>
rect 1040 590 1060 610
rect 1350 510 1370 530
<< poly >>
rect 995 360 1005 410
<< polycont >>
rect 610 375 635 400
rect 655 375 680 400
rect 920 375 945 400
rect 970 375 995 400
<< locali >>
rect 335 830 1120 870
rect 490 735 530 830
rect 800 735 840 830
rect 600 400 695 410
rect 600 375 610 400
rect 635 375 655 400
rect 680 375 695 400
rect 600 360 695 375
rect 760 400 1005 410
rect 760 375 920 400
rect 945 375 970 400
rect 995 375 1005 400
rect 760 360 1005 375
rect 560 40 600 130
rect 870 40 910 130
rect 300 0 1155 40
<< viali >>
rect 260 630 280 650
rect 1040 630 1060 650
rect 260 590 280 610
rect 1040 590 1060 610
rect 1350 510 1370 530
rect 1350 470 1370 490
rect 610 375 635 400
rect 655 375 680 400
rect 920 375 945 400
rect 970 375 995 400
rect 1350 260 1370 280
rect 1350 220 1370 240
rect 1350 180 1370 200
<< metal1 >>
rect 250 650 290 660
rect 250 630 260 650
rect 280 640 290 650
rect 1030 650 1070 660
rect 1030 640 1040 650
rect 280 630 1040 640
rect 1060 630 1070 650
rect 250 620 1070 630
rect 0 580 195 620
rect 250 610 1560 620
rect 250 590 260 610
rect 280 600 1040 610
rect 280 590 290 600
rect 250 580 290 590
rect 155 405 195 580
rect 490 410 530 600
rect 1030 590 1040 600
rect 1060 590 1560 610
rect 1030 580 1560 590
rect 1340 530 1380 540
rect 1340 520 1350 530
rect 945 510 1350 520
rect 1370 510 1380 530
rect 945 490 1380 510
rect 945 475 1350 490
rect 945 410 990 475
rect 1340 470 1350 475
rect 1370 470 1380 490
rect 1340 460 1380 470
rect 490 400 720 410
rect 490 375 610 400
rect 635 375 655 400
rect 680 375 720 400
rect 490 360 720 375
rect 910 400 1005 410
rect 910 375 920 400
rect 945 375 970 400
rect 995 375 1005 400
rect 910 360 1005 375
rect 1110 360 1250 405
rect 1110 250 1150 360
rect 0 210 1150 250
rect 1340 280 1380 290
rect 1340 260 1350 280
rect 1370 260 1380 280
rect 1340 250 1380 260
rect 1340 240 1560 250
rect 1340 220 1350 240
rect 1370 220 1560 240
rect 1340 210 1560 220
rect 1340 200 1380 210
rect 1340 180 1350 200
rect 1370 180 1380 200
rect 1340 170 1380 180
use aux_inv_dco  aux_inv_dco_0
timestamp 1730450942
transform 1 0 600 0 1 440
box -130 -350 180 340
use aux_inv_dco  aux_inv_dco_1
timestamp 1730450942
transform 1 0 910 0 1 440
box -130 -350 180 340
use main_inv_dco  main_inv_dco_0
timestamp 1730450826
transform 1 0 130 0 1 440
box -130 -440 340 430
use main_inv_dco  main_inv_dco_1
timestamp 1730450826
transform 1 0 1220 0 1 440
box -130 -440 340 430
<< labels >>
rlabel metal1 0 600 0 600 7 inp
port 1 w
rlabel metal1 0 230 0 230 7 inn
port 2 w
rlabel metal1 1560 600 1560 600 3 outp
port 3 e
rlabel metal1 1560 230 1560 230 3 outn
port 4 e
rlabel locali 490 870 490 870 1 VDDA
port 5 n
rlabel locali 485 0 485 0 5 VGND
port 6 s
<< end >>
