magic
tech sky130A
magscale 1 2
timestamp 1731030357
<< nwell >>
rect 1066 186309 185970 186630
rect 1066 185221 185970 185787
rect 1066 184133 185970 184699
rect 1066 183045 185970 183611
rect 1066 181957 185970 182523
rect 1066 180869 185970 181435
rect 1066 179781 185970 180347
rect 1066 178693 185970 179259
rect 1066 177605 185970 178171
rect 1066 176517 185970 177083
rect 1066 175429 185970 175995
rect 1066 174341 185970 174907
rect 1066 173253 185970 173819
rect 1066 172165 185970 172731
rect 1066 171077 185970 171643
rect 1066 169989 185970 170555
rect 1066 168901 185970 169467
rect 1066 167813 185970 168379
rect 1066 166725 185970 167291
rect 1066 165637 185970 166203
rect 1066 164549 185970 165115
rect 1066 163461 185970 164027
rect 1066 162373 185970 162939
rect 1066 161285 185970 161851
rect 1066 160197 185970 160763
rect 1066 159109 185970 159675
rect 1066 158021 185970 158587
rect 1066 156933 185970 157499
rect 1066 155845 185970 156411
rect 1066 154757 185970 155323
rect 1066 153669 185970 154235
rect 1066 152581 185970 153147
rect 1066 151493 185970 152059
rect 1066 150405 185970 150971
rect 1066 149317 185970 149883
rect 1066 148229 185970 148795
rect 1066 147141 185970 147707
rect 1066 146053 185970 146619
rect 1066 144965 185970 145531
rect 1066 143877 185970 144443
rect 1066 142789 185970 143355
rect 1066 141701 185970 142267
rect 1066 140613 185970 141179
rect 1066 139525 185970 140091
rect 1066 138437 185970 139003
rect 1066 137349 185970 137915
rect 1066 136261 185970 136827
rect 1066 135173 185970 135739
rect 1066 134085 185970 134651
rect 1066 132997 185970 133563
rect 1066 131909 185970 132475
rect 1066 130821 185970 131387
rect 1066 129733 185970 130299
rect 1066 128645 185970 129211
rect 1066 127557 185970 128123
rect 1066 126469 185970 127035
rect 1066 125381 185970 125947
rect 1066 124293 185970 124859
rect 1066 123205 185970 123771
rect 1066 122117 185970 122683
rect 1066 121029 185970 121595
rect 1066 119941 185970 120507
rect 1066 118853 185970 119419
rect 1066 117765 185970 118331
rect 1066 116677 185970 117243
rect 1066 115589 185970 116155
rect 1066 114501 185970 115067
rect 1066 113413 185970 113979
rect 1066 112325 185970 112891
rect 1066 111237 185970 111803
rect 1066 110149 185970 110715
rect 1066 109061 185970 109627
rect 1066 107973 185970 108539
rect 1066 106885 185970 107451
rect 1066 105797 185970 106363
rect 1066 104709 185970 105275
rect 1066 103621 185970 104187
rect 1066 102533 185970 103099
rect 1066 101445 185970 102011
rect 1066 100357 185970 100923
rect 1066 99269 185970 99835
rect 1066 98181 185970 98747
rect 1066 97093 185970 97659
rect 1066 96005 185970 96571
rect 1066 94917 185970 95483
rect 1066 93829 185970 94395
rect 1066 92741 185970 93307
rect 1066 91653 185970 92219
rect 1066 90565 185970 91131
rect 1066 89477 185970 90043
rect 1066 88389 185970 88955
rect 1066 87301 185970 87867
rect 1066 86213 185970 86779
rect 1066 85125 185970 85691
rect 1066 84037 185970 84603
rect 1066 82949 185970 83515
rect 1066 81861 185970 82427
rect 1066 80773 185970 81339
rect 1066 79685 185970 80251
rect 1066 78597 185970 79163
rect 1066 77509 185970 78075
rect 1066 76421 185970 76987
rect 1066 75333 185970 75899
rect 1066 74245 185970 74811
rect 1066 73157 185970 73723
rect 1066 72069 185970 72635
rect 1066 70981 185970 71547
rect 1066 69893 185970 70459
rect 1066 68805 185970 69371
rect 1066 67717 185970 68283
rect 1066 66629 185970 67195
rect 1066 65541 185970 66107
rect 1066 64453 185970 65019
rect 1066 63365 185970 63931
rect 1066 62277 185970 62843
rect 1066 61189 185970 61755
rect 1066 60101 185970 60667
rect 1066 59013 185970 59579
rect 1066 57925 185970 58491
rect 1066 56837 185970 57403
rect 1066 55749 185970 56315
rect 1066 54661 185970 55227
rect 1066 53573 185970 54139
rect 1066 52485 185970 53051
rect 1066 51397 185970 51963
rect 1066 50309 185970 50875
rect 1066 49221 185970 49787
rect 1066 48133 185970 48699
rect 1066 47045 185970 47611
rect 1066 45957 185970 46523
rect 1066 44869 185970 45435
rect 1066 43781 185970 44347
rect 1066 42693 185970 43259
rect 1066 41605 185970 42171
rect 1066 40517 185970 41083
rect 1066 39429 185970 39995
rect 1066 38341 185970 38907
rect 1066 37253 185970 37819
rect 1066 36165 185970 36731
rect 1066 35077 185970 35643
rect 1066 33989 185970 34555
rect 1066 32901 185970 33467
rect 1066 31813 185970 32379
rect 1066 30725 185970 31291
rect 1066 29637 185970 30203
rect 1066 28549 185970 29115
rect 1066 27461 185970 28027
rect 1066 26373 185970 26939
rect 1066 25285 185970 25851
rect 1066 24197 185970 24763
rect 1066 23109 185970 23675
rect 1066 22021 185970 22587
rect 1066 20933 185970 21499
rect 1066 19845 185970 20411
rect 1066 18757 185970 19323
rect 1066 17669 185970 18235
rect 1066 16581 185970 17147
rect 1066 15493 185970 16059
rect 1066 14405 185970 14971
rect 1066 13317 185970 13883
rect 1066 12229 185970 12795
rect 1066 11141 185970 11707
rect 1066 10053 185970 10619
rect 1066 8965 185970 9531
rect 1066 7877 185970 8443
rect 1066 6789 185970 7355
rect 1066 5701 185970 6267
rect 1066 4613 185970 5179
rect 1066 3525 185970 4091
rect 1066 2437 185970 3003
<< obsli1 >>
rect 1104 2159 185932 186609
<< obsm1 >>
rect 1104 1368 185932 186640
<< metal2 >>
rect 1490 0 1546 800
rect 3790 0 3846 800
rect 6090 0 6146 800
rect 8390 0 8446 800
rect 10690 0 10746 800
rect 12990 0 13046 800
rect 15290 0 15346 800
rect 17590 0 17646 800
rect 19890 0 19946 800
rect 22190 0 22246 800
rect 24490 0 24546 800
rect 26790 0 26846 800
rect 29090 0 29146 800
rect 31390 0 31446 800
rect 33690 0 33746 800
rect 35990 0 36046 800
rect 38290 0 38346 800
rect 40590 0 40646 800
rect 42890 0 42946 800
rect 45190 0 45246 800
rect 47490 0 47546 800
rect 49790 0 49846 800
rect 52090 0 52146 800
rect 54390 0 54446 800
rect 56690 0 56746 800
rect 58990 0 59046 800
rect 61290 0 61346 800
rect 63590 0 63646 800
rect 65890 0 65946 800
rect 68190 0 68246 800
rect 70490 0 70546 800
rect 72790 0 72846 800
rect 75090 0 75146 800
rect 77390 0 77446 800
rect 79690 0 79746 800
rect 81990 0 82046 800
rect 84290 0 84346 800
rect 86590 0 86646 800
rect 88890 0 88946 800
rect 91190 0 91246 800
rect 93490 0 93546 800
rect 95790 0 95846 800
rect 98090 0 98146 800
rect 100390 0 100446 800
rect 102690 0 102746 800
rect 104990 0 105046 800
rect 107290 0 107346 800
rect 109590 0 109646 800
rect 111890 0 111946 800
rect 114190 0 114246 800
rect 116490 0 116546 800
rect 118790 0 118846 800
rect 121090 0 121146 800
rect 123390 0 123446 800
rect 125690 0 125746 800
rect 127990 0 128046 800
rect 130290 0 130346 800
rect 132590 0 132646 800
rect 134890 0 134946 800
rect 137190 0 137246 800
rect 139490 0 139546 800
rect 141790 0 141846 800
rect 144090 0 144146 800
rect 146390 0 146446 800
rect 148690 0 148746 800
rect 150990 0 151046 800
rect 153290 0 153346 800
rect 155590 0 155646 800
rect 157890 0 157946 800
rect 160190 0 160246 800
rect 162490 0 162546 800
rect 164790 0 164846 800
rect 167090 0 167146 800
rect 169390 0 169446 800
rect 171690 0 171746 800
rect 173990 0 174046 800
rect 176290 0 176346 800
rect 178590 0 178646 800
rect 180890 0 180946 800
rect 183190 0 183246 800
rect 185490 0 185546 800
<< obsm2 >>
rect 1490 856 185532 186629
rect 1602 734 3734 856
rect 3902 734 6034 856
rect 6202 734 8334 856
rect 8502 734 10634 856
rect 10802 734 12934 856
rect 13102 734 15234 856
rect 15402 734 17534 856
rect 17702 734 19834 856
rect 20002 734 22134 856
rect 22302 734 24434 856
rect 24602 734 26734 856
rect 26902 734 29034 856
rect 29202 734 31334 856
rect 31502 734 33634 856
rect 33802 734 35934 856
rect 36102 734 38234 856
rect 38402 734 40534 856
rect 40702 734 42834 856
rect 43002 734 45134 856
rect 45302 734 47434 856
rect 47602 734 49734 856
rect 49902 734 52034 856
rect 52202 734 54334 856
rect 54502 734 56634 856
rect 56802 734 58934 856
rect 59102 734 61234 856
rect 61402 734 63534 856
rect 63702 734 65834 856
rect 66002 734 68134 856
rect 68302 734 70434 856
rect 70602 734 72734 856
rect 72902 734 75034 856
rect 75202 734 77334 856
rect 77502 734 79634 856
rect 79802 734 81934 856
rect 82102 734 84234 856
rect 84402 734 86534 856
rect 86702 734 88834 856
rect 89002 734 91134 856
rect 91302 734 93434 856
rect 93602 734 95734 856
rect 95902 734 98034 856
rect 98202 734 100334 856
rect 100502 734 102634 856
rect 102802 734 104934 856
rect 105102 734 107234 856
rect 107402 734 109534 856
rect 109702 734 111834 856
rect 112002 734 114134 856
rect 114302 734 116434 856
rect 116602 734 118734 856
rect 118902 734 121034 856
rect 121202 734 123334 856
rect 123502 734 125634 856
rect 125802 734 127934 856
rect 128102 734 130234 856
rect 130402 734 132534 856
rect 132702 734 134834 856
rect 135002 734 137134 856
rect 137302 734 139434 856
rect 139602 734 141734 856
rect 141902 734 144034 856
rect 144202 734 146334 856
rect 146502 734 148634 856
rect 148802 734 150934 856
rect 151102 734 153234 856
rect 153402 734 155534 856
rect 155702 734 157834 856
rect 158002 734 160134 856
rect 160302 734 162434 856
rect 162602 734 164734 856
rect 164902 734 167034 856
rect 167202 734 169334 856
rect 169502 734 171634 856
rect 171802 734 173934 856
rect 174102 734 176234 856
rect 176402 734 178534 856
rect 178702 734 180834 856
rect 181002 734 183134 856
rect 183302 734 185434 856
<< obsm3 >>
rect 1485 1942 180123 186625
<< metal4 >>
rect 4208 2128 4528 186640
rect 19568 2128 19888 186640
rect 34928 2128 35248 186640
rect 50288 2128 50608 186640
rect 65648 2128 65968 186640
rect 81008 2128 81328 186640
rect 96368 2128 96688 186640
rect 111728 2128 112048 186640
rect 127088 2128 127408 186640
rect 142448 2128 142768 186640
rect 157808 2128 158128 186640
rect 173168 2128 173488 186640
<< obsm4 >>
rect 3003 2075 4128 171733
rect 4608 2075 19488 171733
rect 19968 2075 34848 171733
rect 35328 2075 50208 171733
rect 50688 2075 65568 171733
rect 66048 2075 80928 171733
rect 81408 2075 96288 171733
rect 96768 2075 111648 171733
rect 112128 2075 127008 171733
rect 127488 2075 142368 171733
rect 142848 2075 157728 171733
rect 158208 2075 173088 171733
rect 173568 2075 179157 171733
<< labels >>
rlabel metal2 s 31390 0 31446 800 6 becStatus[0]
port 1 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 becStatus[1]
port 2 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 becStatus[2]
port 3 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 becStatus[3]
port 4 nsew signal output
rlabel metal2 s 1490 0 1546 800 6 clk
port 5 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 data_in[0]
port 6 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 data_in[10]
port 7 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 data_in[11]
port 8 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 data_in[12]
port 9 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 data_in[13]
port 10 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 data_in[14]
port 11 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 data_in[15]
port 12 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 data_in[16]
port 13 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 data_in[17]
port 14 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 data_in[18]
port 15 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 data_in[19]
port 16 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 data_in[1]
port 17 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 data_in[20]
port 18 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 data_in[21]
port 19 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 data_in[22]
port 20 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 data_in[23]
port 21 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 data_in[24]
port 22 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 data_in[25]
port 23 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 data_in[26]
port 24 nsew signal input
rlabel metal2 s 164790 0 164846 800 6 data_in[27]
port 25 nsew signal input
rlabel metal2 s 169390 0 169446 800 6 data_in[28]
port 26 nsew signal input
rlabel metal2 s 173990 0 174046 800 6 data_in[29]
port 27 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 data_in[2]
port 28 nsew signal input
rlabel metal2 s 178590 0 178646 800 6 data_in[30]
port 29 nsew signal input
rlabel metal2 s 183190 0 183246 800 6 data_in[31]
port 30 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 data_in[3]
port 31 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 data_in[4]
port 32 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 data_in[5]
port 33 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 data_in[6]
port 34 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 data_in[7]
port 35 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 data_in[8]
port 36 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 data_in[9]
port 37 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 data_out[0]
port 38 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 data_out[10]
port 39 nsew signal output
rlabel metal2 s 93490 0 93546 800 6 data_out[11]
port 40 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 data_out[12]
port 41 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 data_out[13]
port 42 nsew signal output
rlabel metal2 s 107290 0 107346 800 6 data_out[14]
port 43 nsew signal output
rlabel metal2 s 111890 0 111946 800 6 data_out[15]
port 44 nsew signal output
rlabel metal2 s 116490 0 116546 800 6 data_out[16]
port 45 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 data_out[17]
port 46 nsew signal output
rlabel metal2 s 125690 0 125746 800 6 data_out[18]
port 47 nsew signal output
rlabel metal2 s 130290 0 130346 800 6 data_out[19]
port 48 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 data_out[1]
port 49 nsew signal output
rlabel metal2 s 134890 0 134946 800 6 data_out[20]
port 50 nsew signal output
rlabel metal2 s 139490 0 139546 800 6 data_out[21]
port 51 nsew signal output
rlabel metal2 s 144090 0 144146 800 6 data_out[22]
port 52 nsew signal output
rlabel metal2 s 148690 0 148746 800 6 data_out[23]
port 53 nsew signal output
rlabel metal2 s 153290 0 153346 800 6 data_out[24]
port 54 nsew signal output
rlabel metal2 s 157890 0 157946 800 6 data_out[25]
port 55 nsew signal output
rlabel metal2 s 162490 0 162546 800 6 data_out[26]
port 56 nsew signal output
rlabel metal2 s 167090 0 167146 800 6 data_out[27]
port 57 nsew signal output
rlabel metal2 s 171690 0 171746 800 6 data_out[28]
port 58 nsew signal output
rlabel metal2 s 176290 0 176346 800 6 data_out[29]
port 59 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 data_out[2]
port 60 nsew signal output
rlabel metal2 s 180890 0 180946 800 6 data_out[30]
port 61 nsew signal output
rlabel metal2 s 185490 0 185546 800 6 data_out[31]
port 62 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 data_out[3]
port 63 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 data_out[4]
port 64 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 data_out[5]
port 65 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 data_out[6]
port 66 nsew signal output
rlabel metal2 s 75090 0 75146 800 6 data_out[7]
port 67 nsew signal output
rlabel metal2 s 79690 0 79746 800 6 data_out[8]
port 68 nsew signal output
rlabel metal2 s 84290 0 84346 800 6 data_out[9]
port 69 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 done
port 70 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 enable
port 71 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 ki
port 72 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 load_data
port 73 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 load_status[0]
port 74 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 load_status[1]
port 75 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 load_status[2]
port 76 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 load_status[3]
port 77 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 load_status[4]
port 78 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 load_status[5]
port 79 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 next_key
port 80 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 rst
port 81 nsew signal input
rlabel metal4 s 4208 2128 4528 186640 6 vccd2
port 82 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 186640 6 vccd2
port 82 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 186640 6 vccd2
port 82 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 186640 6 vccd2
port 82 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 186640 6 vccd2
port 82 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 186640 6 vccd2
port 82 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 186640 6 vssd2
port 83 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 186640 6 vssd2
port 83 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 186640 6 vssd2
port 83 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 186640 6 vssd2
port 83 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 186640 6 vssd2
port 83 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 186640 6 vssd2
port 83 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 187041 189185
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 60521196
string GDS_FILE /home/admin/projects/IC5-CASS-2024/openlane/lovers_bec/runs/24_11_08_08_08/results/signoff/bec.magic.gds
string GDS_START 910170
<< end >>

