magic
tech sky130A
magscale 1 2
timestamp 1731514826
<< obsli1 >>
rect 1104 2159 28888 27761
<< obsm1 >>
rect 842 2128 29150 27792
<< metal2 >>
rect 846 0 902 800
rect 1674 0 1730 800
rect 2502 0 2558 800
rect 3330 0 3386 800
rect 4158 0 4214 800
rect 4986 0 5042 800
rect 5814 0 5870 800
rect 6642 0 6698 800
rect 7470 0 7526 800
rect 8298 0 8354 800
rect 9126 0 9182 800
rect 9954 0 10010 800
rect 10782 0 10838 800
rect 11610 0 11666 800
rect 12438 0 12494 800
rect 13266 0 13322 800
rect 14094 0 14150 800
rect 14922 0 14978 800
rect 15750 0 15806 800
rect 16578 0 16634 800
rect 17406 0 17462 800
rect 18234 0 18290 800
rect 19062 0 19118 800
rect 19890 0 19946 800
rect 20718 0 20774 800
rect 21546 0 21602 800
rect 22374 0 22430 800
rect 23202 0 23258 800
rect 24030 0 24086 800
rect 24858 0 24914 800
rect 25686 0 25742 800
rect 26514 0 26570 800
rect 27342 0 27398 800
rect 28170 0 28226 800
rect 28998 0 29054 800
<< obsm2 >>
rect 848 856 29144 27781
rect 958 734 1618 856
rect 1786 734 2446 856
rect 2614 734 3274 856
rect 3442 734 4102 856
rect 4270 734 4930 856
rect 5098 734 5758 856
rect 5926 734 6586 856
rect 6754 734 7414 856
rect 7582 734 8242 856
rect 8410 734 9070 856
rect 9238 734 9898 856
rect 10066 734 10726 856
rect 10894 734 11554 856
rect 11722 734 12382 856
rect 12550 734 13210 856
rect 13378 734 14038 856
rect 14206 734 14866 856
rect 15034 734 15694 856
rect 15862 734 16522 856
rect 16690 734 17350 856
rect 17518 734 18178 856
rect 18346 734 19006 856
rect 19174 734 19834 856
rect 20002 734 20662 856
rect 20830 734 21490 856
rect 21658 734 22318 856
rect 22486 734 23146 856
rect 23314 734 23974 856
rect 24142 734 24802 856
rect 24970 734 25630 856
rect 25798 734 26458 856
rect 26626 734 27286 856
rect 27454 734 28114 856
rect 28282 734 28942 856
rect 29110 734 29144 856
<< obsm3 >>
rect 4245 2143 29046 27777
<< metal4 >>
rect 4417 2128 4737 27792
rect 7890 2128 8210 27792
rect 11363 2128 11683 27792
rect 14836 2128 15156 27792
rect 18309 2128 18629 27792
rect 21782 2128 22102 27792
rect 25255 2128 25575 27792
rect 28728 2128 29048 27792
<< obsm4 >>
rect 18827 16491 18893 19413
<< labels >>
rlabel metal2 s 3330 0 3386 800 6 a[0]
port 1 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 a[1]
port 2 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 a[2]
port 3 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 a[3]
port 4 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 a[4]
port 5 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 a[5]
port 6 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 a[6]
port 7 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 a[7]
port 8 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 b[0]
port 9 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 b[1]
port 10 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 b[2]
port 11 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 b[3]
port 12 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 b[4]
port 13 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 b[5]
port 14 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 b[6]
port 15 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 b[7]
port 16 nsew signal input
rlabel metal2 s 846 0 902 800 6 clk
port 17 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 control
port 18 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 p[0]
port 19 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 p[10]
port 20 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 p[11]
port 21 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 p[12]
port 22 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 p[13]
port 23 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 p[14]
port 24 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 p[15]
port 25 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 p[1]
port 26 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 p[2]
port 27 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 p[3]
port 28 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 p[4]
port 29 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 p[5]
port 30 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 p[6]
port 31 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 p[7]
port 32 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 p[8]
port 33 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 p[9]
port 34 nsew signal output
rlabel metal2 s 1674 0 1730 800 6 rst
port 35 nsew signal input
rlabel metal4 s 4417 2128 4737 27792 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 11363 2128 11683 27792 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 18309 2128 18629 27792 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 25255 2128 25575 27792 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 7890 2128 8210 27792 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 14836 2128 15156 27792 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 21782 2128 22102 27792 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 28728 2128 29048 27792 6 vssd1
port 37 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2270348
string GDS_FILE /home/cass/projects/IC5-CASS-2024/openlane/vmsu_8bit/runs/24_11_13_23_16/results/signoff/vmsu_8bit_top.magic.gds
string GDS_START 313678
<< end >>

