VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ascon_wrapper
  CLASS BLOCK ;
  FOREIGN ascon_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 540.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 449.050 536.000 449.330 540.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 515.480 600.000 516.080 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 425.720 600.000 426.320 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 335.960 600.000 336.560 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 246.200 600.000 246.800 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 156.440 600.000 157.040 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 66.680 600.000 67.280 ;
    END
  END io_in[5]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 536.000 269.930 540.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 536.000 389.530 540.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 536.000 150.330 540.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 536.000 30.730 540.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 470.600 600.000 471.200 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 380.840 600.000 381.440 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 291.080 600.000 291.680 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 201.320 600.000 201.920 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 111.560 600.000 112.160 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 21.800 600.000 22.400 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 536.000 509.130 540.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 329.450 536.000 329.730 540.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 209.850 536.000 210.130 540.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 90.250 536.000 90.530 540.000 ;
    END
  END io_out[2]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 568.650 536.000 568.930 540.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 527.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 527.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 527.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 527.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 527.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 527.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 527.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 527.920 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 523.545 594.510 526.375 ;
        RECT 5.330 518.105 594.510 520.935 ;
        RECT 5.330 512.665 594.510 515.495 ;
        RECT 5.330 507.225 594.510 510.055 ;
        RECT 5.330 501.785 594.510 504.615 ;
        RECT 5.330 496.345 594.510 499.175 ;
        RECT 5.330 490.905 594.510 493.735 ;
        RECT 5.330 485.465 594.510 488.295 ;
        RECT 5.330 480.025 594.510 482.855 ;
        RECT 5.330 474.585 594.510 477.415 ;
        RECT 5.330 469.145 594.510 471.975 ;
        RECT 5.330 463.705 594.510 466.535 ;
        RECT 5.330 458.265 594.510 461.095 ;
        RECT 5.330 452.825 594.510 455.655 ;
        RECT 5.330 447.385 594.510 450.215 ;
        RECT 5.330 441.945 594.510 444.775 ;
        RECT 5.330 436.505 594.510 439.335 ;
        RECT 5.330 431.065 594.510 433.895 ;
        RECT 5.330 425.625 594.510 428.455 ;
        RECT 5.330 420.185 594.510 423.015 ;
        RECT 5.330 414.745 594.510 417.575 ;
        RECT 5.330 409.305 594.510 412.135 ;
        RECT 5.330 403.865 594.510 406.695 ;
        RECT 5.330 398.425 594.510 401.255 ;
        RECT 5.330 392.985 594.510 395.815 ;
        RECT 5.330 387.545 594.510 390.375 ;
        RECT 5.330 382.105 594.510 384.935 ;
        RECT 5.330 376.665 594.510 379.495 ;
        RECT 5.330 371.225 594.510 374.055 ;
        RECT 5.330 365.785 594.510 368.615 ;
        RECT 5.330 360.345 594.510 363.175 ;
        RECT 5.330 354.905 594.510 357.735 ;
        RECT 5.330 349.465 594.510 352.295 ;
        RECT 5.330 344.025 594.510 346.855 ;
        RECT 5.330 338.585 594.510 341.415 ;
        RECT 5.330 333.145 594.510 335.975 ;
        RECT 5.330 327.705 594.510 330.535 ;
        RECT 5.330 322.265 594.510 325.095 ;
        RECT 5.330 316.825 594.510 319.655 ;
        RECT 5.330 311.385 594.510 314.215 ;
        RECT 5.330 305.945 594.510 308.775 ;
        RECT 5.330 300.505 594.510 303.335 ;
        RECT 5.330 295.065 594.510 297.895 ;
        RECT 5.330 289.625 594.510 292.455 ;
        RECT 5.330 284.185 594.510 287.015 ;
        RECT 5.330 278.745 594.510 281.575 ;
        RECT 5.330 273.305 594.510 276.135 ;
        RECT 5.330 267.865 594.510 270.695 ;
        RECT 5.330 262.425 594.510 265.255 ;
        RECT 5.330 256.985 594.510 259.815 ;
        RECT 5.330 251.545 594.510 254.375 ;
        RECT 5.330 246.105 594.510 248.935 ;
        RECT 5.330 240.665 594.510 243.495 ;
        RECT 5.330 235.225 594.510 238.055 ;
        RECT 5.330 229.785 594.510 232.615 ;
        RECT 5.330 224.345 594.510 227.175 ;
        RECT 5.330 218.905 594.510 221.735 ;
        RECT 5.330 213.465 594.510 216.295 ;
        RECT 5.330 208.025 594.510 210.855 ;
        RECT 5.330 202.585 594.510 205.415 ;
        RECT 5.330 197.145 594.510 199.975 ;
        RECT 5.330 191.705 594.510 194.535 ;
        RECT 5.330 186.265 594.510 189.095 ;
        RECT 5.330 180.825 594.510 183.655 ;
        RECT 5.330 175.385 594.510 178.215 ;
        RECT 5.330 169.945 594.510 172.775 ;
        RECT 5.330 164.505 594.510 167.335 ;
        RECT 5.330 159.065 594.510 161.895 ;
        RECT 5.330 153.625 594.510 156.455 ;
        RECT 5.330 148.185 594.510 151.015 ;
        RECT 5.330 142.745 594.510 145.575 ;
        RECT 5.330 137.305 594.510 140.135 ;
        RECT 5.330 131.865 594.510 134.695 ;
        RECT 5.330 126.425 594.510 129.255 ;
        RECT 5.330 120.985 594.510 123.815 ;
        RECT 5.330 115.545 594.510 118.375 ;
        RECT 5.330 110.105 594.510 112.935 ;
        RECT 5.330 104.665 594.510 107.495 ;
        RECT 5.330 99.225 594.510 102.055 ;
        RECT 5.330 93.785 594.510 96.615 ;
        RECT 5.330 88.345 594.510 91.175 ;
        RECT 5.330 82.905 594.510 85.735 ;
        RECT 5.330 77.465 594.510 80.295 ;
        RECT 5.330 72.025 594.510 74.855 ;
        RECT 5.330 66.585 594.510 69.415 ;
        RECT 5.330 61.145 594.510 63.975 ;
        RECT 5.330 55.705 594.510 58.535 ;
        RECT 5.330 50.265 594.510 53.095 ;
        RECT 5.330 44.825 594.510 47.655 ;
        RECT 5.330 39.385 594.510 42.215 ;
        RECT 5.330 33.945 594.510 36.775 ;
        RECT 5.330 28.505 594.510 31.335 ;
        RECT 5.330 23.065 594.510 25.895 ;
        RECT 5.330 17.625 594.510 20.455 ;
        RECT 5.330 12.185 594.510 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 594.320 527.765 ;
      LAYER met1 ;
        RECT 5.520 10.640 594.710 527.920 ;
      LAYER met2 ;
        RECT 19.880 535.720 30.170 536.000 ;
        RECT 31.010 535.720 89.970 536.000 ;
        RECT 90.810 535.720 149.770 536.000 ;
        RECT 150.610 535.720 209.570 536.000 ;
        RECT 210.410 535.720 269.370 536.000 ;
        RECT 270.210 535.720 329.170 536.000 ;
        RECT 330.010 535.720 388.970 536.000 ;
        RECT 389.810 535.720 448.770 536.000 ;
        RECT 449.610 535.720 508.570 536.000 ;
        RECT 509.410 535.720 568.370 536.000 ;
        RECT 569.210 535.720 594.690 536.000 ;
        RECT 19.880 10.695 594.690 535.720 ;
      LAYER met3 ;
        RECT 21.050 516.480 596.000 527.845 ;
        RECT 21.050 515.080 595.600 516.480 ;
        RECT 21.050 471.600 596.000 515.080 ;
        RECT 21.050 470.200 595.600 471.600 ;
        RECT 21.050 426.720 596.000 470.200 ;
        RECT 21.050 425.320 595.600 426.720 ;
        RECT 21.050 381.840 596.000 425.320 ;
        RECT 21.050 380.440 595.600 381.840 ;
        RECT 21.050 336.960 596.000 380.440 ;
        RECT 21.050 335.560 595.600 336.960 ;
        RECT 21.050 292.080 596.000 335.560 ;
        RECT 21.050 290.680 595.600 292.080 ;
        RECT 21.050 247.200 596.000 290.680 ;
        RECT 21.050 245.800 595.600 247.200 ;
        RECT 21.050 202.320 596.000 245.800 ;
        RECT 21.050 200.920 595.600 202.320 ;
        RECT 21.050 157.440 596.000 200.920 ;
        RECT 21.050 156.040 595.600 157.440 ;
        RECT 21.050 112.560 596.000 156.040 ;
        RECT 21.050 111.160 595.600 112.560 ;
        RECT 21.050 67.680 596.000 111.160 ;
        RECT 21.050 66.280 595.600 67.680 ;
        RECT 21.050 22.800 596.000 66.280 ;
        RECT 21.050 21.400 595.600 22.800 ;
        RECT 21.050 10.715 596.000 21.400 ;
      LAYER met4 ;
        RECT 72.055 36.895 97.440 499.625 ;
        RECT 99.840 36.895 174.240 499.625 ;
        RECT 176.640 36.895 251.040 499.625 ;
        RECT 253.440 36.895 327.840 499.625 ;
        RECT 330.240 36.895 404.640 499.625 ;
        RECT 407.040 36.895 481.440 499.625 ;
        RECT 483.840 36.895 558.240 499.625 ;
        RECT 560.640 36.895 578.385 499.625 ;
      LAYER met5 ;
        RECT 122.940 170.900 421.700 342.500 ;
  END
END ascon_wrapper
END LIBRARY

